//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 0 0 1 0 0 1 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968;
  XNOR2_X1  g000(.A(KEYINPUT0), .B(G57gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G85gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G1gat), .B(G29gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(G134gat), .ZN(new_n206));
  INV_X1    g005(.A(G127gat), .ZN(new_n207));
  INV_X1    g006(.A(G120gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G113gat), .ZN(new_n209));
  INV_X1    g008(.A(G113gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G120gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n207), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI211_X1 g013(.A(KEYINPUT1), .B(G127gat), .C1(new_n209), .C2(new_n211), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n206), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G141gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n217), .A2(G148gat), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT73), .B(G141gat), .ZN(new_n220));
  INV_X1    g019(.A(G148gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G162gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G155gat), .ZN(new_n224));
  INV_X1    g023(.A(G155gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G162gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n228), .B1(KEYINPUT74), .B2(G162gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n221), .A2(G141gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n228), .B1(new_n218), .B2(new_n231), .ZN(new_n232));
  AOI22_X1  g031(.A1(new_n222), .A2(new_n230), .B1(new_n232), .B2(new_n227), .ZN(new_n233));
  XNOR2_X1  g032(.A(G113gat), .B(G120gat), .ZN(new_n234));
  OAI21_X1  g033(.A(G127gat), .B1(new_n234), .B2(KEYINPUT1), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n212), .A2(new_n213), .A3(new_n207), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(new_n236), .A3(G134gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n216), .A2(new_n233), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT75), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT75), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n216), .A2(new_n233), .A3(new_n240), .A4(new_n237), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(KEYINPUT4), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT76), .ZN(new_n243));
  OR2_X1    g042(.A1(new_n238), .A2(KEYINPUT4), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT76), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n239), .A2(new_n245), .A3(KEYINPUT4), .A4(new_n241), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n243), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G225gat), .A2(G233gat), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n249), .A2(KEYINPUT5), .ZN(new_n250));
  INV_X1    g049(.A(new_n233), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n216), .A2(new_n237), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n233), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n252), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n247), .A2(new_n250), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n239), .B(new_n241), .C1(new_n258), .C2(new_n249), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n259), .B(new_n256), .C1(new_n258), .C2(new_n238), .ZN(new_n260));
  INV_X1    g059(.A(new_n253), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n239), .B(new_n241), .C1(new_n261), .C2(new_n233), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n249), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n260), .A2(KEYINPUT5), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n205), .B1(new_n257), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT6), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n257), .A2(new_n264), .A3(new_n205), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT77), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT6), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n265), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n268), .B1(new_n267), .B2(new_n269), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n266), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G78gat), .B(G106gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n275), .B(KEYINPUT31), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(G50gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT78), .ZN(new_n278));
  AND2_X1   g077(.A1(G197gat), .A2(G204gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(G197gat), .A2(G204gat), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT22), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G211gat), .A2(G218gat), .ZN(new_n282));
  INV_X1    g081(.A(G211gat), .ZN(new_n283));
  INV_X1    g082(.A(G218gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n281), .A2(new_n282), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n280), .ZN(new_n287));
  NAND2_X1  g086(.A1(G197gat), .A2(G204gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n283), .A2(new_n284), .A3(KEYINPUT22), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(new_n282), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n286), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT29), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n293), .B1(new_n255), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT29), .B1(new_n286), .B2(new_n292), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n251), .B1(new_n297), .B2(KEYINPUT3), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT81), .ZN(new_n299));
  INV_X1    g098(.A(G228gat), .ZN(new_n300));
  INV_X1    g099(.A(G233gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT81), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n251), .B(new_n303), .C1(KEYINPUT3), .C2(new_n297), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n296), .A2(new_n299), .A3(new_n302), .A4(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G22gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n286), .A2(new_n292), .A3(KEYINPUT79), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n287), .A2(new_n288), .B1(new_n290), .B2(new_n282), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT79), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT29), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT80), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n307), .A2(new_n310), .A3(KEYINPUT80), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n313), .A2(new_n254), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n295), .B1(new_n315), .B2(new_n251), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n305), .B(new_n306), .C1(new_n316), .C2(new_n302), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT3), .B1(new_n311), .B2(new_n312), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n233), .B1(new_n319), .B2(new_n314), .ZN(new_n320));
  OAI22_X1  g119(.A1(new_n320), .A2(new_n295), .B1(new_n300), .B2(new_n301), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n306), .B1(new_n321), .B2(new_n305), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n278), .B1(new_n318), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n305), .B1(new_n316), .B2(new_n302), .ZN(new_n324));
  OR3_X1    g123(.A1(new_n324), .A2(KEYINPUT82), .A3(G22gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(G22gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n326), .A2(KEYINPUT82), .A3(new_n317), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n323), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(new_n277), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT78), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n323), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT27), .B(G183gat), .ZN(new_n334));
  INV_X1    g133(.A(G190gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT69), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT28), .ZN(new_n338));
  NAND2_X1  g137(.A1(G169gat), .A2(G176gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT65), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n344));
  OR3_X1    g143(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G183gat), .A2(G190gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n334), .A2(new_n348), .A3(new_n335), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n338), .A2(new_n346), .A3(new_n347), .A4(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  OR3_X1    g150(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AND3_X1   g153(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT66), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT66), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n358), .B1(new_n341), .B2(new_n342), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n354), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n347), .ZN(new_n362));
  NAND3_X1  g161(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT67), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g164(.A1(KEYINPUT67), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n362), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT25), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n360), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n362), .A2(new_n363), .B1(new_n341), .B2(new_n342), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n371), .B1(new_n372), .B2(new_n354), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT68), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n362), .A2(new_n363), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n375), .A2(new_n354), .A3(new_n343), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n370), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT66), .B1(new_n355), .B2(new_n356), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n341), .A2(new_n358), .A3(new_n342), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n380), .A2(KEYINPUT25), .A3(new_n367), .A4(new_n354), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT68), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n377), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n351), .B1(new_n374), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(G226gat), .A2(G233gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n294), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n377), .A2(new_n381), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n350), .ZN(new_n388));
  OAI22_X1  g187(.A1(new_n384), .A2(new_n386), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n293), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT72), .ZN(new_n392));
  INV_X1    g191(.A(new_n385), .ZN(new_n393));
  AOI211_X1 g192(.A(new_n392), .B(new_n393), .C1(new_n388), .C2(new_n294), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT72), .B1(new_n384), .B2(new_n385), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n393), .B1(new_n388), .B2(new_n294), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n394), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n391), .B1(new_n398), .B2(new_n390), .ZN(new_n399));
  XOR2_X1   g198(.A(G8gat), .B(G36gat), .Z(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(G64gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n401), .B(G92gat), .Z(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n391), .B(new_n402), .C1(new_n398), .C2(new_n390), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(KEYINPUT30), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT30), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n399), .A2(new_n407), .A3(new_n403), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n377), .A2(new_n381), .A3(new_n382), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n382), .B1(new_n377), .B2(new_n381), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n350), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n253), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n261), .B(new_n350), .C1(new_n410), .C2(new_n411), .ZN(new_n414));
  NAND2_X1  g213(.A1(G227gat), .A2(G233gat), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(KEYINPUT34), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT70), .B(G71gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(G99gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(G15gat), .B(G43gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n415), .B1(new_n413), .B2(new_n414), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n421), .B1(new_n422), .B2(KEYINPUT33), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT32), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n413), .A2(new_n414), .ZN(new_n427));
  INV_X1    g226(.A(new_n415), .ZN(new_n428));
  AOI221_X4 g227(.A(new_n424), .B1(KEYINPUT33), .B2(new_n421), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n417), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n427), .A2(new_n428), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT32), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT33), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n432), .A2(new_n434), .A3(new_n421), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT34), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n416), .B(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n423), .A2(new_n425), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n435), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n430), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n274), .A2(new_n333), .A3(new_n409), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT35), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT89), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(KEYINPUT89), .A3(KEYINPUT35), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT83), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n405), .A2(KEYINPUT30), .ZN(new_n447));
  INV_X1    g246(.A(new_n394), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n392), .B1(new_n412), .B2(new_n393), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n448), .B1(new_n449), .B2(new_n396), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n293), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n402), .B1(new_n451), .B2(new_n391), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n408), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n446), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n406), .A2(KEYINPUT83), .A3(new_n408), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n455), .A2(new_n333), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT35), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n267), .A2(new_n269), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n266), .B1(new_n459), .B2(new_n265), .ZN(new_n460));
  OR2_X1    g259(.A1(new_n430), .A2(KEYINPUT71), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n430), .A2(new_n439), .A3(KEYINPUT71), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n457), .A2(new_n458), .A3(new_n460), .A4(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n444), .A2(new_n445), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT85), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n466), .B1(new_n262), .B2(new_n249), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n262), .A2(new_n249), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n247), .A2(new_n256), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n468), .B1(new_n469), .B2(new_n249), .ZN(new_n470));
  OAI211_X1 g269(.A(KEYINPUT39), .B(new_n467), .C1(new_n470), .C2(new_n466), .ZN(new_n471));
  XNOR2_X1  g270(.A(KEYINPUT84), .B(KEYINPUT39), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n469), .A2(new_n249), .A3(new_n472), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n471), .A2(KEYINPUT40), .A3(new_n205), .A4(new_n473), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n474), .A2(new_n271), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n455), .A2(new_n456), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n471), .A2(new_n205), .A3(new_n473), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT40), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n475), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT86), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n481), .B1(new_n398), .B2(new_n293), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n389), .A2(new_n293), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n450), .A2(KEYINPUT86), .A3(new_n390), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT37), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT38), .ZN(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT87), .B(KEYINPUT37), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n403), .B1(new_n399), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n486), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT88), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n451), .A2(KEYINPUT37), .A3(new_n391), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n487), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n493), .A2(new_n460), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT88), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n486), .A2(new_n495), .A3(new_n487), .A4(new_n489), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n491), .A2(new_n494), .A3(new_n404), .A4(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n480), .A2(new_n497), .A3(new_n333), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n333), .B1(new_n274), .B2(new_n409), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT36), .B1(new_n461), .B2(new_n462), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n440), .A2(new_n501), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n499), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n465), .A2(new_n504), .ZN(new_n505));
  XOR2_X1   g304(.A(G71gat), .B(G78gat), .Z(new_n506));
  INV_X1    g305(.A(KEYINPUT9), .ZN(new_n507));
  XNOR2_X1  g306(.A(G57gat), .B(G64gat), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  XOR2_X1   g308(.A(G57gat), .B(G64gat), .Z(new_n510));
  AOI21_X1  g309(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT93), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G71gat), .B(G78gat), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n515), .B1(new_n512), .B2(new_n511), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n509), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT102), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G85gat), .A2(G92gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n521));
  XOR2_X1   g320(.A(new_n520), .B(new_n521), .Z(new_n522));
  XOR2_X1   g321(.A(KEYINPUT97), .B(G92gat), .Z(new_n523));
  INV_X1    g322(.A(G85gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  XOR2_X1   g324(.A(G99gat), .B(G106gat), .Z(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(G99gat), .ZN(new_n528));
  INV_X1    g327(.A(G106gat), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT8), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n522), .A2(new_n525), .A3(new_n527), .A4(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(KEYINPUT97), .B(G92gat), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n530), .B1(new_n532), .B2(G85gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n520), .B(new_n521), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n526), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n509), .B(KEYINPUT102), .C1(new_n516), .C2(new_n514), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n519), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G230gat), .A2(G233gat), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n517), .A2(new_n531), .A3(new_n518), .A4(new_n535), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n538), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT103), .B(KEYINPUT10), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n543), .B1(new_n538), .B2(new_n541), .ZN(new_n544));
  INV_X1    g343(.A(new_n536), .ZN(new_n545));
  INV_X1    g344(.A(new_n517), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n545), .A2(KEYINPUT10), .A3(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n542), .B1(new_n548), .B2(new_n540), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT107), .ZN(new_n550));
  XOR2_X1   g349(.A(KEYINPUT106), .B(G148gat), .Z(new_n551));
  XNOR2_X1  g350(.A(G176gat), .B(G204gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(KEYINPUT105), .B(G120gat), .Z(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n549), .A2(new_n550), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n550), .B1(new_n549), .B2(new_n555), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n548), .A2(KEYINPUT104), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT104), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n560), .B1(new_n544), .B2(new_n547), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n540), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n542), .ZN(new_n563));
  NOR3_X1   g362(.A1(new_n562), .A2(new_n555), .A3(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n558), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(G15gat), .B(G22gat), .Z(new_n567));
  INV_X1    g366(.A(G1gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT92), .ZN(new_n570));
  AOI21_X1  g369(.A(G8gat), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT16), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(G1gat), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n569), .B1(new_n573), .B2(new_n567), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n571), .B(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT14), .ZN(new_n577));
  OR3_X1    g376(.A1(new_n577), .A2(G29gat), .A3(G36gat), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n577), .B1(G29gat), .B2(G36gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(KEYINPUT91), .B(G36gat), .ZN(new_n580));
  INV_X1    g379(.A(G29gat), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n578), .B(new_n579), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G43gat), .B(G50gat), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n583), .A2(KEYINPUT90), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(KEYINPUT90), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n584), .A2(KEYINPUT15), .A3(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n583), .A2(KEYINPUT15), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n582), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n586), .A2(new_n582), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n576), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n591), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT17), .B1(new_n593), .B2(new_n589), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT17), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT90), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n583), .B(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n587), .B1(new_n597), .B2(KEYINPUT15), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n595), .B(new_n591), .C1(new_n598), .C2(new_n582), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n594), .A2(new_n599), .A3(new_n575), .ZN(new_n600));
  NAND2_X1  g399(.A1(G229gat), .A2(G233gat), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n592), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT18), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n575), .B1(new_n589), .B2(new_n593), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n592), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n601), .B(KEYINPUT13), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n592), .A2(new_n600), .A3(KEYINPUT18), .A4(new_n601), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n604), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT11), .B(G169gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(G197gat), .ZN(new_n613));
  XOR2_X1   g412(.A(G113gat), .B(G141gat), .Z(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n604), .A2(new_n609), .A3(new_n616), .A4(new_n610), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n566), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  OR3_X1    g422(.A1(new_n575), .A2(KEYINPUT21), .A3(new_n546), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n546), .A2(KEYINPUT21), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n546), .A2(KEYINPUT21), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n625), .A2(new_n575), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G127gat), .B(G155gat), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n629), .B(KEYINPUT94), .Z(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n624), .A2(new_n627), .A3(new_n630), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G231gat), .A2(G233gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(new_n283), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(KEYINPUT95), .B(G183gat), .Z(new_n638));
  XOR2_X1   g437(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n636), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n632), .A2(new_n633), .A3(new_n641), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n637), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n640), .B1(new_n637), .B2(new_n642), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n536), .B(KEYINPUT98), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n648), .A2(new_n594), .A3(new_n599), .ZN(new_n649));
  XNOR2_X1  g448(.A(G190gat), .B(G218gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT99), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(KEYINPUT100), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n590), .A2(new_n545), .A3(new_n591), .ZN(new_n653));
  AND2_X1   g452(.A1(G232gat), .A2(G233gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(KEYINPUT41), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n649), .A2(new_n652), .A3(new_n653), .A4(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n651), .A2(KEYINPUT100), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n647), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n649), .A2(new_n655), .ZN(new_n661));
  INV_X1    g460(.A(new_n657), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n661), .A2(new_n662), .A3(new_n652), .A4(new_n653), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n656), .A2(new_n657), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(new_n664), .A3(KEYINPUT101), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n654), .A2(KEYINPUT41), .ZN(new_n666));
  XNOR2_X1  g465(.A(G134gat), .B(G162gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n660), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n668), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n647), .B(new_n670), .C1(new_n658), .C2(new_n659), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n623), .A2(new_n646), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n505), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(new_n274), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(new_n568), .ZN(G1324gat));
  INV_X1    g476(.A(new_n476), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n680));
  INV_X1    g479(.A(G8gat), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n572), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n679), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT42), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(new_n681), .B2(new_n679), .ZN(G1325gat));
  INV_X1    g484(.A(new_n675), .ZN(new_n686));
  AOI21_X1  g485(.A(G15gat), .B1(new_n686), .B2(new_n463), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n500), .A2(new_n502), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n675), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n687), .B1(G15gat), .B2(new_n689), .ZN(G1326gat));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n333), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT43), .B(G22gat), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  AOI21_X1  g492(.A(new_n672), .B1(new_n465), .B2(new_n504), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n623), .A2(new_n645), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n274), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n696), .A2(new_n581), .A3(new_n697), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n698), .A2(KEYINPUT108), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(KEYINPUT108), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT45), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n694), .B(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n705), .A2(new_n697), .A3(new_n695), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(G29gat), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n699), .A2(KEYINPUT45), .A3(new_n700), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n703), .A2(new_n707), .A3(new_n708), .ZN(G1328gat));
  NAND3_X1  g508(.A1(new_n696), .A2(new_n476), .A3(new_n580), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(KEYINPUT46), .Z(new_n711));
  NAND3_X1  g510(.A1(new_n705), .A2(new_n476), .A3(new_n695), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT109), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n711), .B1(new_n714), .B2(new_n580), .ZN(G1329gat));
  INV_X1    g514(.A(new_n688), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n705), .A2(new_n716), .A3(new_n695), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G43gat), .ZN(new_n718));
  INV_X1    g517(.A(G43gat), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n696), .A2(new_n719), .A3(new_n463), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT110), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT47), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n718), .B(new_n720), .C1(new_n722), .C2(KEYINPUT47), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(G1330gat));
  INV_X1    g525(.A(G50gat), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n331), .B1(new_n277), .B2(new_n328), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n696), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n694), .A2(new_n704), .ZN(new_n730));
  AOI211_X1 g529(.A(KEYINPUT44), .B(new_n672), .C1(new_n465), .C2(new_n504), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n728), .B(new_n695), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT112), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(G50gat), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n732), .A2(new_n733), .ZN(new_n736));
  OAI211_X1 g535(.A(KEYINPUT48), .B(new_n729), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n732), .A2(G50gat), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT48), .B1(new_n738), .B2(new_n729), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI211_X1 g540(.A(KEYINPUT111), .B(KEYINPUT48), .C1(new_n738), .C2(new_n729), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n737), .B1(new_n741), .B2(new_n742), .ZN(G1331gat));
  INV_X1    g542(.A(KEYINPUT114), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n645), .A2(new_n566), .A3(new_n672), .A4(new_n621), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT113), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n744), .B1(new_n505), .B2(new_n747), .ZN(new_n748));
  AOI211_X1 g547(.A(KEYINPUT114), .B(new_n746), .C1(new_n465), .C2(new_n504), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n697), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(G57gat), .ZN(G1332gat));
  INV_X1    g551(.A(new_n750), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n678), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n754), .B(KEYINPUT115), .Z(new_n755));
  NOR2_X1   g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1333gat));
  AND3_X1   g557(.A1(new_n441), .A2(KEYINPUT89), .A3(KEYINPUT35), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT89), .B1(new_n441), .B2(KEYINPUT35), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI22_X1  g560(.A1(new_n761), .A2(new_n464), .B1(new_n498), .B2(new_n503), .ZN(new_n762));
  OAI21_X1  g561(.A(KEYINPUT114), .B1(new_n762), .B2(new_n746), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n505), .A2(new_n744), .A3(new_n747), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n763), .A2(new_n463), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT116), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT116), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n763), .A2(new_n767), .A3(new_n463), .A4(new_n764), .ZN(new_n768));
  AOI21_X1  g567(.A(G71gat), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(G71gat), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n750), .B2(new_n716), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT50), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n767), .B1(new_n750), .B2(new_n463), .ZN(new_n773));
  INV_X1    g572(.A(new_n463), .ZN(new_n774));
  NOR4_X1   g573(.A1(new_n748), .A2(new_n749), .A3(KEYINPUT116), .A4(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n770), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n777));
  INV_X1    g576(.A(new_n771), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n772), .A2(new_n779), .ZN(G1334gat));
  NAND2_X1  g579(.A1(new_n750), .A2(new_n728), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g581(.A1(new_n645), .A2(new_n620), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n566), .B(new_n783), .C1(new_n730), .C2(new_n731), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n784), .A2(new_n524), .A3(new_n274), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT117), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n786), .B1(new_n762), .B2(new_n672), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n694), .A2(KEYINPUT117), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n787), .A2(new_n788), .A3(new_n783), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT51), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n787), .A2(new_n791), .A3(new_n788), .A4(new_n783), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n790), .A2(new_n792), .A3(new_n697), .A4(new_n566), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n785), .B1(new_n793), .B2(new_n524), .ZN(G1336gat));
  NOR2_X1   g593(.A1(new_n678), .A2(G92gat), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n790), .A2(new_n792), .A3(new_n566), .A4(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n532), .B1(new_n784), .B2(new_n678), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT52), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n796), .A2(new_n800), .A3(new_n797), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(G1337gat));
  OAI21_X1  g601(.A(G99gat), .B1(new_n784), .B2(new_n688), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n790), .A2(new_n792), .A3(new_n528), .A4(new_n566), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n804), .B2(new_n774), .ZN(G1338gat));
  NOR2_X1   g604(.A1(new_n333), .A2(G106gat), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n790), .A2(new_n792), .A3(new_n566), .A4(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(G106gat), .B1(new_n784), .B2(new_n333), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT53), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n807), .A2(new_n811), .A3(new_n808), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(G1339gat));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n814), .B(new_n539), .C1(new_n544), .C2(new_n547), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n815), .A2(new_n555), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n548), .A2(new_n540), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT54), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n816), .B1(new_n562), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n564), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n816), .B(KEYINPUT55), .C1(new_n562), .C2(new_n818), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n821), .A2(new_n822), .A3(new_n620), .A4(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n606), .A2(new_n608), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n601), .B1(new_n592), .B2(new_n600), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n615), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n619), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n828), .B1(new_n558), .B2(new_n564), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n824), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n672), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n669), .A2(new_n671), .A3(new_n828), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n831), .A2(new_n834), .A3(KEYINPUT119), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT119), .ZN(new_n836));
  AOI22_X1  g635(.A1(new_n824), .A2(new_n829), .B1(new_n669), .B2(new_n671), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n832), .A2(new_n833), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n835), .A2(new_n839), .A3(new_n646), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n645), .A2(new_n672), .A3(new_n621), .A4(new_n565), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(KEYINPUT120), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n840), .A2(new_n846), .A3(new_n843), .ZN(new_n847));
  AND4_X1   g646(.A1(new_n333), .A2(new_n845), .A3(new_n440), .A4(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n476), .A2(new_n274), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n210), .A3(new_n620), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n840), .A2(new_n846), .A3(new_n843), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n846), .B1(new_n840), .B2(new_n843), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n852), .A2(new_n853), .A3(new_n774), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n697), .A3(new_n457), .ZN(new_n855));
  OAI21_X1  g654(.A(G113gat), .B1(new_n855), .B2(new_n621), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n851), .A2(new_n856), .ZN(G1340gat));
  NAND3_X1  g656(.A1(new_n850), .A2(new_n208), .A3(new_n566), .ZN(new_n858));
  OAI21_X1  g657(.A(G120gat), .B1(new_n855), .B2(new_n565), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1341gat));
  NOR3_X1   g659(.A1(new_n855), .A2(new_n207), .A3(new_n646), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n850), .A2(new_n645), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n861), .B1(new_n862), .B2(new_n207), .ZN(G1342gat));
  NAND3_X1  g662(.A1(new_n850), .A2(new_n206), .A3(new_n673), .ZN(new_n864));
  XNOR2_X1  g663(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(G134gat), .B1(new_n855), .B2(new_n672), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n864), .A2(new_n865), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(G1343gat));
  AND2_X1   g668(.A1(new_n688), .A2(new_n849), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n646), .B1(new_n837), .B2(new_n838), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n843), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(KEYINPUT57), .B1(new_n872), .B2(new_n333), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n845), .A2(new_n728), .A3(new_n847), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n870), .B(new_n873), .C1(new_n874), .C2(KEYINPUT57), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n220), .B1(new_n875), .B2(new_n621), .ZN(new_n876));
  INV_X1    g675(.A(new_n874), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n870), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n620), .A2(new_n217), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n876), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT58), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT58), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n876), .B(new_n882), .C1(new_n878), .C2(new_n879), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n883), .ZN(G1344gat));
  NAND4_X1  g683(.A1(new_n877), .A2(new_n221), .A3(new_n566), .A4(new_n870), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n874), .A2(KEYINPUT57), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n870), .B(KEYINPUT122), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n841), .A2(KEYINPUT123), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n841), .A2(KEYINPUT123), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n889), .A2(new_n871), .A3(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n892), .A3(new_n728), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n887), .A2(new_n566), .A3(new_n888), .A4(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n221), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n893), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n897), .B1(new_n874), .B2(KEYINPUT57), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n898), .A2(KEYINPUT124), .A3(new_n566), .A4(new_n888), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n886), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n886), .B1(new_n875), .B2(new_n565), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n901), .A2(new_n221), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n885), .B1(new_n900), .B2(new_n902), .ZN(G1345gat));
  OAI21_X1  g702(.A(new_n225), .B1(new_n878), .B2(new_n646), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n875), .A2(new_n225), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(new_n646), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(G1346gat));
  XOR2_X1   g706(.A(KEYINPUT74), .B(G162gat), .Z(new_n908));
  OAI21_X1  g707(.A(new_n908), .B1(new_n878), .B2(new_n672), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n875), .A2(new_n908), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(new_n672), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(G1347gat));
  INV_X1    g711(.A(G169gat), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n678), .A2(new_n697), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n848), .A2(new_n913), .A3(new_n620), .A4(new_n914), .ZN(new_n915));
  NOR4_X1   g714(.A1(new_n852), .A2(new_n853), .A3(new_n728), .A4(new_n774), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(new_n914), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n917), .A2(new_n621), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n915), .B1(new_n919), .B2(new_n913), .ZN(G1348gat));
  INV_X1    g719(.A(G176gat), .ZN(new_n921));
  NOR4_X1   g720(.A1(new_n917), .A2(new_n921), .A3(new_n565), .A4(new_n918), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n848), .A2(new_n914), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n921), .B1(new_n923), .B2(new_n565), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n922), .B1(new_n926), .B2(new_n927), .ZN(G1349gat));
  NAND4_X1  g727(.A1(new_n854), .A2(new_n333), .A3(new_n645), .A4(new_n914), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(KEYINPUT126), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT126), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n916), .A2(new_n931), .A3(new_n645), .A4(new_n914), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n930), .A2(G183gat), .A3(new_n932), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n848), .A2(new_n334), .A3(new_n645), .A4(new_n914), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT60), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT60), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n933), .A2(new_n937), .A3(new_n934), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1350gat));
  NAND3_X1  g738(.A1(new_n916), .A2(new_n673), .A3(new_n914), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT61), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n940), .A2(new_n941), .A3(G190gat), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n941), .B1(new_n940), .B2(G190gat), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n673), .A2(new_n335), .ZN(new_n944));
  OAI22_X1  g743(.A1(new_n942), .A2(new_n943), .B1(new_n923), .B2(new_n944), .ZN(G1351gat));
  NOR3_X1   g744(.A1(new_n874), .A2(new_n716), .A3(new_n918), .ZN(new_n946));
  INV_X1    g745(.A(G197gat), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(new_n947), .A3(new_n620), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n918), .A2(new_n716), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n898), .A2(new_n620), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n948), .B1(new_n950), .B2(new_n947), .ZN(G1352gat));
  INV_X1    g750(.A(G204gat), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n946), .A2(new_n952), .A3(new_n566), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n898), .A2(new_n566), .A3(new_n949), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n954), .B(new_n955), .C1(new_n952), .C2(new_n956), .ZN(G1353gat));
  NAND3_X1  g756(.A1(new_n898), .A2(new_n645), .A3(new_n949), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(G211gat), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n959), .A2(new_n960), .A3(KEYINPUT63), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n946), .A2(new_n283), .A3(new_n645), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(KEYINPUT63), .ZN(new_n963));
  OR2_X1    g762(.A1(new_n960), .A2(KEYINPUT63), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n958), .A2(G211gat), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n961), .A2(new_n962), .A3(new_n965), .ZN(G1354gat));
  NAND3_X1  g765(.A1(new_n946), .A2(new_n284), .A3(new_n673), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n898), .A2(new_n673), .A3(new_n949), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n967), .B1(new_n968), .B2(new_n284), .ZN(G1355gat));
endmodule


