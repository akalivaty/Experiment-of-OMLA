//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1233, new_n1234, new_n1235, new_n1236, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n208), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT64), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n219), .A2(KEYINPUT65), .A3(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G226), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n201), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  INV_X1    g0024(.A(G77), .ZN(new_n225));
  INV_X1    g0025(.A(G244), .ZN(new_n226));
  OAI22_X1  g0026(.A1(new_n203), .A2(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n223), .B(new_n227), .C1(G116), .C2(G270), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n221), .A2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(KEYINPUT65), .B1(new_n219), .B2(new_n220), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n210), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n213), .B1(new_n216), .B2(new_n217), .C1(new_n231), .C2(KEYINPUT1), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G226), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  AND2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  OAI211_X1 g0051(.A(new_n208), .B(G87), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT83), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n259), .A2(KEYINPUT83), .A3(new_n208), .A4(G87), .ZN(new_n260));
  AND3_X1   g0060(.A1(new_n254), .A2(new_n260), .A3(KEYINPUT22), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT22), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n252), .A2(new_n253), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT84), .ZN(new_n264));
  INV_X1    g0064(.A(G107), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G20), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n264), .B1(new_n266), .B2(KEYINPUT23), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT23), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(new_n265), .A3(G20), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n208), .A2(G33), .A3(G116), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n266), .A2(new_n264), .A3(KEYINPUT23), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n263), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(KEYINPUT24), .B1(new_n261), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n254), .A2(new_n260), .A3(KEYINPUT22), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT24), .ZN(new_n277));
  INV_X1    g0077(.A(new_n273), .ZN(new_n278));
  NOR3_X1   g0078(.A1(new_n278), .A2(new_n267), .A3(new_n271), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n276), .A2(new_n277), .A3(new_n279), .A4(new_n263), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n214), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n265), .ZN(new_n287));
  XNOR2_X1  g0087(.A(new_n287), .B(KEYINPUT25), .ZN(new_n288));
  INV_X1    g0088(.A(new_n283), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n207), .A2(KEYINPUT72), .A3(G33), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT72), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(new_n256), .B2(G1), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n289), .A2(new_n290), .A3(new_n285), .A4(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(new_n265), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n288), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G1698), .ZN(new_n296));
  OAI211_X1 g0096(.A(G250), .B(new_n296), .C1(new_n250), .C2(new_n251), .ZN(new_n297));
  OAI211_X1 g0097(.A(G257), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G294), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G41), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n207), .B(G45), .C1(new_n303), .C2(KEYINPUT5), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT5), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n306), .A2(G41), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n301), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G264), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT73), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(new_n306), .B2(G41), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n303), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G274), .ZN(new_n315));
  AND2_X1   g0115(.A1(G1), .A2(G13), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G41), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n305), .A2(new_n314), .A3(new_n318), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n302), .A2(new_n310), .A3(G179), .A4(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT85), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n302), .A2(new_n310), .A3(new_n319), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n320), .A2(new_n321), .B1(new_n323), .B2(G169), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n284), .A2(new_n295), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n301), .A2(new_n300), .B1(new_n309), .B2(G264), .ZN(new_n326));
  AOI21_X1  g0126(.A(G200), .B1(new_n326), .B2(new_n319), .ZN(new_n327));
  INV_X1    g0127(.A(G190), .ZN(new_n328));
  AND4_X1   g0128(.A1(new_n328), .A2(new_n302), .A3(new_n310), .A4(new_n319), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n289), .B1(new_n275), .B2(new_n280), .ZN(new_n331));
  INV_X1    g0131(.A(new_n295), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(KEYINPUT86), .B1(new_n325), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n324), .A2(new_n322), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n331), .B2(new_n332), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n284), .B(new_n295), .C1(new_n329), .C2(new_n327), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT86), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n285), .A2(G50), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n283), .B1(new_n207), .B2(G20), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n341), .B1(new_n342), .B2(G50), .ZN(new_n343));
  NOR2_X1   g0143(.A1(G20), .A2(G33), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G150), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT8), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G58), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n208), .A2(G33), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI211_X1 g0153(.A(new_n347), .B(new_n353), .C1(G20), .C2(new_n204), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n343), .B1(new_n354), .B2(new_n289), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n296), .A2(G222), .ZN(new_n356));
  INV_X1    g0156(.A(G223), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n259), .B(new_n356), .C1(new_n357), .C2(new_n296), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n358), .B(new_n301), .C1(G77), .C2(new_n259), .ZN(new_n359));
  INV_X1    g0159(.A(G45), .ZN(new_n360));
  AOI21_X1  g0160(.A(G1), .B1(new_n303), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n317), .A2(G1), .A3(G13), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(new_n362), .A3(G274), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n301), .A2(new_n361), .ZN(new_n364));
  XOR2_X1   g0164(.A(KEYINPUT66), .B(G226), .Z(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n359), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  OR2_X1    g0167(.A1(new_n367), .A2(KEYINPUT67), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(KEYINPUT67), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n355), .B1(new_n370), .B2(G169), .ZN(new_n371));
  AOI21_X1  g0171(.A(G179), .B1(new_n368), .B2(new_n369), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n370), .A2(G190), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n355), .A2(KEYINPUT9), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT9), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n376), .B(new_n343), .C1(new_n354), .C2(new_n289), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n368), .A2(G200), .A3(new_n369), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n374), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT10), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT10), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n374), .A2(new_n378), .A3(new_n382), .A4(new_n379), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n373), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT16), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n257), .A2(new_n208), .A3(new_n258), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT7), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n257), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n258), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n203), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n202), .A2(new_n203), .ZN(new_n392));
  NOR2_X1   g0192(.A1(G58), .A2(G68), .ZN(new_n393));
  OAI21_X1  g0193(.A(G20), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n344), .A2(G159), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n386), .B1(new_n391), .B2(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n250), .A2(new_n251), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT7), .B1(new_n398), .B2(new_n208), .ZN(new_n399));
  INV_X1    g0199(.A(new_n390), .ZN(new_n400));
  OAI21_X1  g0200(.A(G68), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n396), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(KEYINPUT16), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n397), .A2(new_n403), .A3(new_n283), .ZN(new_n404));
  INV_X1    g0204(.A(new_n351), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n405), .A2(new_n285), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n406), .B1(new_n342), .B2(new_n405), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT18), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n357), .A2(new_n296), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n222), .A2(G1698), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n410), .B(new_n411), .C1(new_n250), .C2(new_n251), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G87), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n362), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n362), .A2(G232), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n363), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G169), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(G179), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n408), .A2(new_n409), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n409), .B1(new_n408), .B2(new_n422), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n328), .A2(KEYINPUT70), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n328), .A2(KEYINPUT70), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(KEYINPUT71), .B1(new_n419), .B2(new_n429), .ZN(new_n430));
  NOR4_X1   g0230(.A1(new_n414), .A2(new_n417), .A3(KEYINPUT71), .A4(new_n429), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(G200), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n419), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n430), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT17), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n435), .A2(new_n436), .A3(new_n404), .A4(new_n407), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n414), .A2(new_n417), .A3(new_n429), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT71), .ZN(new_n439));
  OAI22_X1  g0239(.A1(new_n438), .A2(new_n439), .B1(G200), .B2(new_n418), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n404), .B(new_n407), .C1(new_n440), .C2(new_n431), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT17), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n425), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n203), .A2(G20), .ZN(new_n445));
  OAI221_X1 g0245(.A(new_n445), .B1(new_n352), .B2(new_n225), .C1(new_n345), .C2(new_n201), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n446), .A2(new_n283), .ZN(new_n447));
  OR2_X1    g0247(.A1(new_n447), .A2(KEYINPUT11), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(KEYINPUT11), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT12), .ZN(new_n450));
  INV_X1    g0250(.A(G13), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n450), .A2(new_n451), .A3(G1), .ZN(new_n452));
  INV_X1    g0252(.A(new_n445), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n452), .A2(new_n453), .B1(new_n450), .B2(new_n285), .ZN(new_n454));
  OAI21_X1  g0254(.A(G68), .B1(new_n342), .B2(new_n450), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n448), .A2(new_n449), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n296), .A2(G226), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT68), .B1(new_n398), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT68), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n259), .A2(new_n459), .A3(G226), .A4(new_n296), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  OAI211_X1 g0261(.A(G232), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G97), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n362), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n364), .A2(G238), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n363), .ZN(new_n468));
  OAI21_X1  g0268(.A(KEYINPUT13), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n467), .A2(new_n363), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT13), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n464), .B1(new_n460), .B2(new_n458), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n470), .B(new_n471), .C1(new_n472), .C2(new_n362), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT14), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n474), .A2(new_n475), .A3(G169), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n469), .A2(new_n473), .A3(G179), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n475), .B1(new_n474), .B2(G169), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n456), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n469), .A2(new_n473), .A3(G190), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT69), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT69), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n469), .A2(new_n473), .A3(new_n483), .A4(G190), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n456), .B1(G200), .B2(new_n474), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n480), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G238), .A2(G1698), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n259), .B(new_n489), .C1(new_n237), .C2(G1698), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n490), .B(new_n301), .C1(G107), .C2(new_n259), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n364), .A2(G244), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(new_n363), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G200), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n342), .A2(G77), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(G77), .B2(new_n285), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G20), .A2(G77), .ZN(new_n497));
  XNOR2_X1  g0297(.A(KEYINPUT15), .B(G87), .ZN(new_n498));
  OAI221_X1 g0298(.A(new_n497), .B1(new_n498), .B2(new_n352), .C1(new_n351), .C2(new_n345), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n496), .B1(new_n283), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n494), .B(new_n500), .C1(new_n328), .C2(new_n493), .ZN(new_n501));
  INV_X1    g0301(.A(G169), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n493), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n499), .A2(new_n283), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n504), .B(new_n495), .C1(G77), .C2(new_n285), .ZN(new_n505));
  INV_X1    g0305(.A(G179), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n491), .A2(new_n506), .A3(new_n363), .A4(new_n492), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n503), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n501), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NOR4_X1   g0310(.A1(new_n385), .A2(new_n444), .A3(new_n488), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G283), .ZN(new_n512));
  INV_X1    g0312(.A(G97), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n512), .B(new_n208), .C1(G33), .C2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(G116), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G20), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n283), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT81), .ZN(new_n518));
  OR2_X1    g0318(.A1(new_n518), .A2(KEYINPUT20), .ZN(new_n519));
  OR2_X1    g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n292), .A2(new_n290), .A3(new_n285), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n521), .A2(new_n283), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G116), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n286), .A2(new_n515), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n518), .A2(KEYINPUT20), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n517), .A2(new_n519), .A3(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n520), .A2(new_n523), .A3(new_n524), .A4(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(G303), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n257), .A2(new_n528), .A3(new_n258), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G264), .A2(G1698), .ZN(new_n530));
  INV_X1    g0330(.A(G257), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n530), .B1(new_n531), .B2(G1698), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n529), .B(new_n301), .C1(new_n398), .C2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n319), .ZN(new_n534));
  OAI211_X1 g0334(.A(G270), .B(new_n362), .C1(new_n304), .C2(new_n307), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT80), .ZN(new_n536));
  OR2_X1    g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n536), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n534), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n527), .B1(new_n539), .B2(new_n429), .ZN(new_n540));
  XNOR2_X1  g0340(.A(new_n535), .B(new_n536), .ZN(new_n541));
  INV_X1    g0341(.A(new_n534), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G200), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(G169), .A3(new_n527), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT21), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n541), .A2(G179), .A3(new_n542), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n527), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n543), .A2(KEYINPUT21), .A3(G169), .A4(new_n527), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n545), .A2(new_n548), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT82), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n550), .A2(new_n551), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT82), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n554), .A2(new_n555), .A3(new_n548), .A4(new_n545), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT6), .ZN(new_n558));
  NOR3_X1   g0358(.A1(new_n558), .A2(new_n513), .A3(G107), .ZN(new_n559));
  XNOR2_X1  g0359(.A(G97), .B(G107), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n559), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  OAI22_X1  g0361(.A1(new_n561), .A2(new_n208), .B1(new_n225), .B2(new_n345), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n265), .B1(new_n389), .B2(new_n390), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n283), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n285), .A2(G97), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n522), .B2(G97), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT4), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n568), .A2(G1698), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n569), .B(G244), .C1(new_n251), .C2(new_n250), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n226), .B1(new_n257), .B2(new_n258), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n570), .B(new_n512), .C1(new_n571), .C2(KEYINPUT4), .ZN(new_n572));
  OAI21_X1  g0372(.A(G250), .B1(new_n250), .B2(new_n251), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n296), .B1(new_n573), .B2(KEYINPUT4), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n301), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(G257), .B(new_n362), .C1(new_n304), .C2(new_n307), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n319), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT74), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n319), .A2(KEYINPUT74), .A3(new_n576), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n575), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n567), .B1(G200), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT75), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n575), .A2(new_n579), .A3(new_n580), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n583), .B1(new_n584), .B2(G190), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n581), .A2(KEYINPUT75), .A3(new_n328), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n582), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  XOR2_X1   g0387(.A(KEYINPUT15), .B(G87), .Z(new_n588));
  INV_X1    g0388(.A(KEYINPUT78), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n498), .A2(KEYINPUT78), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(KEYINPUT79), .B1(new_n592), .B2(new_n293), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT79), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n522), .A2(new_n594), .A3(new_n590), .A4(new_n591), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n588), .A2(new_n285), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n259), .A2(new_n208), .A3(G68), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT19), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n352), .B2(new_n513), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n208), .B1(new_n463), .B2(new_n599), .ZN(new_n601));
  INV_X1    g0401(.A(G87), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(new_n513), .A3(new_n265), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n601), .A2(KEYINPUT77), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT77), .B1(new_n601), .B2(new_n603), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n598), .B(new_n600), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n597), .B1(new_n606), .B2(new_n283), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n596), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n224), .A2(new_n296), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n226), .A2(G1698), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n609), .B(new_n610), .C1(new_n250), .C2(new_n251), .ZN(new_n611));
  NAND2_X1  g0411(.A1(G33), .A2(G116), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(KEYINPUT76), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT76), .B1(new_n611), .B2(new_n612), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n614), .A2(new_n615), .A3(new_n362), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n207), .A2(G45), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n617), .A2(G274), .ZN(new_n618));
  AOI21_X1  g0418(.A(G250), .B1(new_n207), .B2(G45), .ZN(new_n619));
  NOR3_X1   g0419(.A1(new_n618), .A2(new_n301), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n502), .B1(new_n616), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n611), .A2(new_n612), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT76), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n362), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n620), .B1(new_n624), .B2(new_n613), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n506), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n608), .A2(new_n621), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(G200), .B1(new_n616), .B2(new_n620), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n521), .A2(new_n602), .A3(new_n283), .ZN(new_n629));
  AOI211_X1 g0429(.A(new_n597), .B(new_n629), .C1(new_n606), .C2(new_n283), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n625), .A2(G190), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n628), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n581), .A2(new_n502), .B1(new_n564), .B2(new_n566), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n584), .A2(new_n506), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n587), .A2(new_n633), .A3(new_n636), .ZN(new_n637));
  AND4_X1   g0437(.A1(new_n340), .A2(new_n511), .A3(new_n557), .A4(new_n637), .ZN(G372));
  INV_X1    g0438(.A(new_n508), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n487), .A2(new_n639), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n640), .A2(new_n480), .B1(new_n442), .B2(new_n437), .ZN(new_n641));
  INV_X1    g0441(.A(new_n425), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n381), .A2(new_n383), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n373), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n511), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT87), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n627), .A2(new_n632), .A3(new_n635), .A4(new_n634), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT26), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n648), .A2(new_n647), .A3(new_n649), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n554), .A2(new_n548), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(new_n325), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n587), .A2(new_n633), .A3(new_n337), .A4(new_n636), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n627), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n645), .B1(new_n646), .B2(new_n659), .ZN(G369));
  INV_X1    g0460(.A(KEYINPUT89), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n662));
  AOI21_X1  g0462(.A(KEYINPUT88), .B1(new_n662), .B2(KEYINPUT27), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n662), .A2(KEYINPUT88), .A3(KEYINPUT27), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(G213), .B1(new_n662), .B2(KEYINPUT27), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(G343), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n527), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(new_n554), .B2(new_n548), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n672), .B1(new_n557), .B2(new_n671), .ZN(new_n673));
  INV_X1    g0473(.A(G330), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n661), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n553), .A2(new_n556), .B1(new_n527), .B2(new_n670), .ZN(new_n676));
  OAI211_X1 g0476(.A(KEYINPUT89), .B(G330), .C1(new_n676), .C2(new_n672), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n670), .B1(new_n331), .B2(new_n332), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n340), .A2(new_n679), .B1(new_n325), .B2(new_n670), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n340), .A2(new_n655), .A3(new_n669), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n325), .A2(new_n669), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n682), .A2(new_n686), .ZN(G399));
  INV_X1    g0487(.A(new_n211), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G41), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(new_n207), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n603), .A2(G116), .ZN(new_n691));
  INV_X1    g0491(.A(new_n217), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n690), .A2(new_n691), .B1(new_n692), .B2(new_n689), .ZN(new_n693));
  XOR2_X1   g0493(.A(new_n693), .B(KEYINPUT28), .Z(new_n694));
  XNOR2_X1  g0494(.A(KEYINPUT90), .B(KEYINPUT31), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT30), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n539), .A2(new_n625), .A3(G179), .A4(new_n326), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n696), .B1(new_n697), .B2(new_n581), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n625), .A2(new_n326), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n699), .A2(KEYINPUT30), .A3(new_n549), .A4(new_n584), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n539), .A2(G179), .ZN(new_n701));
  INV_X1    g0501(.A(new_n625), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n701), .A2(new_n323), .A3(new_n581), .A4(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n698), .A2(new_n700), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n670), .ZN(new_n705));
  MUX2_X1   g0505(.A(new_n695), .B(KEYINPUT31), .S(new_n705), .Z(new_n706));
  NAND4_X1  g0506(.A1(new_n340), .A2(new_n557), .A3(new_n637), .A4(new_n669), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n674), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n669), .B1(new_n654), .B2(new_n658), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n648), .B(KEYINPUT26), .ZN(new_n712));
  OAI211_X1 g0512(.A(KEYINPUT29), .B(new_n669), .C1(new_n658), .C2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n708), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n694), .B1(new_n714), .B2(G1), .ZN(G364));
  NAND2_X1  g0515(.A1(new_n208), .A2(G13), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT91), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G45), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n690), .A2(new_n718), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n676), .A2(G330), .A3(new_n672), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n719), .B1(new_n678), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n208), .A2(new_n506), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G200), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n428), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n723), .A2(G190), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI22_X1  g0527(.A1(new_n725), .A2(new_n201), .B1(new_n727), .B2(new_n203), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n208), .A2(G190), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(new_n506), .A3(G200), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n730), .A2(KEYINPUT94), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(KEYINPUT94), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G107), .ZN(new_n735));
  NOR4_X1   g0535(.A1(new_n208), .A2(new_n328), .A3(new_n433), .A4(G179), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n398), .B1(new_n736), .B2(G87), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n722), .A2(new_n433), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n428), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n735), .B(new_n737), .C1(new_n202), .C2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n738), .A2(G190), .ZN(new_n742));
  AOI211_X1 g0542(.A(new_n728), .B(new_n741), .C1(G77), .C2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n506), .A2(new_n433), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT93), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n208), .B1(new_n746), .B2(G190), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n743), .B1(new_n513), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n746), .A2(new_n729), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G159), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT32), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(G329), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n734), .A2(G283), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n742), .A2(G311), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n259), .B1(new_n736), .B2(G303), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n753), .A2(new_n754), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  AOI22_X1  g0557(.A1(G322), .A2(new_n739), .B1(new_n724), .B2(G326), .ZN(new_n758));
  INV_X1    g0558(.A(G317), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(KEYINPUT33), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n759), .A2(KEYINPUT33), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n726), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G294), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n758), .B(new_n762), .C1(new_n747), .C2(new_n763), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n748), .A2(new_n752), .B1(new_n757), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n214), .B1(G20), .B2(new_n502), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n211), .A2(new_n398), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(new_n360), .B2(new_n692), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(new_n245), .B2(new_n360), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n688), .A2(new_n398), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n770), .A2(G355), .B1(new_n515), .B2(new_n688), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n772), .A2(KEYINPUT92), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G13), .A2(G33), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G20), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n766), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n778), .B1(new_n772), .B2(KEYINPUT92), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n765), .A2(new_n766), .B1(new_n773), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n673), .A2(new_n776), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n719), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n721), .A2(new_n783), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n784), .A2(KEYINPUT95), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(KEYINPUT95), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(new_n786), .ZN(G396));
  NAND2_X1  g0587(.A1(new_n670), .A2(new_n505), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n509), .A2(KEYINPUT97), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n501), .A2(new_n788), .A3(new_n508), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT97), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n508), .A2(new_n669), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n793), .A2(KEYINPUT98), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(KEYINPUT98), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n789), .A2(new_n792), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n709), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n796), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n669), .B(new_n798), .C1(new_n654), .C2(new_n658), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n797), .A2(new_n708), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n719), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(KEYINPUT99), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT99), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(new_n800), .B2(new_n719), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n708), .B1(new_n797), .B2(new_n799), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n802), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n719), .ZN(new_n807));
  INV_X1    g0607(.A(new_n766), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n775), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n807), .B1(G77), .B2(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT96), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n724), .A2(G137), .B1(new_n742), .B2(G159), .ZN(new_n812));
  INV_X1    g0612(.A(G143), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n812), .B1(new_n813), .B2(new_n740), .C1(new_n346), .C2(new_n727), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT34), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n734), .A2(G68), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n398), .B1(new_n736), .B2(G50), .ZN(new_n817));
  INV_X1    g0617(.A(G132), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n816), .B(new_n817), .C1(new_n818), .C2(new_n749), .ZN(new_n819));
  INV_X1    g0619(.A(new_n747), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n819), .B1(G58), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n733), .A2(new_n602), .ZN(new_n822));
  INV_X1    g0622(.A(new_n736), .ZN(new_n823));
  INV_X1    g0623(.A(new_n742), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n398), .B1(new_n823), .B2(new_n265), .C1(new_n824), .C2(new_n515), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n822), .B(new_n825), .C1(G311), .C2(new_n750), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n739), .A2(G294), .B1(new_n726), .B2(G283), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n528), .B2(new_n725), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(G97), .B2(new_n820), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n815), .A2(new_n821), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n811), .B1(new_n808), .B2(new_n830), .C1(new_n798), .C2(new_n775), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(KEYINPUT100), .B1(new_n806), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT100), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n804), .A2(new_n805), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n834), .B(new_n831), .C1(new_n835), .C2(new_n802), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n833), .A2(new_n836), .ZN(G384));
  NOR2_X1   g0637(.A1(new_n717), .A2(new_n207), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT40), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n704), .A2(KEYINPUT31), .A3(new_n670), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT106), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n705), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n704), .A2(KEYINPUT106), .A3(new_n670), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n842), .A2(new_n695), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n707), .A2(new_n840), .A3(new_n844), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n485), .A2(new_n486), .ZN(new_n846));
  INV_X1    g0646(.A(new_n479), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n847), .A2(new_n477), .A3(new_n476), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n456), .B(new_n670), .C1(new_n846), .C2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n456), .A2(new_n670), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n480), .A2(new_n487), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n796), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT38), .ZN(new_n853));
  INV_X1    g0653(.A(new_n407), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT103), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n391), .B2(new_n396), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n401), .A2(KEYINPUT103), .A3(new_n402), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n856), .A2(new_n857), .A3(new_n386), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n391), .A2(new_n396), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n289), .B1(new_n859), .B2(KEYINPUT16), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n854), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n668), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(new_n425), .B2(new_n443), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT37), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n408), .A2(new_n422), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n408), .A2(new_n668), .ZN(new_n868));
  AND4_X1   g0668(.A1(new_n866), .A2(new_n867), .A3(new_n868), .A4(new_n441), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n441), .B1(new_n861), .B2(new_n862), .ZN(new_n870));
  INV_X1    g0670(.A(new_n422), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n861), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT37), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n869), .B1(new_n873), .B2(KEYINPUT104), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT104), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n875), .B(KEYINPUT37), .C1(new_n870), .C2(new_n872), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n853), .B(new_n865), .C1(new_n874), .C2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n873), .A2(KEYINPUT104), .ZN(new_n878));
  INV_X1    g0678(.A(new_n869), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n878), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n865), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT38), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n845), .B(new_n852), .C1(new_n877), .C2(new_n882), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n845), .A2(new_n852), .A3(KEYINPUT40), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n880), .A2(KEYINPUT38), .A3(new_n881), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n867), .A2(new_n868), .A3(new_n441), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n886), .B(new_n866), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n868), .B1(new_n425), .B2(new_n443), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n853), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n839), .A2(new_n883), .B1(new_n884), .B2(new_n890), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n511), .A2(new_n845), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n674), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n892), .B2(new_n891), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT107), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n880), .A2(new_n881), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n853), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n897), .B1(new_n899), .B2(new_n885), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n885), .A2(new_n897), .A3(new_n889), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT105), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n848), .A2(new_n456), .A3(new_n669), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT39), .B1(new_n877), .B2(new_n882), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT105), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n885), .A2(new_n897), .A3(new_n889), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n902), .A2(new_n904), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n849), .A2(new_n851), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n508), .A2(new_n670), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n911), .B1(new_n799), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n899), .A2(new_n885), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n914), .A2(new_n915), .B1(new_n642), .B2(new_n862), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n909), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n711), .A2(new_n511), .A3(new_n713), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n645), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n917), .B(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n838), .B1(new_n896), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n896), .B2(new_n920), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n561), .B(KEYINPUT101), .Z(new_n923));
  NOR2_X1   g0723(.A1(new_n923), .A2(KEYINPUT35), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n924), .A2(new_n515), .A3(new_n216), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n926), .A2(KEYINPUT102), .B1(KEYINPUT35), .B2(new_n923), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(KEYINPUT102), .B2(new_n926), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT36), .ZN(new_n929));
  NOR3_X1   g0729(.A1(new_n392), .A2(new_n217), .A3(new_n225), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n203), .A2(G50), .ZN(new_n931));
  OAI211_X1 g0731(.A(G1), .B(new_n451), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n922), .A2(new_n929), .A3(new_n932), .ZN(G367));
  NAND2_X1  g0733(.A1(new_n670), .A2(new_n567), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n587), .A2(new_n636), .A3(new_n934), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n935), .A2(new_n336), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n670), .B1(new_n936), .B2(new_n636), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n655), .A2(new_n669), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n339), .B2(new_n334), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n634), .A2(new_n635), .A3(new_n670), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n935), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n937), .B1(new_n942), .B2(KEYINPUT42), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n942), .A2(KEYINPUT42), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n630), .A2(new_n669), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n633), .A2(new_n945), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n945), .A2(new_n627), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n943), .A2(new_n944), .B1(KEYINPUT43), .B2(new_n948), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n941), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n682), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n949), .A2(new_n950), .ZN(new_n954));
  AND3_X1   g0754(.A1(new_n951), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n953), .B1(new_n951), .B2(new_n954), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n689), .B(KEYINPUT41), .Z(new_n958));
  INV_X1    g0758(.A(new_n658), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n652), .A2(new_n653), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n670), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n713), .B1(new_n961), .B2(KEYINPUT29), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n939), .B1(new_n680), .B2(new_n938), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n678), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n708), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n340), .A2(new_n679), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n325), .A2(new_n670), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n966), .A2(new_n967), .A3(new_n938), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n683), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n969), .A2(new_n675), .A3(new_n677), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n962), .A2(new_n964), .A3(new_n965), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(KEYINPUT109), .ZN(new_n972));
  XOR2_X1   g0772(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n973));
  NAND3_X1  g0773(.A1(new_n686), .A2(new_n941), .A3(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n973), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n685), .B2(new_n952), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(KEYINPUT44), .B1(new_n686), .B2(new_n941), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT44), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n685), .A2(new_n979), .A3(new_n952), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n977), .A2(new_n682), .A3(new_n978), .A4(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT109), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n714), .A2(new_n982), .A3(new_n964), .A4(new_n970), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n978), .A2(new_n974), .A3(new_n980), .A4(new_n976), .ZN(new_n984));
  INV_X1    g0784(.A(new_n682), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n972), .A2(new_n981), .A3(new_n983), .A4(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n958), .B1(new_n987), .B2(new_n714), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n718), .A2(G1), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n957), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n241), .A2(new_n211), .A3(new_n398), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n778), .B1(new_n688), .B2(new_n588), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n719), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n776), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n725), .A2(new_n813), .B1(new_n824), .B2(new_n201), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(G159), .B2(new_n726), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n747), .A2(new_n203), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n734), .A2(G77), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n398), .B1(new_n739), .B2(G150), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n996), .A2(new_n998), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(G137), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n749), .A2(new_n1002), .B1(new_n202), .B2(new_n823), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT110), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n733), .A2(new_n513), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(G317), .B2(new_n750), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n823), .A2(new_n515), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1007), .A2(KEYINPUT46), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n1007), .A2(KEYINPUT46), .B1(new_n726), .B2(G294), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1006), .A2(new_n398), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n724), .A2(G311), .B1(new_n742), .B2(G283), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n528), .B2(new_n740), .C1(new_n747), .C2(new_n265), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n1001), .A2(new_n1004), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT47), .Z(new_n1014));
  OAI221_X1 g0814(.A(new_n993), .B1(new_n994), .B2(new_n948), .C1(new_n1014), .C2(new_n808), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n990), .A2(new_n1015), .ZN(G387));
  AND2_X1   g0816(.A1(new_n972), .A2(new_n983), .ZN(new_n1017));
  AND2_X1   g0817(.A1(new_n964), .A2(new_n970), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n689), .B1(new_n1018), .B2(new_n714), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1018), .A2(new_n989), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT111), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1018), .A2(KEYINPUT111), .A3(new_n989), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n211), .A2(G107), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n351), .A2(G50), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT50), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n691), .ZN(new_n1030));
  AOI211_X1 g0830(.A(G45), .B(new_n1030), .C1(G68), .C2(G77), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n767), .B(new_n1032), .C1(new_n238), .C2(G45), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1027), .B(new_n1033), .C1(new_n1030), .C2(new_n770), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n807), .B1(new_n1034), .B2(new_n778), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n259), .B1(new_n750), .B2(G326), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n724), .A2(G322), .B1(new_n726), .B2(G311), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n528), .B2(new_n824), .C1(new_n759), .C2(new_n740), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT48), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n820), .A2(G283), .B1(G294), .B2(new_n736), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT49), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1036), .B1(new_n515), .B2(new_n733), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n259), .B1(new_n823), .B2(new_n225), .C1(new_n824), .C2(new_n203), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1048), .A2(new_n1005), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n346), .B2(new_n749), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n747), .A2(new_n592), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n724), .A2(G159), .B1(new_n726), .B2(new_n405), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(new_n201), .C2(new_n740), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n1045), .A2(new_n1047), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1035), .B1(new_n1054), .B2(new_n766), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n680), .A2(new_n776), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n1026), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1021), .A2(new_n1058), .ZN(G393));
  AOI21_X1  g0859(.A(KEYINPUT112), .B1(new_n984), .B2(new_n985), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(new_n981), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n689), .B(new_n987), .C1(new_n1061), .C2(new_n1017), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n777), .B1(new_n513), .B2(new_n211), .C1(new_n248), .C2(new_n767), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n807), .A2(new_n1063), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT113), .Z(new_n1065));
  OAI22_X1  g0865(.A1(new_n727), .A2(new_n528), .B1(new_n824), .B2(new_n763), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G311), .A2(new_n739), .B1(new_n724), .B2(G317), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT52), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1066), .B(new_n1068), .C1(G116), .C2(new_n820), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n750), .A2(G322), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n259), .B1(new_n736), .B2(G283), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1070), .A2(new_n735), .A3(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT114), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G150), .A2(new_n724), .B1(new_n739), .B2(G159), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT51), .Z(new_n1075));
  OAI22_X1  g0875(.A1(new_n749), .A2(new_n813), .B1(new_n733), .B2(new_n602), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n398), .B1(new_n736), .B2(G68), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1077), .B1(new_n824), .B2(new_n351), .C1(new_n201), .C2(new_n727), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1076), .B(new_n1078), .C1(G77), .C2(new_n820), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1069), .A2(new_n1073), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1065), .B1(new_n1080), .B2(new_n808), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n952), .B2(new_n776), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n1061), .B2(new_n989), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1062), .A2(new_n1083), .ZN(G390));
  NAND2_X1  g0884(.A1(new_n845), .A2(G330), .ZN(new_n1085));
  NOR3_X1   g0885(.A1(new_n1085), .A2(new_n796), .A3(new_n911), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n799), .A2(new_n913), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n904), .B1(new_n1087), .B2(new_n910), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n902), .B2(new_n908), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n798), .B(new_n669), .C1(new_n658), .C2(new_n712), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1090), .A2(new_n913), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n890), .B(new_n903), .C1(new_n1091), .C2(new_n911), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1086), .B1(new_n1089), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1087), .A2(new_n910), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n903), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n906), .B1(new_n905), .B2(new_n907), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n708), .A2(new_n910), .A3(new_n798), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1099), .A2(new_n1092), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1094), .A2(new_n1101), .A3(new_n989), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT115), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1094), .A2(new_n1101), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n910), .B1(new_n708), .B2(new_n798), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1087), .B1(new_n1086), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n911), .B1(new_n1085), .B2(new_n796), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1107), .A2(new_n1091), .A3(new_n1100), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n918), .B(new_n645), .C1(new_n646), .C2(new_n1085), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1104), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1110), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1094), .A2(new_n1101), .A3(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1113), .A2(new_n689), .A3(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n774), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n807), .B1(new_n405), .B2(new_n809), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n816), .B1(new_n763), .B2(new_n749), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT116), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n398), .B1(new_n823), .B2(new_n602), .C1(new_n824), .C2(new_n513), .ZN(new_n1121));
  INV_X1    g0921(.A(G283), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n725), .A2(new_n1122), .B1(new_n727), .B2(new_n265), .ZN(new_n1123));
  OR3_X1    g0923(.A1(new_n1120), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n747), .A2(new_n225), .B1(new_n515), .B2(new_n740), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT117), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n750), .A2(G125), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n398), .B(new_n1127), .C1(G128), .C2(new_n724), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n736), .A2(G150), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1129), .B(KEYINPUT53), .Z(new_n1130));
  OAI211_X1 g0930(.A(new_n1128), .B(new_n1130), .C1(new_n201), .C2(new_n733), .ZN(new_n1131));
  XOR2_X1   g0931(.A(KEYINPUT54), .B(G143), .Z(new_n1132));
  AOI22_X1  g0932(.A1(G137), .A2(new_n726), .B1(new_n742), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(G159), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1133), .B1(new_n818), .B2(new_n740), .C1(new_n747), .C2(new_n1134), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n1124), .A2(new_n1126), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1118), .B1(new_n1136), .B2(new_n766), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT118), .Z(new_n1138));
  NAND2_X1  g0938(.A1(new_n1117), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1103), .A2(new_n1116), .A3(new_n1139), .ZN(G378));
  OAI21_X1  g0940(.A(new_n807), .B1(G50), .B2(new_n809), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n733), .A2(new_n202), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1143), .B1(new_n1122), .B2(new_n749), .C1(new_n592), .C2(new_n824), .ZN(new_n1144));
  AOI211_X1 g0944(.A(G41), .B(new_n259), .C1(new_n736), .C2(G77), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n513), .B2(new_n727), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n265), .A2(new_n740), .B1(new_n725), .B2(new_n515), .ZN(new_n1147));
  NOR4_X1   g0947(.A1(new_n1144), .A2(new_n997), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  OR2_X1    g0948(.A1(new_n1148), .A2(KEYINPUT58), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(G125), .A2(new_n724), .B1(new_n739), .B2(G128), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G137), .B2(new_n742), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n726), .A2(G132), .B1(new_n736), .B2(new_n1132), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1152), .B(new_n1153), .C1(new_n346), .C2(new_n747), .ZN(new_n1154));
  OR2_X1    g0954(.A1(new_n1154), .A2(KEYINPUT59), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(KEYINPUT59), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n256), .B(new_n303), .C1(new_n733), .C2(new_n1134), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G124), .B2(new_n750), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1155), .A2(new_n1156), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1148), .A2(KEYINPUT58), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n201), .B1(new_n250), .B2(G41), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1149), .A2(new_n1159), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1141), .B1(new_n1162), .B2(new_n766), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n355), .A2(new_n668), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1164), .A2(KEYINPUT55), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(KEYINPUT55), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n384), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n384), .A2(new_n1167), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  OR3_X1    g0971(.A1(new_n1168), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1171), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1163), .B1(new_n1174), .B2(new_n775), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT120), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n883), .A2(new_n839), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n884), .A2(new_n890), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1177), .A2(new_n1178), .A3(G330), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1174), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1177), .A2(new_n1174), .A3(new_n1178), .A4(G330), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT121), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n909), .B2(new_n916), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1176), .B1(new_n1189), .B2(new_n989), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1115), .A2(new_n1111), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT57), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1182), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1174), .B1(new_n891), .B2(G330), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n917), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1181), .A2(new_n909), .A3(new_n916), .A4(new_n1182), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1192), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1191), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1198), .A2(KEYINPUT122), .A3(new_n689), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1115), .A2(new_n1111), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1192), .B1(new_n1200), .B2(new_n1188), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT122), .B1(new_n1198), .B2(new_n689), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1190), .B1(new_n1202), .B2(new_n1203), .ZN(G375));
  INV_X1    g1004(.A(new_n958), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1110), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1112), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  XOR2_X1   g1007(.A(new_n1207), .B(KEYINPUT123), .Z(new_n1208));
  NAND2_X1  g1008(.A1(new_n911), .A2(new_n774), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n807), .B1(G68), .B2(new_n809), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n724), .A2(G132), .B1(new_n726), .B2(new_n1132), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n398), .B1(new_n736), .B2(G159), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(new_n1002), .C2(new_n740), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1142), .B(new_n1213), .C1(G128), .C2(new_n750), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n747), .A2(new_n201), .B1(new_n346), .B2(new_n824), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT124), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n398), .B1(new_n823), .B2(new_n513), .C1(new_n824), .C2(new_n265), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G77), .B2(new_n734), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n725), .A2(new_n763), .B1(new_n727), .B2(new_n515), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G283), .B2(new_n739), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n750), .A2(G303), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1219), .A2(new_n1051), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1217), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1210), .B1(new_n1224), .B2(new_n766), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1109), .A2(new_n989), .B1(new_n1209), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1208), .A2(new_n1226), .ZN(G381));
  NAND4_X1  g1027(.A1(new_n990), .A2(new_n1062), .A3(new_n1015), .A4(new_n1083), .ZN(new_n1228));
  INV_X1    g1028(.A(G396), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1021), .A2(new_n1058), .A3(new_n1229), .ZN(new_n1230));
  OR3_X1    g1030(.A1(G381), .A2(G384), .A3(new_n1230), .ZN(new_n1231));
  OR4_X1    g1031(.A1(G378), .A2(G375), .A3(new_n1228), .A4(new_n1231), .ZN(G407));
  INV_X1    g1032(.A(G378), .ZN(new_n1233));
  INV_X1    g1033(.A(G213), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1234), .A2(G343), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1233), .A2(new_n1235), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G407), .B(G213), .C1(G375), .C2(new_n1236), .ZN(G409));
  INV_X1    g1037(.A(KEYINPUT61), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(G387), .A2(G390), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1026), .A2(new_n1057), .ZN(new_n1240));
  OAI21_X1  g1040(.A(G396), .B1(new_n1240), .B2(new_n1020), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1230), .A2(new_n1241), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1239), .A2(new_n1242), .A3(new_n1228), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1242), .B1(new_n1239), .B2(new_n1228), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(G378), .B(new_n1190), .C1(new_n1202), .C2(new_n1203), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1189), .A2(new_n1205), .A3(new_n1191), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1176), .B1(new_n1248), .B2(new_n989), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1233), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1235), .B1(new_n1246), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1235), .A2(G2897), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1206), .ZN(new_n1255));
  OAI21_X1  g1055(.A(KEYINPUT60), .B1(new_n1255), .B2(new_n1114), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT60), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1206), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1256), .A2(new_n689), .A3(new_n1258), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1259), .A2(new_n836), .A3(new_n833), .A4(new_n1226), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT126), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1257), .B1(new_n1112), .B2(new_n1206), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1258), .A2(new_n689), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1226), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(G384), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1260), .A2(new_n1261), .A3(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1261), .B1(new_n1260), .B2(new_n1265), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1254), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1260), .A2(new_n1265), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT126), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1260), .A2(new_n1261), .A3(new_n1265), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1270), .A2(new_n1253), .A3(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1268), .A2(new_n1272), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1238), .B(new_n1245), .C1(new_n1252), .C2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1269), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n1235), .B(new_n1276), .C1(new_n1246), .C2(new_n1251), .ZN(new_n1277));
  OAI21_X1  g1077(.A(KEYINPUT63), .B1(new_n1277), .B2(KEYINPUT125), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1252), .A2(new_n1269), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT125), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1275), .A2(new_n1278), .A3(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT62), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1252), .A2(new_n1284), .A3(new_n1269), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1238), .B1(new_n1252), .B2(new_n1273), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1284), .B1(new_n1252), .B2(new_n1269), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n1285), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1283), .B1(new_n1288), .B2(new_n1245), .ZN(G405));
  INV_X1    g1089(.A(KEYINPUT127), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1246), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1245), .A2(new_n1291), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1293), .A2(new_n1290), .A3(new_n1246), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1276), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1292), .A2(new_n1269), .A3(new_n1294), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1296), .A2(new_n1233), .A3(G375), .A4(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(G375), .A2(new_n1233), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1292), .A2(new_n1269), .A3(new_n1294), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1269), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1299), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1298), .A2(new_n1302), .ZN(G402));
endmodule


