

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U557 ( .A1(n812), .A2(n811), .ZN(n522) );
  OR2_X1 U558 ( .A1(n777), .A2(n776), .ZN(n523) );
  OR2_X1 U559 ( .A1(n777), .A2(n766), .ZN(n524) );
  AND2_X1 U560 ( .A1(n774), .A2(n773), .ZN(n525) );
  INV_X1 U561 ( .A(KEYINPUT95), .ZN(n705) );
  XNOR2_X1 U562 ( .A(n692), .B(n732), .ZN(n704) );
  NAND2_X1 U563 ( .A1(n524), .A2(n946), .ZN(n767) );
  OR2_X1 U564 ( .A1(n768), .A2(n767), .ZN(n774) );
  NOR2_X2 U565 ( .A1(n530), .A2(G2105), .ZN(n892) );
  NOR2_X1 U566 ( .A1(G651), .A2(n622), .ZN(n641) );
  NOR2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  XOR2_X2 U568 ( .A(KEYINPUT17), .B(n526), .Z(n889) );
  NAND2_X1 U569 ( .A1(G137), .A2(n889), .ZN(n528) );
  INV_X1 U570 ( .A(G2104), .ZN(n530) );
  INV_X1 U571 ( .A(G2105), .ZN(n533) );
  NOR2_X1 U572 ( .A1(n530), .A2(n533), .ZN(n884) );
  NAND2_X1 U573 ( .A1(G113), .A2(n884), .ZN(n527) );
  NAND2_X1 U574 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U575 ( .A(n529), .B(KEYINPUT66), .ZN(n538) );
  NAND2_X1 U576 ( .A1(G101), .A2(n892), .ZN(n531) );
  XNOR2_X1 U577 ( .A(n531), .B(KEYINPUT65), .ZN(n532) );
  XNOR2_X1 U578 ( .A(n532), .B(KEYINPUT23), .ZN(n536) );
  NOR2_X1 U579 ( .A1(n533), .A2(G2104), .ZN(n534) );
  XNOR2_X1 U580 ( .A(n534), .B(KEYINPUT64), .ZN(n885) );
  NAND2_X1 U581 ( .A1(G125), .A2(n885), .ZN(n535) );
  NAND2_X1 U582 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X2 U583 ( .A1(n538), .A2(n537), .ZN(G160) );
  NOR2_X1 U584 ( .A1(G543), .A2(G651), .ZN(n646) );
  NAND2_X1 U585 ( .A1(G90), .A2(n646), .ZN(n540) );
  XOR2_X1 U586 ( .A(G543), .B(KEYINPUT0), .Z(n622) );
  INV_X1 U587 ( .A(G651), .ZN(n544) );
  NOR2_X1 U588 ( .A1(n622), .A2(n544), .ZN(n650) );
  NAND2_X1 U589 ( .A1(G77), .A2(n650), .ZN(n539) );
  NAND2_X1 U590 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U591 ( .A(n541), .B(KEYINPUT9), .ZN(n543) );
  NAND2_X1 U592 ( .A1(G52), .A2(n641), .ZN(n542) );
  NAND2_X1 U593 ( .A1(n543), .A2(n542), .ZN(n548) );
  NOR2_X1 U594 ( .A1(G543), .A2(n544), .ZN(n545) );
  XOR2_X1 U595 ( .A(KEYINPUT1), .B(n545), .Z(n642) );
  NAND2_X1 U596 ( .A1(n642), .A2(G64), .ZN(n546) );
  XOR2_X1 U597 ( .A(KEYINPUT70), .B(n546), .Z(n547) );
  NOR2_X1 U598 ( .A1(n548), .A2(n547), .ZN(G171) );
  AND2_X1 U599 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U600 ( .A(G120), .ZN(G236) );
  INV_X1 U601 ( .A(G132), .ZN(G219) );
  INV_X1 U602 ( .A(G82), .ZN(G220) );
  NAND2_X1 U603 ( .A1(n646), .A2(G89), .ZN(n549) );
  XNOR2_X1 U604 ( .A(n549), .B(KEYINPUT4), .ZN(n551) );
  NAND2_X1 U605 ( .A1(G76), .A2(n650), .ZN(n550) );
  NAND2_X1 U606 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U607 ( .A(KEYINPUT5), .B(n552), .ZN(n558) );
  NAND2_X1 U608 ( .A1(n642), .A2(G63), .ZN(n553) );
  XOR2_X1 U609 ( .A(KEYINPUT75), .B(n553), .Z(n555) );
  NAND2_X1 U610 ( .A1(n641), .A2(G51), .ZN(n554) );
  NAND2_X1 U611 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U612 ( .A(KEYINPUT6), .B(n556), .Z(n557) );
  NAND2_X1 U613 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U614 ( .A(KEYINPUT7), .B(n559), .ZN(G168) );
  XOR2_X1 U615 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U616 ( .A1(G7), .A2(G661), .ZN(n560) );
  XNOR2_X1 U617 ( .A(n560), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U618 ( .A(G223), .ZN(n830) );
  NAND2_X1 U619 ( .A1(n830), .A2(G567), .ZN(n561) );
  XOR2_X1 U620 ( .A(KEYINPUT11), .B(n561), .Z(G234) );
  NAND2_X1 U621 ( .A1(G56), .A2(n642), .ZN(n562) );
  XOR2_X1 U622 ( .A(KEYINPUT14), .B(n562), .Z(n569) );
  NAND2_X1 U623 ( .A1(G81), .A2(n646), .ZN(n563) );
  XOR2_X1 U624 ( .A(KEYINPUT73), .B(n563), .Z(n564) );
  XNOR2_X1 U625 ( .A(n564), .B(KEYINPUT12), .ZN(n566) );
  NAND2_X1 U626 ( .A1(G68), .A2(n650), .ZN(n565) );
  NAND2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U628 ( .A(KEYINPUT13), .B(n567), .Z(n568) );
  NOR2_X1 U629 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U630 ( .A1(n641), .A2(G43), .ZN(n570) );
  NAND2_X1 U631 ( .A1(n571), .A2(n570), .ZN(n968) );
  INV_X1 U632 ( .A(G860), .ZN(n593) );
  OR2_X1 U633 ( .A1(n968), .A2(n593), .ZN(G153) );
  INV_X1 U634 ( .A(G171), .ZN(G301) );
  NAND2_X1 U635 ( .A1(G868), .A2(G301), .ZN(n581) );
  NAND2_X1 U636 ( .A1(G92), .A2(n646), .ZN(n573) );
  NAND2_X1 U637 ( .A1(G66), .A2(n642), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(KEYINPUT74), .B(n574), .ZN(n578) );
  NAND2_X1 U640 ( .A1(G54), .A2(n641), .ZN(n576) );
  NAND2_X1 U641 ( .A1(G79), .A2(n650), .ZN(n575) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U644 ( .A(KEYINPUT15), .B(n579), .Z(n960) );
  INV_X1 U645 ( .A(n960), .ZN(n903) );
  INV_X1 U646 ( .A(G868), .ZN(n653) );
  NAND2_X1 U647 ( .A1(n903), .A2(n653), .ZN(n580) );
  NAND2_X1 U648 ( .A1(n581), .A2(n580), .ZN(G284) );
  NAND2_X1 U649 ( .A1(G65), .A2(n642), .ZN(n582) );
  XNOR2_X1 U650 ( .A(n582), .B(KEYINPUT72), .ZN(n589) );
  NAND2_X1 U651 ( .A1(G53), .A2(n641), .ZN(n584) );
  NAND2_X1 U652 ( .A1(G78), .A2(n650), .ZN(n583) );
  NAND2_X1 U653 ( .A1(n584), .A2(n583), .ZN(n587) );
  NAND2_X1 U654 ( .A1(G91), .A2(n646), .ZN(n585) );
  XNOR2_X1 U655 ( .A(KEYINPUT71), .B(n585), .ZN(n586) );
  NOR2_X1 U656 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U657 ( .A1(n589), .A2(n588), .ZN(G299) );
  NOR2_X1 U658 ( .A1(G868), .A2(G299), .ZN(n590) );
  XNOR2_X1 U659 ( .A(n590), .B(KEYINPUT76), .ZN(n592) );
  NOR2_X1 U660 ( .A1(n653), .A2(G286), .ZN(n591) );
  NOR2_X1 U661 ( .A1(n592), .A2(n591), .ZN(G297) );
  NAND2_X1 U662 ( .A1(n593), .A2(G559), .ZN(n594) );
  NAND2_X1 U663 ( .A1(n594), .A2(n960), .ZN(n595) );
  XNOR2_X1 U664 ( .A(n595), .B(KEYINPUT77), .ZN(n596) );
  XOR2_X1 U665 ( .A(KEYINPUT16), .B(n596), .Z(G148) );
  NOR2_X1 U666 ( .A1(G868), .A2(n968), .ZN(n599) );
  NAND2_X1 U667 ( .A1(n960), .A2(G868), .ZN(n597) );
  NOR2_X1 U668 ( .A1(G559), .A2(n597), .ZN(n598) );
  NOR2_X1 U669 ( .A1(n599), .A2(n598), .ZN(G282) );
  NAND2_X1 U670 ( .A1(G99), .A2(n892), .ZN(n601) );
  NAND2_X1 U671 ( .A1(G111), .A2(n884), .ZN(n600) );
  NAND2_X1 U672 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U673 ( .A(KEYINPUT78), .B(n602), .ZN(n607) );
  NAND2_X1 U674 ( .A1(G123), .A2(n885), .ZN(n603) );
  XNOR2_X1 U675 ( .A(n603), .B(KEYINPUT18), .ZN(n605) );
  NAND2_X1 U676 ( .A1(G135), .A2(n889), .ZN(n604) );
  NAND2_X1 U677 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U678 ( .A1(n607), .A2(n606), .ZN(n928) );
  XNOR2_X1 U679 ( .A(n928), .B(G2096), .ZN(n609) );
  INV_X1 U680 ( .A(G2100), .ZN(n608) );
  NAND2_X1 U681 ( .A1(n609), .A2(n608), .ZN(G156) );
  NAND2_X1 U682 ( .A1(n960), .A2(G559), .ZN(n663) );
  XNOR2_X1 U683 ( .A(n968), .B(n663), .ZN(n610) );
  NOR2_X1 U684 ( .A1(n610), .A2(G860), .ZN(n618) );
  NAND2_X1 U685 ( .A1(G93), .A2(n646), .ZN(n612) );
  NAND2_X1 U686 ( .A1(G80), .A2(n650), .ZN(n611) );
  NAND2_X1 U687 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U688 ( .A1(G67), .A2(n642), .ZN(n613) );
  XNOR2_X1 U689 ( .A(KEYINPUT79), .B(n613), .ZN(n614) );
  NOR2_X1 U690 ( .A1(n615), .A2(n614), .ZN(n617) );
  NAND2_X1 U691 ( .A1(n641), .A2(G55), .ZN(n616) );
  NAND2_X1 U692 ( .A1(n617), .A2(n616), .ZN(n655) );
  XOR2_X1 U693 ( .A(n618), .B(n655), .Z(G145) );
  NAND2_X1 U694 ( .A1(G49), .A2(n641), .ZN(n620) );
  NAND2_X1 U695 ( .A1(G74), .A2(G651), .ZN(n619) );
  NAND2_X1 U696 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U697 ( .A1(n642), .A2(n621), .ZN(n624) );
  NAND2_X1 U698 ( .A1(n622), .A2(G87), .ZN(n623) );
  NAND2_X1 U699 ( .A1(n624), .A2(n623), .ZN(G288) );
  NAND2_X1 U700 ( .A1(G86), .A2(n646), .ZN(n626) );
  NAND2_X1 U701 ( .A1(G61), .A2(n642), .ZN(n625) );
  NAND2_X1 U702 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U703 ( .A1(n650), .A2(G73), .ZN(n627) );
  XOR2_X1 U704 ( .A(KEYINPUT2), .B(n627), .Z(n628) );
  NOR2_X1 U705 ( .A1(n629), .A2(n628), .ZN(n631) );
  NAND2_X1 U706 ( .A1(n641), .A2(G48), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n631), .A2(n630), .ZN(G305) );
  NAND2_X1 U708 ( .A1(n641), .A2(G47), .ZN(n632) );
  XNOR2_X1 U709 ( .A(n632), .B(KEYINPUT68), .ZN(n639) );
  NAND2_X1 U710 ( .A1(G85), .A2(n646), .ZN(n634) );
  NAND2_X1 U711 ( .A1(G72), .A2(n650), .ZN(n633) );
  NAND2_X1 U712 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U713 ( .A1(G60), .A2(n642), .ZN(n635) );
  XNOR2_X1 U714 ( .A(KEYINPUT67), .B(n635), .ZN(n636) );
  NOR2_X1 U715 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U717 ( .A(KEYINPUT69), .B(n640), .Z(G290) );
  NAND2_X1 U718 ( .A1(G50), .A2(n641), .ZN(n644) );
  NAND2_X1 U719 ( .A1(G62), .A2(n642), .ZN(n643) );
  NAND2_X1 U720 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U721 ( .A(KEYINPUT80), .B(n645), .ZN(n649) );
  NAND2_X1 U722 ( .A1(G88), .A2(n646), .ZN(n647) );
  XNOR2_X1 U723 ( .A(KEYINPUT81), .B(n647), .ZN(n648) );
  NOR2_X1 U724 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U725 ( .A1(n650), .A2(G75), .ZN(n651) );
  NAND2_X1 U726 ( .A1(n652), .A2(n651), .ZN(G303) );
  INV_X1 U727 ( .A(G303), .ZN(G166) );
  AND2_X1 U728 ( .A1(n653), .A2(n655), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n654), .B(KEYINPUT83), .ZN(n666) );
  XNOR2_X1 U730 ( .A(KEYINPUT19), .B(G288), .ZN(n656) );
  XNOR2_X1 U731 ( .A(n656), .B(n655), .ZN(n659) );
  XOR2_X1 U732 ( .A(G290), .B(G299), .Z(n657) );
  XNOR2_X1 U733 ( .A(G305), .B(n657), .ZN(n658) );
  XNOR2_X1 U734 ( .A(n659), .B(n658), .ZN(n661) );
  XNOR2_X1 U735 ( .A(n968), .B(G166), .ZN(n660) );
  XNOR2_X1 U736 ( .A(n661), .B(n660), .ZN(n900) );
  XOR2_X1 U737 ( .A(n900), .B(KEYINPUT82), .Z(n662) );
  XNOR2_X1 U738 ( .A(n663), .B(n662), .ZN(n664) );
  NAND2_X1 U739 ( .A1(G868), .A2(n664), .ZN(n665) );
  NAND2_X1 U740 ( .A1(n666), .A2(n665), .ZN(G295) );
  NAND2_X1 U741 ( .A1(G2078), .A2(G2084), .ZN(n667) );
  XOR2_X1 U742 ( .A(KEYINPUT20), .B(n667), .Z(n668) );
  NAND2_X1 U743 ( .A1(G2090), .A2(n668), .ZN(n670) );
  XNOR2_X1 U744 ( .A(KEYINPUT21), .B(KEYINPUT84), .ZN(n669) );
  XNOR2_X1 U745 ( .A(n670), .B(n669), .ZN(n671) );
  NAND2_X1 U746 ( .A1(G2072), .A2(n671), .ZN(G158) );
  XNOR2_X1 U747 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U748 ( .A1(G220), .A2(G219), .ZN(n672) );
  XOR2_X1 U749 ( .A(KEYINPUT22), .B(n672), .Z(n673) );
  NOR2_X1 U750 ( .A1(G218), .A2(n673), .ZN(n674) );
  XOR2_X1 U751 ( .A(KEYINPUT85), .B(n674), .Z(n675) );
  NAND2_X1 U752 ( .A1(G96), .A2(n675), .ZN(n835) );
  NAND2_X1 U753 ( .A1(n835), .A2(G2106), .ZN(n679) );
  NAND2_X1 U754 ( .A1(G69), .A2(G108), .ZN(n676) );
  NOR2_X1 U755 ( .A1(G236), .A2(n676), .ZN(n677) );
  NAND2_X1 U756 ( .A1(G57), .A2(n677), .ZN(n834) );
  NAND2_X1 U757 ( .A1(n834), .A2(G567), .ZN(n678) );
  NAND2_X1 U758 ( .A1(n679), .A2(n678), .ZN(n837) );
  NAND2_X1 U759 ( .A1(G661), .A2(G483), .ZN(n680) );
  NOR2_X1 U760 ( .A1(n837), .A2(n680), .ZN(n833) );
  NAND2_X1 U761 ( .A1(n833), .A2(G36), .ZN(G176) );
  NAND2_X1 U762 ( .A1(G102), .A2(n892), .ZN(n682) );
  NAND2_X1 U763 ( .A1(G138), .A2(n889), .ZN(n681) );
  NAND2_X1 U764 ( .A1(n682), .A2(n681), .ZN(n686) );
  NAND2_X1 U765 ( .A1(G114), .A2(n884), .ZN(n684) );
  NAND2_X1 U766 ( .A1(G126), .A2(n885), .ZN(n683) );
  NAND2_X1 U767 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U768 ( .A1(n686), .A2(n685), .ZN(G164) );
  NOR2_X1 U769 ( .A1(G164), .A2(G1384), .ZN(n779) );
  NAND2_X1 U770 ( .A1(G160), .A2(G40), .ZN(n778) );
  XOR2_X1 U771 ( .A(KEYINPUT92), .B(n778), .Z(n687) );
  NAND2_X2 U772 ( .A1(n779), .A2(n687), .ZN(n732) );
  INV_X1 U773 ( .A(G1996), .ZN(n1008) );
  NOR2_X1 U774 ( .A1(n732), .A2(n1008), .ZN(n688) );
  XOR2_X1 U775 ( .A(n688), .B(KEYINPUT26), .Z(n699) );
  AND2_X1 U776 ( .A1(n732), .A2(G1341), .ZN(n689) );
  NOR2_X1 U777 ( .A1(n689), .A2(n968), .ZN(n698) );
  AND2_X1 U778 ( .A1(n698), .A2(n960), .ZN(n690) );
  NAND2_X1 U779 ( .A1(n699), .A2(n690), .ZN(n696) );
  NAND2_X1 U780 ( .A1(G1348), .A2(n732), .ZN(n691) );
  XNOR2_X1 U781 ( .A(n691), .B(KEYINPUT96), .ZN(n694) );
  INV_X1 U782 ( .A(KEYINPUT94), .ZN(n692) );
  NAND2_X1 U783 ( .A1(G2067), .A2(n704), .ZN(n693) );
  NAND2_X1 U784 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U785 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U786 ( .A(KEYINPUT97), .B(n697), .ZN(n702) );
  AND2_X1 U787 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U788 ( .A1(n960), .A2(n700), .ZN(n701) );
  NOR2_X1 U789 ( .A1(n702), .A2(n701), .ZN(n710) );
  NAND2_X1 U790 ( .A1(G2072), .A2(n704), .ZN(n703) );
  XOR2_X1 U791 ( .A(KEYINPUT27), .B(n703), .Z(n708) );
  INV_X1 U792 ( .A(n704), .ZN(n717) );
  NAND2_X1 U793 ( .A1(n717), .A2(G1956), .ZN(n706) );
  XNOR2_X1 U794 ( .A(n706), .B(n705), .ZN(n707) );
  NAND2_X1 U795 ( .A1(n708), .A2(n707), .ZN(n712) );
  NOR2_X1 U796 ( .A1(G299), .A2(n712), .ZN(n709) );
  NOR2_X1 U797 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U798 ( .A(n711), .B(KEYINPUT98), .ZN(n715) );
  NAND2_X1 U799 ( .A1(G299), .A2(n712), .ZN(n713) );
  XOR2_X1 U800 ( .A(KEYINPUT28), .B(n713), .Z(n714) );
  NOR2_X1 U801 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U802 ( .A(n716), .B(KEYINPUT29), .ZN(n722) );
  XNOR2_X1 U803 ( .A(G1961), .B(KEYINPUT93), .ZN(n975) );
  NAND2_X1 U804 ( .A1(n732), .A2(n975), .ZN(n720) );
  XNOR2_X1 U805 ( .A(G2078), .B(KEYINPUT25), .ZN(n1007) );
  INV_X1 U806 ( .A(n717), .ZN(n718) );
  NAND2_X1 U807 ( .A1(n1007), .A2(n718), .ZN(n719) );
  NAND2_X1 U808 ( .A1(n720), .A2(n719), .ZN(n723) );
  NAND2_X1 U809 ( .A1(G171), .A2(n723), .ZN(n721) );
  NAND2_X1 U810 ( .A1(n722), .A2(n721), .ZN(n747) );
  NOR2_X1 U811 ( .A1(G171), .A2(n723), .ZN(n724) );
  XOR2_X1 U812 ( .A(KEYINPUT100), .B(n724), .Z(n730) );
  NAND2_X1 U813 ( .A1(G8), .A2(n732), .ZN(n777) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n777), .ZN(n749) );
  NOR2_X1 U815 ( .A1(G2084), .A2(n732), .ZN(n745) );
  NOR2_X1 U816 ( .A1(n749), .A2(n745), .ZN(n725) );
  NAND2_X1 U817 ( .A1(G8), .A2(n725), .ZN(n726) );
  XNOR2_X1 U818 ( .A(KEYINPUT30), .B(n726), .ZN(n727) );
  NOR2_X1 U819 ( .A1(G168), .A2(n727), .ZN(n728) );
  XNOR2_X1 U820 ( .A(KEYINPUT99), .B(n728), .ZN(n729) );
  NAND2_X1 U821 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U822 ( .A(n731), .B(KEYINPUT31), .ZN(n746) );
  INV_X1 U823 ( .A(G8), .ZN(n737) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n732), .ZN(n734) );
  NOR2_X1 U825 ( .A1(G1971), .A2(n777), .ZN(n733) );
  NOR2_X1 U826 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U827 ( .A1(n735), .A2(G303), .ZN(n736) );
  OR2_X1 U828 ( .A1(n737), .A2(n736), .ZN(n739) );
  AND2_X1 U829 ( .A1(n746), .A2(n739), .ZN(n738) );
  NAND2_X1 U830 ( .A1(n747), .A2(n738), .ZN(n742) );
  INV_X1 U831 ( .A(n739), .ZN(n740) );
  OR2_X1 U832 ( .A1(n740), .A2(G286), .ZN(n741) );
  NAND2_X1 U833 ( .A1(n742), .A2(n741), .ZN(n744) );
  XOR2_X1 U834 ( .A(KEYINPUT32), .B(KEYINPUT101), .Z(n743) );
  XNOR2_X1 U835 ( .A(n744), .B(n743), .ZN(n753) );
  NAND2_X1 U836 ( .A1(G8), .A2(n745), .ZN(n751) );
  AND2_X1 U837 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U838 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U839 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n753), .A2(n752), .ZN(n771) );
  NOR2_X1 U841 ( .A1(G1971), .A2(G303), .ZN(n754) );
  NOR2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n951) );
  NOR2_X1 U843 ( .A1(n754), .A2(n951), .ZN(n755) );
  NAND2_X1 U844 ( .A1(n771), .A2(n755), .ZN(n760) );
  INV_X1 U845 ( .A(n777), .ZN(n758) );
  NAND2_X1 U846 ( .A1(G288), .A2(G1976), .ZN(n756) );
  XOR2_X1 U847 ( .A(KEYINPUT102), .B(n756), .Z(n953) );
  NOR2_X1 U848 ( .A1(KEYINPUT103), .A2(n953), .ZN(n757) );
  AND2_X1 U849 ( .A1(n758), .A2(n757), .ZN(n759) );
  AND2_X1 U850 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U851 ( .A1(KEYINPUT33), .A2(n761), .ZN(n768) );
  INV_X1 U852 ( .A(KEYINPUT103), .ZN(n763) );
  NAND2_X1 U853 ( .A1(n951), .A2(KEYINPUT33), .ZN(n762) );
  NAND2_X1 U854 ( .A1(n763), .A2(n762), .ZN(n765) );
  NAND2_X1 U855 ( .A1(n951), .A2(KEYINPUT103), .ZN(n764) );
  NAND2_X1 U856 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U857 ( .A(G1981), .B(G305), .Z(n946) );
  NOR2_X1 U858 ( .A1(G2090), .A2(G303), .ZN(n769) );
  NAND2_X1 U859 ( .A1(G8), .A2(n769), .ZN(n770) );
  NAND2_X1 U860 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U861 ( .A1(n772), .A2(n777), .ZN(n773) );
  NOR2_X1 U862 ( .A1(G1981), .A2(G305), .ZN(n775) );
  XOR2_X1 U863 ( .A(n775), .B(KEYINPUT24), .Z(n776) );
  NAND2_X1 U864 ( .A1(n525), .A2(n523), .ZN(n813) );
  XNOR2_X1 U865 ( .A(G1986), .B(G290), .ZN(n952) );
  NOR2_X1 U866 ( .A1(n779), .A2(n778), .ZN(n824) );
  AND2_X1 U867 ( .A1(n952), .A2(n824), .ZN(n812) );
  XNOR2_X1 U868 ( .A(G2067), .B(KEYINPUT37), .ZN(n780) );
  XNOR2_X1 U869 ( .A(n780), .B(KEYINPUT86), .ZN(n822) );
  NAND2_X1 U870 ( .A1(G104), .A2(n892), .ZN(n782) );
  NAND2_X1 U871 ( .A1(G140), .A2(n889), .ZN(n781) );
  NAND2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n784) );
  XOR2_X1 U873 ( .A(KEYINPUT34), .B(KEYINPUT87), .Z(n783) );
  XNOR2_X1 U874 ( .A(n784), .B(n783), .ZN(n789) );
  NAND2_X1 U875 ( .A1(G116), .A2(n884), .ZN(n786) );
  NAND2_X1 U876 ( .A1(G128), .A2(n885), .ZN(n785) );
  NAND2_X1 U877 ( .A1(n786), .A2(n785), .ZN(n787) );
  XOR2_X1 U878 ( .A(KEYINPUT35), .B(n787), .Z(n788) );
  NOR2_X1 U879 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U880 ( .A(KEYINPUT36), .B(n790), .ZN(n881) );
  NOR2_X1 U881 ( .A1(n822), .A2(n881), .ZN(n929) );
  NAND2_X1 U882 ( .A1(n824), .A2(n929), .ZN(n820) );
  NAND2_X1 U883 ( .A1(G117), .A2(n884), .ZN(n792) );
  NAND2_X1 U884 ( .A1(G129), .A2(n885), .ZN(n791) );
  NAND2_X1 U885 ( .A1(n792), .A2(n791), .ZN(n795) );
  NAND2_X1 U886 ( .A1(n892), .A2(G105), .ZN(n793) );
  XOR2_X1 U887 ( .A(KEYINPUT38), .B(n793), .Z(n794) );
  NOR2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n797) );
  NAND2_X1 U889 ( .A1(n889), .A2(G141), .ZN(n796) );
  NAND2_X1 U890 ( .A1(n797), .A2(n796), .ZN(n876) );
  NAND2_X1 U891 ( .A1(G1996), .A2(n876), .ZN(n798) );
  XNOR2_X1 U892 ( .A(n798), .B(KEYINPUT89), .ZN(n807) );
  NAND2_X1 U893 ( .A1(G131), .A2(n889), .ZN(n800) );
  NAND2_X1 U894 ( .A1(G119), .A2(n885), .ZN(n799) );
  NAND2_X1 U895 ( .A1(n800), .A2(n799), .ZN(n804) );
  NAND2_X1 U896 ( .A1(G95), .A2(n892), .ZN(n802) );
  NAND2_X1 U897 ( .A1(G107), .A2(n884), .ZN(n801) );
  NAND2_X1 U898 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U900 ( .A(n805), .B(KEYINPUT88), .Z(n875) );
  AND2_X1 U901 ( .A1(G1991), .A2(n875), .ZN(n806) );
  NOR2_X1 U902 ( .A1(n807), .A2(n806), .ZN(n922) );
  XOR2_X1 U903 ( .A(n824), .B(KEYINPUT90), .Z(n808) );
  NOR2_X1 U904 ( .A1(n922), .A2(n808), .ZN(n817) );
  INV_X1 U905 ( .A(n817), .ZN(n809) );
  NAND2_X1 U906 ( .A1(n820), .A2(n809), .ZN(n810) );
  XOR2_X1 U907 ( .A(KEYINPUT91), .B(n810), .Z(n811) );
  NAND2_X1 U908 ( .A1(n813), .A2(n522), .ZN(n827) );
  NOR2_X1 U909 ( .A1(G1996), .A2(n876), .ZN(n924) );
  NOR2_X1 U910 ( .A1(G1986), .A2(G290), .ZN(n814) );
  NOR2_X1 U911 ( .A1(G1991), .A2(n875), .ZN(n927) );
  NOR2_X1 U912 ( .A1(n814), .A2(n927), .ZN(n815) );
  XNOR2_X1 U913 ( .A(n815), .B(KEYINPUT104), .ZN(n816) );
  NOR2_X1 U914 ( .A1(n817), .A2(n816), .ZN(n818) );
  NOR2_X1 U915 ( .A1(n924), .A2(n818), .ZN(n819) );
  XNOR2_X1 U916 ( .A(KEYINPUT39), .B(n819), .ZN(n821) );
  NAND2_X1 U917 ( .A1(n821), .A2(n820), .ZN(n823) );
  NAND2_X1 U918 ( .A1(n822), .A2(n881), .ZN(n921) );
  NAND2_X1 U919 ( .A1(n823), .A2(n921), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U921 ( .A1(n827), .A2(n826), .ZN(n829) );
  XOR2_X1 U922 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n828) );
  XNOR2_X1 U923 ( .A(n829), .B(n828), .ZN(G329) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n830), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U926 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U928 ( .A1(n833), .A2(n832), .ZN(G188) );
  XOR2_X1 U929 ( .A(G69), .B(KEYINPUT106), .Z(G235) );
  XNOR2_X1 U930 ( .A(G108), .B(KEYINPUT115), .ZN(G238) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  NOR2_X1 U933 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U934 ( .A(n836), .B(KEYINPUT107), .ZN(G261) );
  INV_X1 U935 ( .A(G261), .ZN(G325) );
  INV_X1 U936 ( .A(n837), .ZN(G319) );
  XOR2_X1 U937 ( .A(G2100), .B(G2678), .Z(n839) );
  XNOR2_X1 U938 ( .A(KEYINPUT42), .B(KEYINPUT108), .ZN(n838) );
  XNOR2_X1 U939 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U940 ( .A(KEYINPUT109), .B(G2090), .Z(n841) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2072), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U943 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U944 ( .A(KEYINPUT43), .B(G2096), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(n847) );
  XOR2_X1 U946 ( .A(G2078), .B(G2084), .Z(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(G227) );
  XOR2_X1 U948 ( .A(G1976), .B(G1956), .Z(n849) );
  XNOR2_X1 U949 ( .A(G1986), .B(G1966), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U951 ( .A(n850), .B(KEYINPUT41), .Z(n852) );
  XNOR2_X1 U952 ( .A(G1961), .B(G1971), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U954 ( .A(G2474), .B(G1981), .Z(n854) );
  XNOR2_X1 U955 ( .A(G1996), .B(G1991), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n856), .B(n855), .ZN(G229) );
  NAND2_X1 U958 ( .A1(G100), .A2(n892), .ZN(n858) );
  NAND2_X1 U959 ( .A1(G112), .A2(n884), .ZN(n857) );
  NAND2_X1 U960 ( .A1(n858), .A2(n857), .ZN(n865) );
  NAND2_X1 U961 ( .A1(G124), .A2(n885), .ZN(n859) );
  XOR2_X1 U962 ( .A(KEYINPUT44), .B(n859), .Z(n862) );
  NAND2_X1 U963 ( .A1(n889), .A2(G136), .ZN(n860) );
  XOR2_X1 U964 ( .A(KEYINPUT110), .B(n860), .Z(n861) );
  NOR2_X1 U965 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U966 ( .A(n863), .B(KEYINPUT111), .ZN(n864) );
  NOR2_X1 U967 ( .A1(n865), .A2(n864), .ZN(G162) );
  NAND2_X1 U968 ( .A1(G106), .A2(n892), .ZN(n867) );
  NAND2_X1 U969 ( .A1(G142), .A2(n889), .ZN(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U971 ( .A(n868), .B(KEYINPUT45), .ZN(n873) );
  NAND2_X1 U972 ( .A1(G118), .A2(n884), .ZN(n870) );
  NAND2_X1 U973 ( .A1(G130), .A2(n885), .ZN(n869) );
  NAND2_X1 U974 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U975 ( .A(KEYINPUT112), .B(n871), .Z(n872) );
  NAND2_X1 U976 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U977 ( .A(n874), .B(G164), .ZN(n880) );
  XNOR2_X1 U978 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n878) );
  XNOR2_X1 U979 ( .A(n876), .B(n875), .ZN(n877) );
  XNOR2_X1 U980 ( .A(n878), .B(n877), .ZN(n879) );
  XNOR2_X1 U981 ( .A(n880), .B(n879), .ZN(n883) );
  XNOR2_X1 U982 ( .A(n881), .B(n928), .ZN(n882) );
  XNOR2_X1 U983 ( .A(n883), .B(n882), .ZN(n896) );
  NAND2_X1 U984 ( .A1(G115), .A2(n884), .ZN(n887) );
  NAND2_X1 U985 ( .A1(G127), .A2(n885), .ZN(n886) );
  NAND2_X1 U986 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U987 ( .A(n888), .B(KEYINPUT47), .ZN(n891) );
  NAND2_X1 U988 ( .A1(G139), .A2(n889), .ZN(n890) );
  NAND2_X1 U989 ( .A1(n891), .A2(n890), .ZN(n895) );
  NAND2_X1 U990 ( .A1(G103), .A2(n892), .ZN(n893) );
  XNOR2_X1 U991 ( .A(KEYINPUT113), .B(n893), .ZN(n894) );
  NOR2_X1 U992 ( .A1(n895), .A2(n894), .ZN(n932) );
  XOR2_X1 U993 ( .A(n896), .B(n932), .Z(n898) );
  XNOR2_X1 U994 ( .A(G160), .B(G162), .ZN(n897) );
  XNOR2_X1 U995 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U996 ( .A1(G37), .A2(n899), .ZN(G395) );
  XOR2_X1 U997 ( .A(KEYINPUT114), .B(n900), .Z(n902) );
  XNOR2_X1 U998 ( .A(G171), .B(G286), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n905), .ZN(G397) );
  XOR2_X1 U1002 ( .A(G2451), .B(G2430), .Z(n907) );
  XNOR2_X1 U1003 ( .A(G2438), .B(G2443), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n913) );
  XOR2_X1 U1005 ( .A(G2435), .B(G2454), .Z(n909) );
  XNOR2_X1 U1006 ( .A(G1348), .B(G1341), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(n909), .B(n908), .ZN(n911) );
  XOR2_X1 U1008 ( .A(G2446), .B(G2427), .Z(n910) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1010 ( .A(n913), .B(n912), .Z(n914) );
  NAND2_X1 U1011 ( .A1(G14), .A2(n914), .ZN(n920) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n920), .ZN(n917) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(KEYINPUT49), .B(n915), .ZN(n916) );
  NOR2_X1 U1015 ( .A1(n917), .A2(n916), .ZN(n919) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1017 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(G57), .ZN(G237) );
  INV_X1 U1020 ( .A(n920), .ZN(G401) );
  NAND2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n941) );
  XOR2_X1 U1022 ( .A(G2090), .B(G162), .Z(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1024 ( .A(KEYINPUT51), .B(n925), .Z(n939) );
  XOR2_X1 U1025 ( .A(G160), .B(G2084), .Z(n926) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n931) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n937) );
  XOR2_X1 U1029 ( .A(G2072), .B(n932), .Z(n934) );
  XOR2_X1 U1030 ( .A(G164), .B(G2078), .Z(n933) );
  NOR2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1032 ( .A(KEYINPUT50), .B(n935), .Z(n936) );
  NOR2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1036 ( .A(KEYINPUT52), .B(n942), .ZN(n944) );
  INV_X1 U1037 ( .A(KEYINPUT55), .ZN(n943) );
  NAND2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1039 ( .A1(n945), .A2(G29), .ZN(n1030) );
  XNOR2_X1 U1040 ( .A(G16), .B(KEYINPUT56), .ZN(n974) );
  XNOR2_X1 U1041 ( .A(G1966), .B(G168), .ZN(n947) );
  NAND2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(n948), .B(KEYINPUT57), .ZN(n972) );
  XOR2_X1 U1044 ( .A(G1956), .B(KEYINPUT123), .Z(n949) );
  XNOR2_X1 U1045 ( .A(G299), .B(n949), .ZN(n950) );
  NOR2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n955) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n958) );
  XOR2_X1 U1049 ( .A(G1971), .B(G166), .Z(n956) );
  XNOR2_X1 U1050 ( .A(KEYINPUT124), .B(n956), .ZN(n957) );
  NOR2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1052 ( .A(KEYINPUT125), .B(n959), .Z(n966) );
  XNOR2_X1 U1053 ( .A(G1348), .B(n960), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(n961), .B(KEYINPUT121), .ZN(n963) );
  XOR2_X1 U1055 ( .A(G1961), .B(G171), .Z(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(KEYINPUT122), .B(n964), .ZN(n965) );
  NAND2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(KEYINPUT126), .B(n967), .ZN(n970) );
  XNOR2_X1 U1060 ( .A(G1341), .B(n968), .ZN(n969) );
  NOR2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1062 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1063 ( .A1(n974), .A2(n973), .ZN(n1000) );
  INV_X1 U1064 ( .A(G16), .ZN(n998) );
  XNOR2_X1 U1065 ( .A(G5), .B(n975), .ZN(n993) );
  XOR2_X1 U1066 ( .A(G1348), .B(KEYINPUT59), .Z(n976) );
  XNOR2_X1 U1067 ( .A(G4), .B(n976), .ZN(n978) );
  XNOR2_X1 U1068 ( .A(G20), .B(G1956), .ZN(n977) );
  NOR2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n982) );
  XNOR2_X1 U1070 ( .A(G1341), .B(G19), .ZN(n980) );
  XNOR2_X1 U1071 ( .A(G1981), .B(G6), .ZN(n979) );
  NOR2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1074 ( .A(n983), .B(KEYINPUT60), .ZN(n991) );
  XNOR2_X1 U1075 ( .A(G1971), .B(G22), .ZN(n985) );
  XNOR2_X1 U1076 ( .A(G23), .B(G1976), .ZN(n984) );
  NOR2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n988) );
  XNOR2_X1 U1078 ( .A(G1986), .B(KEYINPUT127), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(n986), .B(G24), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1081 ( .A(KEYINPUT58), .B(n989), .ZN(n990) );
  NOR2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(G21), .B(G1966), .ZN(n994) );
  NOR2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(KEYINPUT61), .B(n996), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1028) );
  XOR2_X1 U1089 ( .A(G1991), .B(G25), .Z(n1001) );
  NAND2_X1 U1090 ( .A1(n1001), .A2(G28), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(n1002), .B(KEYINPUT117), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(G2067), .B(G26), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(G33), .B(G2072), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1013) );
  XOR2_X1 U1096 ( .A(n1007), .B(G27), .Z(n1010) );
  XOR2_X1 U1097 ( .A(n1008), .B(G32), .Z(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1099 ( .A(KEYINPUT118), .B(n1011), .Z(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1101 ( .A(KEYINPUT53), .B(n1014), .Z(n1018) );
  XNOR2_X1 U1102 ( .A(KEYINPUT54), .B(G34), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(n1015), .B(KEYINPUT119), .ZN(n1016) );
  XNOR2_X1 U1104 ( .A(G2084), .B(n1016), .ZN(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(KEYINPUT116), .B(G2090), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(G35), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1109 ( .A(n1022), .B(KEYINPUT55), .ZN(n1024) );
  INV_X1 U1110 ( .A(G29), .ZN(n1023) );
  NAND2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(G11), .A2(n1025), .ZN(n1026) );
  XNOR2_X1 U1113 ( .A(KEYINPUT120), .B(n1026), .ZN(n1027) );
  NOR2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1031), .Z(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

