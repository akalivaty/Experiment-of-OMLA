//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 1 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n765,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891;
  XOR2_X1   g000(.A(G15gat), .B(G22gat), .Z(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(new_n206), .B2(G1gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT90), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n204), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G8gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G43gat), .B(G50gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n212), .B(KEYINPUT87), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT15), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT15), .ZN(new_n215));
  INV_X1    g014(.A(G50gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n216), .A2(KEYINPUT89), .A3(G43gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G43gat), .B2(new_n216), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT89), .B1(new_n216), .B2(G43gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n215), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  OR3_X1    g019(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n221), .A2(new_n222), .B1(G29gat), .B2(G36gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n214), .A2(new_n220), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G29gat), .A2(G36gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT88), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n221), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n222), .B1(new_n221), .B2(new_n226), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n225), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n229), .A2(KEYINPUT15), .A3(new_n213), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n231), .A2(KEYINPUT17), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT17), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n233), .B1(new_n224), .B2(new_n230), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n211), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n211), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(new_n231), .ZN(new_n237));
  NAND2_X1  g036(.A1(G229gat), .A2(G233gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT18), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n236), .B(new_n231), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n238), .B(KEYINPUT91), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(KEYINPUT13), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n235), .A2(KEYINPUT18), .A3(new_n237), .A4(new_n238), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n241), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT11), .B(G169gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(G197gat), .ZN(new_n249));
  XOR2_X1   g048(.A(G113gat), .B(G141gat), .Z(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(KEYINPUT12), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n247), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n241), .A2(new_n252), .A3(new_n245), .A4(new_n246), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(KEYINPUT92), .ZN(new_n257));
  OR2_X1    g056(.A1(G183gat), .A2(G190gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(G183gat), .A2(G190gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(KEYINPUT24), .A3(new_n259), .ZN(new_n260));
  OR2_X1    g059(.A1(new_n259), .A2(KEYINPUT24), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT65), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G169gat), .A2(G176gat), .ZN(new_n263));
  INV_X1    g062(.A(G169gat), .ZN(new_n264));
  INV_X1    g063(.A(G176gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT23), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n263), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT64), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n262), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n266), .A2(new_n267), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT25), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n273), .B1(new_n269), .B2(new_n268), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n260), .A2(KEYINPUT65), .A3(new_n261), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n271), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n276), .A2(KEYINPUT66), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT25), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n272), .A3(new_n261), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n278), .B1(new_n279), .B2(new_n268), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n276), .A2(KEYINPUT66), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n277), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT28), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT67), .ZN(new_n284));
  XOR2_X1   g083(.A(new_n284), .B(KEYINPUT68), .Z(new_n285));
  XOR2_X1   g084(.A(KEYINPUT27), .B(G183gat), .Z(new_n286));
  OAI22_X1  g085(.A1(new_n286), .A2(G190gat), .B1(KEYINPUT67), .B2(new_n283), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n285), .B(new_n287), .ZN(new_n288));
  OR2_X1    g087(.A1(new_n266), .A2(KEYINPUT26), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n266), .A2(KEYINPUT26), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n289), .A2(new_n290), .A3(new_n263), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n288), .A2(new_n259), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n282), .A2(new_n292), .ZN(new_n293));
  XOR2_X1   g092(.A(G127gat), .B(G134gat), .Z(new_n294));
  XNOR2_X1  g093(.A(G113gat), .B(G120gat), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n294), .B1(KEYINPUT1), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT69), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT1), .ZN(new_n299));
  INV_X1    g098(.A(new_n294), .ZN(new_n300));
  XOR2_X1   g099(.A(KEYINPUT70), .B(G113gat), .Z(new_n301));
  INV_X1    g100(.A(G120gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n302), .A2(G113gat), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n299), .B(new_n300), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n298), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n293), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G227gat), .ZN(new_n308));
  INV_X1    g107(.A(G233gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n298), .A2(new_n305), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n282), .A2(new_n292), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n307), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT34), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT34), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n307), .A2(new_n316), .A3(new_n311), .A4(new_n313), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n313), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n312), .B1(new_n282), .B2(new_n292), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n310), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n318), .A2(KEYINPUT32), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT33), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G15gat), .B(G43gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(G71gat), .B(G99gat), .ZN(new_n326));
  XOR2_X1   g125(.A(new_n325), .B(new_n326), .Z(new_n327));
  NAND2_X1  g126(.A1(new_n321), .A2(KEYINPUT32), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n328), .A2(new_n315), .A3(new_n317), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n322), .A2(new_n324), .A3(new_n327), .A4(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n324), .A2(new_n327), .ZN(new_n331));
  INV_X1    g130(.A(new_n329), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n328), .B1(new_n317), .B2(new_n315), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  XOR2_X1   g133(.A(G155gat), .B(G162gat), .Z(new_n335));
  XNOR2_X1  g134(.A(G141gat), .B(G148gat), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT2), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n337), .B1(new_n338), .B2(G162gat), .ZN(new_n339));
  OR3_X1    g138(.A1(new_n335), .A2(new_n336), .A3(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n335), .B1(KEYINPUT2), .B2(new_n336), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G197gat), .B(G204gat), .ZN(new_n343));
  AND2_X1   g142(.A1(G211gat), .A2(G218gat), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n343), .B1(KEYINPUT22), .B2(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(G211gat), .A2(G218gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n345), .B(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n349), .A2(KEYINPUT29), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n350), .A2(KEYINPUT79), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT3), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n352), .B1(new_n350), .B2(KEYINPUT79), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n342), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(G228gat), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n355), .A2(new_n309), .ZN(new_n356));
  INV_X1    g155(.A(new_n349), .ZN(new_n357));
  INV_X1    g156(.A(new_n342), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n352), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT29), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n357), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n354), .A2(new_n356), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT80), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n350), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n358), .B1(new_n366), .B2(new_n352), .ZN(new_n367));
  OAI22_X1  g166(.A1(new_n367), .A2(new_n361), .B1(new_n355), .B2(new_n309), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n354), .A2(KEYINPUT80), .A3(new_n356), .A4(new_n362), .ZN(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT31), .B(G50gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n370), .B(KEYINPUT78), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n371), .B(G78gat), .ZN(new_n372));
  INV_X1    g171(.A(G106gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n365), .A2(new_n368), .A3(new_n369), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(G22gat), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n375), .A2(G22gat), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n365), .A2(new_n368), .A3(new_n369), .ZN(new_n379));
  INV_X1    g178(.A(new_n374), .ZN(new_n380));
  AND2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI22_X1  g180(.A1(new_n377), .A2(new_n378), .B1(new_n381), .B2(KEYINPUT81), .ZN(new_n382));
  INV_X1    g181(.A(new_n378), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT81), .B1(new_n379), .B2(new_n380), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n384), .A3(new_n376), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n330), .A2(new_n334), .A3(new_n382), .A4(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  XOR2_X1   g186(.A(KEYINPUT77), .B(KEYINPUT6), .Z(new_n388));
  NAND3_X1  g187(.A1(new_n312), .A2(KEYINPUT74), .A3(new_n358), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n358), .A2(new_n298), .A3(new_n305), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT74), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT4), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n342), .A2(KEYINPUT3), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n359), .A2(new_n306), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT4), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n390), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT5), .ZN(new_n399));
  NAND2_X1  g198(.A1(G225gat), .A2(G233gat), .ZN(new_n400));
  XOR2_X1   g199(.A(new_n400), .B(KEYINPUT73), .Z(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n394), .A2(new_n398), .A3(new_n399), .A4(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT76), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n393), .A2(KEYINPUT4), .B1(new_n397), .B2(new_n390), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n406), .A2(KEYINPUT76), .A3(new_n399), .A4(new_n402), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(KEYINPUT0), .B(G57gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(G85gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(G1gat), .B(G29gat), .ZN(new_n411));
  XOR2_X1   g210(.A(new_n410), .B(new_n411), .Z(new_n412));
  NAND2_X1  g211(.A1(new_n306), .A2(new_n342), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT75), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n389), .B(new_n392), .C1(new_n415), .C2(new_n401), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n401), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n416), .B(new_n396), .C1(new_n415), .C2(new_n390), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n418), .A3(KEYINPUT5), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n408), .A2(new_n412), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n412), .B1(new_n408), .B2(new_n419), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n388), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OR2_X1    g221(.A1(new_n421), .A2(new_n388), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT30), .ZN(new_n424));
  INV_X1    g223(.A(G226gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n425), .A2(new_n309), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n282), .A2(new_n427), .A3(new_n292), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n282), .A2(new_n292), .B1(new_n360), .B2(new_n427), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n349), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n427), .A2(new_n360), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n293), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n433), .A2(new_n357), .A3(new_n428), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  XOR2_X1   g234(.A(G8gat), .B(G36gat), .Z(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(G64gat), .ZN(new_n437));
  INV_X1    g236(.A(G92gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n424), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n435), .A2(new_n439), .ZN(new_n441));
  INV_X1    g240(.A(new_n439), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n431), .A2(new_n434), .A3(KEYINPUT30), .A4(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n440), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n422), .A2(new_n423), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT85), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n387), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n422), .A2(new_n423), .A3(new_n445), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT85), .B1(new_n449), .B2(new_n386), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(KEYINPUT35), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT35), .ZN(new_n452));
  OAI211_X1 g251(.A(KEYINPUT85), .B(new_n452), .C1(new_n449), .C2(new_n386), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n382), .A2(new_n385), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  XOR2_X1   g255(.A(new_n413), .B(KEYINPUT75), .Z(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n402), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT39), .B1(new_n458), .B2(new_n393), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT82), .ZN(new_n460));
  OR2_X1    g259(.A1(new_n406), .A2(new_n402), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT82), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n462), .B(KEYINPUT39), .C1(new_n458), .C2(new_n393), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n460), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  OR2_X1    g263(.A1(new_n461), .A2(KEYINPUT39), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(new_n412), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT40), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n421), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n464), .A2(KEYINPUT40), .A3(new_n412), .A4(new_n465), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n468), .A2(new_n469), .A3(new_n444), .A4(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n422), .A2(new_n423), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT37), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n431), .A2(new_n473), .A3(new_n434), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n473), .B1(new_n431), .B2(new_n434), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT38), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n357), .B1(new_n433), .B2(new_n428), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT83), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n473), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n431), .A2(KEYINPUT83), .A3(new_n434), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT84), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT38), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT84), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n481), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n484), .A2(new_n485), .A3(new_n487), .A4(new_n474), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n439), .A2(KEYINPUT38), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n488), .A2(new_n439), .B1(new_n435), .B2(new_n489), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n456), .B(new_n471), .C1(new_n478), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n449), .A2(new_n455), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n334), .A2(new_n330), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT36), .B1(new_n493), .B2(KEYINPUT71), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT71), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT36), .ZN(new_n496));
  AOI211_X1 g295(.A(new_n495), .B(new_n496), .C1(new_n334), .C2(new_n330), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n491), .A2(new_n492), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n454), .A2(KEYINPUT86), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(new_n453), .A3(new_n451), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT86), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n257), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT21), .ZN(new_n505));
  XNOR2_X1  g304(.A(G57gat), .B(G64gat), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G71gat), .B(G78gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n211), .B1(new_n505), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(KEYINPUT93), .ZN(new_n512));
  NAND2_X1  g311(.A1(G231gat), .A2(G233gat), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n513), .B(KEYINPUT94), .Z(new_n514));
  XNOR2_X1  g313(.A(new_n512), .B(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n510), .A2(new_n505), .ZN(new_n516));
  XOR2_X1   g315(.A(G127gat), .B(G155gat), .Z(new_n517));
  XOR2_X1   g316(.A(new_n516), .B(new_n517), .Z(new_n518));
  XNOR2_X1  g317(.A(new_n515), .B(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n520));
  XNOR2_X1  g319(.A(G183gat), .B(G211gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n519), .B(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(G85gat), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT95), .B1(new_n524), .B2(new_n438), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT95), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n526), .A2(G85gat), .A3(G92gat), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n525), .A2(new_n527), .A3(KEYINPUT7), .ZN(new_n528));
  AOI21_X1  g327(.A(KEYINPUT7), .B1(new_n525), .B2(new_n527), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n524), .A2(KEYINPUT96), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT96), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(G85gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n438), .ZN(new_n535));
  INV_X1    g334(.A(G99gat), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT8), .B1(new_n536), .B2(new_n373), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT97), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(G92gat), .B1(new_n531), .B2(new_n533), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT97), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT8), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n541), .B1(G99gat), .B2(G106gat), .ZN(new_n542));
  NOR3_X1   g341(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n530), .B1(new_n538), .B2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G99gat), .B(G106gat), .Z(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n540), .B1(new_n539), .B2(new_n542), .ZN(new_n548));
  XNOR2_X1  g347(.A(KEYINPUT96), .B(G85gat), .ZN(new_n549));
  OAI211_X1 g348(.A(KEYINPUT97), .B(new_n537), .C1(new_n549), .C2(G92gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n551), .A2(new_n545), .A3(new_n530), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n547), .B(new_n552), .C1(new_n232), .C2(new_n234), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n547), .A2(new_n552), .ZN(new_n554));
  AND2_X1   g353(.A1(G232gat), .A2(G233gat), .ZN(new_n555));
  AOI22_X1  g354(.A1(new_n554), .A2(new_n231), .B1(KEYINPUT41), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G134gat), .B(G162gat), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n557), .B(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n555), .A2(KEYINPUT41), .ZN(new_n561));
  XNOR2_X1  g360(.A(G190gat), .B(G218gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n560), .B(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n510), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n554), .A2(KEYINPUT10), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT98), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n544), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n547), .A2(new_n569), .A3(new_n566), .A4(new_n552), .ZN(new_n570));
  AND3_X1   g369(.A1(new_n551), .A2(new_n545), .A3(new_n530), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n545), .B1(new_n551), .B2(new_n530), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT98), .B1(new_n551), .B2(new_n530), .ZN(new_n573));
  OAI22_X1  g372(.A1(new_n571), .A2(new_n572), .B1(new_n573), .B2(new_n510), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT10), .ZN(new_n576));
  AOI21_X1  g375(.A(KEYINPUT99), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT99), .ZN(new_n578));
  AOI211_X1 g377(.A(new_n578), .B(KEYINPUT10), .C1(new_n570), .C2(new_n574), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n567), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G230gat), .A2(G233gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n581), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n570), .A2(new_n574), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G120gat), .B(G148gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(new_n265), .ZN(new_n587));
  INV_X1    g386(.A(G204gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n589), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n582), .A2(new_n584), .A3(new_n591), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n523), .A2(new_n565), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT100), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT100), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n523), .A2(new_n596), .A3(new_n565), .A4(new_n593), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n504), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT101), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT101), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n504), .A2(new_n602), .A3(new_n599), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n472), .A2(KEYINPUT102), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n472), .A2(KEYINPUT102), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g409(.A(KEYINPUT16), .B(G8gat), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n604), .A2(KEYINPUT42), .A3(new_n444), .A4(new_n612), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n504), .A2(new_n602), .A3(new_n599), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n602), .B1(new_n504), .B2(new_n599), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n444), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT103), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT103), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n604), .A2(new_n618), .A3(new_n444), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n612), .A2(KEYINPUT42), .ZN(new_n620));
  AND3_X1   g419(.A1(new_n617), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n210), .A2(KEYINPUT42), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n613), .B1(new_n621), .B2(new_n622), .ZN(G1325gat));
  INV_X1    g422(.A(new_n493), .ZN(new_n624));
  AOI21_X1  g423(.A(G15gat), .B1(new_n604), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n498), .B1(new_n601), .B2(new_n603), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n625), .B1(G15gat), .B2(new_n626), .ZN(G1326gat));
  NAND2_X1  g426(.A1(new_n604), .A2(new_n455), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT43), .B(G22gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(G1327gat));
  INV_X1    g429(.A(new_n593), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n523), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n504), .A2(new_n564), .A3(new_n632), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n633), .A2(G29gat), .A3(new_n607), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n634), .B(KEYINPUT45), .Z(new_n635));
  AOI21_X1  g434(.A(KEYINPUT86), .B1(new_n454), .B2(new_n499), .ZN(new_n636));
  AND4_X1   g435(.A1(KEYINPUT86), .A2(new_n499), .A3(new_n453), .A4(new_n451), .ZN(new_n637));
  OAI211_X1 g436(.A(KEYINPUT44), .B(new_n564), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n501), .A2(new_n564), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT44), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n638), .A2(new_n256), .A3(new_n632), .A4(new_n641), .ZN(new_n642));
  OR3_X1    g441(.A1(new_n642), .A2(KEYINPUT104), .A3(new_n607), .ZN(new_n643));
  OAI21_X1  g442(.A(KEYINPUT104), .B1(new_n642), .B2(new_n607), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n643), .A2(G29gat), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n635), .A2(new_n645), .ZN(G1328gat));
  NOR3_X1   g445(.A1(new_n633), .A2(G36gat), .A3(new_n445), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT46), .ZN(new_n648));
  OAI21_X1  g447(.A(G36gat), .B1(new_n642), .B2(new_n445), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(G1329gat));
  OR3_X1    g449(.A1(new_n633), .A2(G43gat), .A3(new_n493), .ZN(new_n651));
  OAI21_X1  g450(.A(G43gat), .B1(new_n642), .B2(new_n498), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n651), .A2(new_n652), .A3(KEYINPUT47), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(KEYINPUT106), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT106), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n655), .B(G43gat), .C1(new_n642), .C2(new_n498), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n654), .A2(new_n651), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n653), .B1(new_n657), .B2(new_n658), .ZN(G1330gat));
  OAI21_X1  g458(.A(new_n216), .B1(new_n633), .B2(new_n456), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n455), .A2(G50gat), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n660), .B1(new_n642), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT48), .ZN(G1331gat));
  AOI21_X1  g462(.A(new_n256), .B1(new_n454), .B2(new_n499), .ZN(new_n664));
  INV_X1    g463(.A(new_n523), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n665), .A2(new_n564), .A3(new_n593), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n608), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g468(.A(new_n444), .B(KEYINPUT107), .Z(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n671), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT49), .B(G64gat), .Z(new_n673));
  OAI21_X1  g472(.A(new_n672), .B1(new_n671), .B2(new_n673), .ZN(G1333gat));
  INV_X1    g473(.A(new_n667), .ZN(new_n675));
  OAI21_X1  g474(.A(G71gat), .B1(new_n675), .B2(new_n498), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n675), .A2(G71gat), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n676), .B1(new_n493), .B2(new_n677), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g478(.A1(new_n667), .A2(new_n455), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g480(.A1(new_n523), .A2(new_n256), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n501), .A2(new_n564), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n683), .B(KEYINPUT51), .Z(new_n684));
  AND2_X1   g483(.A1(new_n684), .A2(new_n631), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n685), .A2(new_n534), .A3(new_n608), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n638), .A2(new_n631), .A3(new_n641), .A4(new_n682), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n549), .B1(new_n688), .B2(new_n607), .ZN(new_n689));
  AND3_X1   g488(.A1(new_n686), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n687), .B1(new_n686), .B2(new_n689), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(G1336gat));
  AND4_X1   g491(.A1(new_n438), .A2(new_n684), .A3(new_n631), .A4(new_n670), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(KEYINPUT109), .A2(KEYINPUT52), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT52), .ZN(new_n696));
  INV_X1    g495(.A(new_n670), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n696), .B(G92gat), .C1(new_n688), .C2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n694), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n688), .A2(new_n445), .ZN(new_n700));
  AOI22_X1  g499(.A1(new_n693), .A2(KEYINPUT109), .B1(new_n700), .B2(G92gat), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n699), .B1(new_n701), .B2(new_n696), .ZN(G1337gat));
  XOR2_X1   g501(.A(KEYINPUT110), .B(G99gat), .Z(new_n703));
  NAND3_X1  g502(.A1(new_n624), .A2(new_n631), .A3(new_n703), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n704), .B(KEYINPUT111), .Z(new_n705));
  NAND2_X1  g504(.A1(new_n684), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n688), .A2(new_n498), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n706), .B1(new_n707), .B2(new_n703), .ZN(G1338gat));
  NAND3_X1  g507(.A1(new_n685), .A2(new_n373), .A3(new_n455), .ZN(new_n709));
  OAI21_X1  g508(.A(G106gat), .B1(new_n688), .B2(new_n456), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT53), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT53), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n709), .A2(new_n713), .A3(new_n710), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(G1339gat));
  OAI211_X1 g514(.A(new_n583), .B(new_n567), .C1(new_n577), .C2(new_n579), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n582), .A2(KEYINPUT54), .A3(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT54), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n580), .A2(new_n718), .A3(new_n581), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n717), .A2(KEYINPUT55), .A3(new_n589), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n592), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n719), .A2(new_n589), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT55), .B1(new_n722), .B2(new_n717), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT112), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT55), .ZN(new_n725));
  INV_X1    g524(.A(new_n717), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n719), .A2(new_n589), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT112), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n728), .A2(new_n729), .A3(new_n592), .A4(new_n720), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n724), .A2(new_n256), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n238), .B1(new_n235), .B2(new_n237), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n242), .A2(new_n244), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n251), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n255), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n631), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n564), .B1(new_n731), .B2(new_n736), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n564), .A2(new_n735), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n724), .A2(new_n738), .A3(new_n730), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n665), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n594), .A2(new_n256), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n456), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(KEYINPUT113), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT113), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n744), .A2(new_n747), .A3(new_n456), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n624), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n608), .A2(new_n697), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(G113gat), .B1(new_n753), .B2(new_n257), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n607), .B1(new_n741), .B2(new_n743), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n755), .A2(new_n387), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n697), .ZN(new_n757));
  INV_X1    g556(.A(new_n256), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n758), .A2(new_n301), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n754), .B1(new_n757), .B2(new_n759), .ZN(G1340gat));
  OAI21_X1  g559(.A(G120gat), .B1(new_n753), .B2(new_n593), .ZN(new_n761));
  INV_X1    g560(.A(new_n757), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n762), .A2(new_n302), .A3(new_n631), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(G1341gat));
  AOI21_X1  g563(.A(G127gat), .B1(new_n762), .B2(new_n523), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n523), .A2(G127gat), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n765), .B1(new_n752), .B2(new_n766), .ZN(G1342gat));
  OAI21_X1  g566(.A(G134gat), .B1(new_n753), .B2(new_n565), .ZN(new_n768));
  INV_X1    g567(.A(G134gat), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n565), .A2(new_n444), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n756), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT56), .Z(new_n772));
  NAND2_X1  g571(.A1(new_n768), .A2(new_n772), .ZN(G1343gat));
  INV_X1    g572(.A(new_n498), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(new_n456), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n755), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n776), .A2(new_n670), .ZN(new_n777));
  INV_X1    g576(.A(G141gat), .ZN(new_n778));
  INV_X1    g577(.A(new_n257), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT116), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n751), .A2(new_n774), .ZN(new_n782));
  INV_X1    g581(.A(new_n736), .ZN(new_n783));
  OR2_X1    g582(.A1(new_n723), .A2(KEYINPUT115), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n723), .A2(KEYINPUT115), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n257), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n721), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n783), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n739), .B1(new_n788), .B2(new_n564), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n742), .B1(new_n789), .B2(new_n665), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT57), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n790), .A2(new_n791), .A3(new_n456), .ZN(new_n792));
  XOR2_X1   g591(.A(KEYINPUT114), .B(KEYINPUT57), .Z(new_n793));
  AOI21_X1  g592(.A(new_n793), .B1(new_n744), .B2(new_n455), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n782), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n795), .A2(new_n758), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(new_n778), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT58), .B1(new_n781), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(G141gat), .B1(new_n795), .B2(new_n257), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT58), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(new_n800), .A3(new_n780), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n801), .ZN(G1344gat));
  NOR4_X1   g601(.A1(new_n776), .A2(G148gat), .A3(new_n593), .A4(new_n670), .ZN(new_n803));
  XOR2_X1   g602(.A(new_n803), .B(KEYINPUT117), .Z(new_n804));
  INV_X1    g603(.A(KEYINPUT59), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n805), .B(G148gat), .C1(new_n795), .C2(new_n593), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(KEYINPUT118), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n731), .A2(new_n736), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n565), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n523), .B1(new_n809), .B2(new_n739), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n455), .B(new_n793), .C1(new_n810), .C2(new_n742), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT119), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n595), .A2(new_n257), .A3(new_n597), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n738), .A2(new_n787), .A3(new_n728), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n788), .B2(new_n564), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n813), .B1(new_n815), .B2(new_n665), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n791), .B1(new_n816), .B2(new_n456), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n744), .A2(new_n818), .A3(new_n455), .A4(new_n793), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n812), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(new_n631), .A3(new_n782), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n805), .B1(new_n821), .B2(G148gat), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n804), .B1(new_n807), .B2(new_n822), .ZN(G1345gat));
  INV_X1    g622(.A(G155gat), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n795), .A2(new_n824), .A3(new_n665), .ZN(new_n825));
  AOI21_X1  g624(.A(G155gat), .B1(new_n777), .B2(new_n523), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(G1346gat));
  XOR2_X1   g626(.A(KEYINPUT72), .B(G162gat), .Z(new_n828));
  OAI21_X1  g627(.A(new_n828), .B1(new_n795), .B2(new_n565), .ZN(new_n829));
  INV_X1    g628(.A(new_n828), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n770), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n829), .B1(new_n776), .B2(new_n831), .ZN(G1347gat));
  NAND2_X1  g631(.A1(new_n607), .A2(new_n444), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n746), .A2(new_n624), .A3(new_n748), .A4(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n264), .B1(new_n836), .B2(new_n779), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n837), .A2(KEYINPUT121), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(KEYINPUT121), .ZN(new_n839));
  AOI211_X1 g638(.A(new_n608), .B(new_n697), .C1(new_n741), .C2(new_n743), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n387), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n841), .A2(G169gat), .A3(new_n758), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(KEYINPUT120), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n838), .A2(new_n839), .A3(new_n843), .ZN(G1348gat));
  INV_X1    g643(.A(new_n841), .ZN(new_n845));
  AOI21_X1  g644(.A(G176gat), .B1(new_n845), .B2(new_n631), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n835), .A2(new_n593), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n847), .B2(G176gat), .ZN(G1349gat));
  OAI21_X1  g647(.A(G183gat), .B1(new_n835), .B2(new_n665), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n665), .A2(new_n286), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n849), .B1(new_n841), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n852));
  XOR2_X1   g651(.A(new_n851), .B(new_n852), .Z(G1350gat));
  OR3_X1    g652(.A1(new_n841), .A2(G190gat), .A3(new_n565), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT61), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n836), .A2(new_n564), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n856), .B2(G190gat), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n855), .B(G190gat), .C1(new_n835), .C2(new_n565), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n854), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g661(.A(KEYINPUT123), .B(new_n854), .C1(new_n857), .C2(new_n859), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(G1351gat));
  AND2_X1   g663(.A1(new_n840), .A2(new_n775), .ZN(new_n865));
  INV_X1    g664(.A(G197gat), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(new_n866), .A3(new_n256), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n833), .A2(new_n774), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(KEYINPUT125), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT124), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n820), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n812), .A2(new_n817), .A3(KEYINPUT124), .A4(new_n819), .ZN(new_n872));
  AOI211_X1 g671(.A(new_n257), .B(new_n869), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n867), .B1(new_n873), .B2(new_n866), .ZN(G1352gat));
  NAND3_X1  g673(.A1(new_n865), .A2(new_n588), .A3(new_n631), .ZN(new_n875));
  XOR2_X1   g674(.A(new_n875), .B(KEYINPUT62), .Z(new_n876));
  AOI211_X1 g675(.A(new_n593), .B(new_n869), .C1(new_n871), .C2(new_n872), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n588), .B2(new_n877), .ZN(G1353gat));
  INV_X1    g677(.A(new_n869), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n820), .A2(new_n523), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(G211gat), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n881), .B(KEYINPUT63), .Z(new_n882));
  INV_X1    g681(.A(G211gat), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n865), .A2(new_n883), .A3(new_n523), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(G1354gat));
  AOI21_X1  g684(.A(G218gat), .B1(new_n865), .B2(new_n564), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n872), .ZN(new_n887));
  AOI21_X1  g686(.A(KEYINPUT126), .B1(new_n887), .B2(new_n879), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT126), .ZN(new_n889));
  AOI211_X1 g688(.A(new_n889), .B(new_n869), .C1(new_n871), .C2(new_n872), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n888), .A2(new_n890), .A3(new_n565), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n886), .B1(new_n891), .B2(G218gat), .ZN(G1355gat));
endmodule


