//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1283, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342;
  INV_X1    g0000(.A(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G58), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT64), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g0015(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n217), .A2(G20), .A3(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT65), .B(G244), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(new_n202), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G107), .A2(G264), .ZN(new_n226));
  NAND4_X1  g0026(.A1(new_n223), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n209), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n212), .B(new_n220), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT66), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  NAND2_X1  g0039(.A1(G68), .A2(G77), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n203), .A2(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n241), .B(KEYINPUT67), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NAND2_X1  g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n217), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(G222), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n256), .A2(G223), .A3(G1698), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n255), .A2(G77), .ZN(new_n260));
  AND3_X1   g0060(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT68), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n250), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n263), .B1(new_n262), .B2(new_n261), .ZN(new_n264));
  INV_X1    g0064(.A(G274), .ZN(new_n265));
  INV_X1    g0065(.A(new_n213), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n265), .B1(new_n266), .B2(new_n249), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G41), .ZN(new_n269));
  INV_X1    g0069(.A(G45), .ZN(new_n270));
  AOI21_X1  g0070(.A(G1), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(new_n271), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n273), .B1(G226), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n264), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G200), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n279), .B1(new_n264), .B2(new_n276), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n278), .A2(G190), .B1(new_n280), .B2(KEYINPUT73), .ZN(new_n281));
  INV_X1    g0081(.A(G13), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G1), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G20), .ZN(new_n284));
  NAND3_X1  g0084(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n284), .A2(new_n215), .A3(new_n216), .A4(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n206), .A2(G20), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G50), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n286), .A2(new_n288), .B1(G50), .B2(new_n284), .ZN(new_n289));
  XOR2_X1   g0089(.A(new_n289), .B(KEYINPUT70), .Z(new_n290));
  INV_X1    g0090(.A(G50), .ZN(new_n291));
  INV_X1    g0091(.A(G58), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(new_n292), .A3(new_n201), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G20), .A2(G33), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n293), .A2(G20), .B1(G150), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(KEYINPUT8), .B(G58), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT69), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OR3_X1    g0098(.A1(new_n297), .A2(new_n292), .A3(KEYINPUT8), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n207), .A2(G33), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n295), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n215), .A2(new_n216), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n285), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n290), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT9), .ZN(new_n307));
  OR2_X1    g0107(.A1(new_n280), .A2(KEYINPUT73), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n281), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT10), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT10), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n281), .A2(new_n308), .A3(new_n311), .A4(new_n307), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n278), .A2(G169), .ZN(new_n314));
  INV_X1    g0114(.A(new_n306), .ZN(new_n315));
  AND2_X1   g0115(.A1(KEYINPUT71), .A2(G179), .ZN(new_n316));
  NOR2_X1   g0116(.A1(KEYINPUT71), .A2(G179), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n277), .A2(new_n319), .ZN(new_n320));
  OR3_X1    g0120(.A1(new_n314), .A2(new_n315), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n313), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n275), .A2(G232), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(new_n272), .B2(new_n268), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n252), .ZN(new_n326));
  AND2_X1   g0126(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n327));
  NOR2_X1   g0127(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n326), .B1(new_n329), .B2(G33), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G226), .A2(G1698), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT80), .ZN(new_n332));
  INV_X1    g0132(.A(G223), .ZN(new_n333));
  OAI22_X1  g0133(.A1(new_n331), .A2(new_n332), .B1(new_n333), .B2(G1698), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n330), .A2(new_n334), .B1(G33), .B2(G87), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT78), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n253), .ZN(new_n337));
  NAND2_X1  g0137(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(G33), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n252), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n332), .B1(new_n340), .B2(new_n331), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g0142(.A(KEYINPUT81), .B(new_n325), .C1(new_n342), .C2(new_n250), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT81), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n250), .B1(new_n335), .B2(new_n341), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n344), .B1(new_n345), .B2(new_n324), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n279), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n345), .A2(new_n324), .ZN(new_n349));
  INV_X1    g0149(.A(G190), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g0152(.A(G58), .B(G68), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n353), .A2(G20), .B1(G159), .B2(new_n294), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT79), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n340), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n339), .A2(KEYINPUT79), .A3(new_n252), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(new_n207), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT7), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(G20), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n358), .A2(new_n359), .B1(new_n360), .B2(new_n340), .ZN(new_n361));
  OAI211_X1 g0161(.A(KEYINPUT16), .B(new_n354), .C1(new_n361), .C2(new_n201), .ZN(new_n362));
  INV_X1    g0162(.A(new_n360), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n251), .B1(new_n327), .B2(new_n328), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n363), .B1(new_n364), .B2(new_n254), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT7), .B1(new_n255), .B2(new_n207), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n354), .B1(new_n367), .B2(new_n201), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT16), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n362), .A2(new_n370), .A3(new_n304), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n300), .B1(new_n206), .B2(G20), .ZN(new_n372));
  INV_X1    g0172(.A(new_n286), .ZN(new_n373));
  INV_X1    g0173(.A(new_n284), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n372), .A2(new_n373), .B1(new_n374), .B2(new_n300), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT17), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n376), .A2(KEYINPUT82), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n352), .A2(new_n371), .A3(new_n375), .A4(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(G200), .B1(new_n343), .B2(new_n346), .ZN(new_n380));
  INV_X1    g0180(.A(new_n351), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n371), .B(new_n375), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  XOR2_X1   g0182(.A(KEYINPUT82), .B(KEYINPUT17), .Z(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AND2_X1   g0184(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n371), .A2(new_n375), .ZN(new_n387));
  INV_X1    g0187(.A(G169), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n347), .A2(new_n388), .B1(new_n349), .B2(new_n318), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT18), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT18), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n387), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n386), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT76), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n252), .A2(new_n254), .A3(G232), .A4(G1698), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n252), .A2(new_n254), .A3(G226), .A4(new_n257), .ZN(new_n399));
  INV_X1    g0199(.A(G97), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n398), .B(new_n399), .C1(new_n251), .C2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n250), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n275), .A2(G238), .B1(new_n271), .B2(new_n267), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT13), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT13), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n403), .A2(new_n407), .A3(new_n404), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(G179), .A3(new_n408), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n409), .B(KEYINPUT75), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n403), .A2(new_n407), .A3(new_n404), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n407), .B1(new_n403), .B2(new_n404), .ZN(new_n412));
  OAI21_X1  g0212(.A(G169), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT14), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n406), .A2(new_n408), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT14), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n415), .A2(new_n416), .A3(G169), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n397), .B1(new_n410), .B2(new_n418), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n414), .A2(new_n417), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT75), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n409), .B(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n420), .A2(new_n422), .A3(KEYINPUT76), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  OR2_X1    g0224(.A1(new_n286), .A2(KEYINPUT72), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n286), .A2(KEYINPUT72), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n201), .B1(new_n206), .B2(G20), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n374), .A2(new_n201), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT12), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n294), .A2(G50), .B1(G20), .B2(new_n201), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(new_n202), .B2(new_n301), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n304), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT11), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n304), .A2(KEYINPUT11), .A3(new_n432), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n428), .A2(new_n430), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  OR2_X1    g0237(.A1(new_n437), .A2(KEYINPUT77), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(KEYINPUT77), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n424), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n437), .B1(new_n415), .B2(G200), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n406), .A2(G190), .A3(new_n408), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT74), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n444), .A2(new_n445), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n443), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n425), .A2(G77), .A3(new_n287), .A4(new_n426), .ZN(new_n450));
  INV_X1    g0250(.A(new_n294), .ZN(new_n451));
  OAI22_X1  g0251(.A1(new_n296), .A2(new_n451), .B1(new_n207), .B2(new_n202), .ZN(new_n452));
  XNOR2_X1  g0252(.A(KEYINPUT15), .B(G87), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(new_n301), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n304), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n374), .A2(new_n202), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n450), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n256), .A2(G232), .A3(new_n257), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n256), .A2(G238), .A3(G1698), .ZN(new_n459));
  INV_X1    g0259(.A(G107), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n458), .B(new_n459), .C1(new_n460), .C2(new_n256), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n402), .ZN(new_n462));
  INV_X1    g0262(.A(new_n221), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n273), .B1(new_n463), .B2(new_n275), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n457), .B1(G200), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n462), .A2(G190), .A3(new_n464), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n465), .A2(new_n388), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n462), .A2(new_n318), .A3(new_n464), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n469), .A2(new_n470), .A3(new_n457), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NOR4_X1   g0272(.A1(new_n322), .A2(new_n396), .A3(new_n449), .A4(new_n472), .ZN(new_n473));
  XNOR2_X1  g0273(.A(KEYINPUT92), .B(KEYINPUT21), .ZN(new_n474));
  MUX2_X1   g0274(.A(G257), .B(G264), .S(G1698), .Z(new_n475));
  NAND2_X1  g0275(.A1(new_n330), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n255), .A2(G303), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT89), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT89), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n476), .A2(new_n480), .A3(new_n477), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n479), .A2(new_n402), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT5), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT84), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n483), .B1(new_n484), .B2(G41), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n269), .A2(KEYINPUT84), .A3(KEYINPUT5), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n270), .A2(G1), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n268), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n266), .A2(new_n249), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n489), .B1(new_n491), .B2(G270), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n388), .B1(new_n482), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n251), .A2(G1), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n425), .A2(G116), .A3(new_n426), .A4(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(G20), .B1(new_n251), .B2(G97), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G283), .ZN(new_n498));
  INV_X1    g0298(.A(G116), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n497), .A2(new_n498), .B1(G20), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n304), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT20), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n304), .A2(KEYINPUT20), .A3(new_n500), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n283), .A2(G20), .A3(new_n499), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n496), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT91), .B1(new_n493), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n481), .A2(new_n402), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n480), .B1(new_n476), .B2(new_n477), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n492), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AND4_X1   g0311(.A1(KEYINPUT91), .A2(new_n511), .A3(new_n507), .A4(G169), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n474), .B1(new_n508), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n507), .B1(new_n511), .B2(G200), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(new_n350), .B2(new_n511), .ZN(new_n515));
  INV_X1    g0315(.A(new_n507), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n511), .A2(KEYINPUT21), .A3(G169), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n482), .A2(G179), .A3(new_n492), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(KEYINPUT90), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT90), .ZN(new_n521));
  AOI211_X1 g0321(.A(new_n521), .B(new_n516), .C1(new_n517), .C2(new_n518), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n513), .B(new_n515), .C1(new_n520), .C2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  OR2_X1    g0324(.A1(G250), .A2(G1698), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(G257), .B2(new_n257), .ZN(new_n526));
  INV_X1    g0326(.A(G294), .ZN(new_n527));
  OAI22_X1  g0327(.A1(new_n340), .A2(new_n526), .B1(new_n251), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n402), .ZN(new_n529));
  INV_X1    g0329(.A(new_n489), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n488), .A2(G264), .A3(new_n490), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G169), .ZN(new_n533));
  XOR2_X1   g0333(.A(new_n531), .B(KEYINPUT95), .Z(new_n534));
  AOI21_X1  g0334(.A(new_n489), .B1(new_n528), .B2(new_n402), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(G179), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n533), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n304), .ZN(new_n539));
  OAI21_X1  g0339(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT94), .ZN(new_n541));
  XNOR2_X1  g0341(.A(new_n540), .B(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT22), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n207), .A2(G87), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n543), .B1(new_n255), .B2(new_n544), .ZN(new_n545));
  OR3_X1    g0345(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n542), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n339), .A2(KEYINPUT22), .A3(G87), .A4(new_n252), .ZN(new_n549));
  NAND2_X1  g0349(.A1(G33), .A2(G116), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n207), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT93), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n548), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(G20), .B1(new_n549), .B2(new_n550), .ZN(new_n555));
  OAI21_X1  g0355(.A(KEYINPUT93), .B1(new_n555), .B2(new_n547), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT24), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT24), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n554), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n539), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n286), .A2(new_n494), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT25), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n284), .B2(G107), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n374), .A2(KEYINPUT25), .A3(new_n460), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n562), .A2(G107), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n538), .B1(new_n561), .B2(new_n567), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n554), .A2(new_n559), .A3(new_n556), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n559), .B1(new_n554), .B2(new_n556), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n304), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n536), .ZN(new_n572));
  OAI22_X1  g0372(.A1(new_n572), .A2(G200), .B1(G190), .B2(new_n532), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n573), .A3(new_n566), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n284), .A2(G97), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(new_n562), .B2(G97), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n460), .A2(KEYINPUT6), .A3(G97), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n400), .A2(new_n460), .ZN(new_n578));
  NOR2_X1   g0378(.A1(G97), .A2(G107), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n577), .B1(new_n580), .B2(KEYINPUT6), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n581), .A2(G20), .B1(G77), .B2(new_n294), .ZN(new_n582));
  OAI21_X1  g0382(.A(G107), .B1(new_n365), .B2(new_n366), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n539), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT83), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n584), .A2(KEYINPUT83), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n576), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n339), .A2(G244), .A3(new_n257), .A4(new_n252), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT4), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AND2_X1   g0391(.A1(KEYINPUT4), .A2(G244), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n252), .A2(new_n254), .A3(new_n592), .A4(new_n257), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n252), .A2(new_n254), .A3(G250), .A4(G1698), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(new_n594), .A3(new_n498), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n402), .B1(new_n591), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n491), .A2(G257), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(new_n530), .A3(new_n597), .ZN(new_n598));
  OR2_X1    g0398(.A1(new_n598), .A2(new_n319), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n388), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n588), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n587), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n585), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n596), .A2(G190), .A3(new_n530), .A4(new_n597), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n598), .A2(G200), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n603), .A2(new_n576), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n568), .A2(new_n574), .A3(new_n601), .A4(new_n606), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n257), .A2(G238), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n330), .A2(new_n608), .B1(G33), .B2(G116), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n330), .A2(KEYINPUT86), .A3(G244), .A4(G1698), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n339), .A2(G244), .A3(G1698), .A4(new_n252), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT86), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n609), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n402), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n490), .B(G250), .C1(G1), .C2(new_n270), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT85), .ZN(new_n617));
  AND4_X1   g0417(.A1(new_n617), .A2(new_n490), .A3(G274), .A4(new_n487), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n617), .B1(new_n267), .B2(new_n487), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n615), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT87), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n620), .B1(new_n614), .B2(new_n402), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT87), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n318), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n207), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT88), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(G87), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n579), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n628), .A2(KEYINPUT88), .A3(new_n207), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n631), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n339), .A2(new_n207), .A3(G68), .A4(new_n252), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT19), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(new_n301), .B2(new_n400), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n635), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n639), .A2(new_n304), .B1(new_n374), .B2(new_n453), .ZN(new_n640));
  INV_X1    g0440(.A(new_n453), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n562), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT87), .B1(new_n615), .B2(new_n621), .ZN(new_n644));
  AOI211_X1 g0444(.A(new_n623), .B(new_n620), .C1(new_n614), .C2(new_n402), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n627), .B(new_n643), .C1(G169), .C2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n624), .A2(G190), .A3(new_n626), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n562), .A2(G87), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n640), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n648), .B(new_n651), .C1(new_n279), .C2(new_n646), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n607), .A2(new_n653), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n473), .A2(new_n524), .A3(new_n654), .ZN(G372));
  AND3_X1   g0455(.A1(new_n588), .A2(new_n599), .A3(new_n600), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n647), .A2(new_n652), .A3(new_n656), .A4(KEYINPUT26), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT97), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n639), .A2(new_n304), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n374), .A2(new_n453), .ZN(new_n660));
  AND4_X1   g0460(.A1(KEYINPUT96), .A2(new_n659), .A3(new_n660), .A4(new_n649), .ZN(new_n661));
  AOI21_X1  g0461(.A(KEYINPUT96), .B1(new_n640), .B2(new_n649), .ZN(new_n662));
  OAI22_X1  g0462(.A1(new_n661), .A2(new_n662), .B1(new_n279), .B2(new_n625), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n663), .B1(G190), .B2(new_n646), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n643), .B1(new_n625), .B2(G169), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n665), .B1(new_n646), .B2(new_n318), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n658), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n662), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n640), .A2(KEYINPUT96), .A3(new_n649), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n668), .A2(new_n669), .B1(new_n622), .B2(G200), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n648), .ZN(new_n671));
  INV_X1    g0471(.A(new_n665), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n627), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n671), .A2(new_n673), .A3(KEYINPUT97), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n601), .B1(new_n667), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n657), .B1(new_n675), .B2(KEYINPUT26), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n574), .A2(new_n601), .A3(new_n606), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n667), .B2(new_n674), .ZN(new_n678));
  INV_X1    g0478(.A(new_n519), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n513), .A2(new_n568), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n666), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n473), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n321), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n440), .B1(new_n419), .B2(new_n423), .ZN(new_n685));
  INV_X1    g0485(.A(new_n448), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(new_n471), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n395), .B1(new_n688), .B2(new_n385), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n684), .B1(new_n689), .B2(new_n313), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n683), .A2(new_n690), .ZN(G369));
  INV_X1    g0491(.A(new_n283), .ZN(new_n692));
  OR3_X1    g0492(.A1(new_n692), .A2(KEYINPUT27), .A3(G20), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT27), .B1(new_n692), .B2(G20), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(G213), .A3(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(G343), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n568), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n574), .ZN(new_n699));
  INV_X1    g0499(.A(new_n697), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n700), .B1(new_n571), .B2(new_n566), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n698), .B1(new_n703), .B2(new_n568), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n513), .A2(new_n679), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n516), .A2(new_n700), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n523), .B2(new_n706), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n704), .A2(G330), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n698), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n513), .B1(new_n520), .B2(new_n522), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n702), .A2(new_n711), .A3(new_n568), .A4(new_n700), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n709), .A2(new_n710), .A3(new_n712), .ZN(G399));
  INV_X1    g0513(.A(new_n210), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G41), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n633), .A2(G116), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(G1), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n218), .B2(new_n716), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  INV_X1    g0520(.A(G330), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT31), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n722), .B1(new_n654), .B2(new_n524), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT98), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n518), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n596), .A2(new_n597), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n536), .A2(new_n726), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n482), .A2(KEYINPUT98), .A3(G179), .A4(new_n492), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n728), .A2(KEYINPUT30), .A3(new_n646), .A4(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT30), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n725), .A2(new_n729), .A3(new_n727), .ZN(new_n732));
  INV_X1    g0532(.A(new_n646), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n572), .A2(new_n319), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n735), .A2(new_n511), .A3(new_n622), .A4(new_n598), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n730), .A2(new_n722), .A3(new_n734), .A4(new_n736), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n737), .A2(new_n697), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n723), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n700), .A2(new_n722), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n730), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n734), .A2(new_n736), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n742), .B1(KEYINPUT99), .B2(new_n743), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n743), .A2(KEYINPUT99), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n741), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n721), .B1(new_n739), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n682), .A2(new_n700), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT29), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n647), .A2(new_n652), .A3(new_n656), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT26), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT100), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n667), .A2(new_n674), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(KEYINPUT26), .A3(new_n656), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n752), .A2(KEYINPUT100), .A3(new_n753), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n756), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n513), .B(new_n568), .C1(new_n520), .C2(new_n522), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n666), .B1(new_n678), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(KEYINPUT29), .A3(new_n700), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n748), .B1(new_n751), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n720), .B1(new_n765), .B2(G1), .ZN(G364));
  NOR2_X1   g0566(.A1(new_n282), .A2(G20), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n206), .B1(new_n767), .B2(G45), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n715), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n770), .B1(new_n708), .B2(G330), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(G330), .B2(new_n708), .ZN(new_n772));
  INV_X1    g0572(.A(new_n770), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n303), .B1(G20), .B2(new_n388), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n207), .A2(new_n350), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n279), .A2(G179), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n207), .A2(G190), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G179), .A2(G200), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI22_X1  g0583(.A1(G303), .A2(new_n779), .B1(new_n783), .B2(G329), .ZN(new_n784));
  INV_X1    g0584(.A(G283), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n780), .A2(new_n777), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n784), .B(new_n255), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n781), .A2(G190), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G20), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n787), .B1(G294), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n319), .A2(new_n279), .A3(new_n780), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n207), .A2(new_n279), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n319), .A2(new_n350), .A3(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(KEYINPUT33), .B(G317), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n792), .A2(G311), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n319), .A2(new_n279), .A3(new_n776), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n319), .A2(G190), .A3(new_n793), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G322), .A2(new_n799), .B1(new_n801), .B2(G326), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n790), .A2(new_n797), .A3(new_n802), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n291), .A2(new_n800), .B1(new_n798), .B2(new_n292), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(G68), .B2(new_n795), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n256), .B1(new_n786), .B2(new_n460), .C1(new_n632), .C2(new_n778), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(G77), .B2(new_n792), .ZN(new_n807));
  INV_X1    g0607(.A(G159), .ZN(new_n808));
  OAI21_X1  g0608(.A(KEYINPUT32), .B1(new_n782), .B2(new_n808), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n782), .A2(KEYINPUT32), .A3(new_n808), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(G97), .B2(new_n789), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n805), .A2(new_n807), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n775), .B1(new_n803), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n244), .A2(G45), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n356), .A2(new_n357), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n714), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n814), .B(new_n816), .C1(G45), .C2(new_n218), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n714), .A2(new_n255), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n818), .A2(G355), .B1(new_n499), .B2(new_n714), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(G13), .A2(G33), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(G20), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n774), .A2(new_n823), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n773), .B(new_n813), .C1(new_n820), .C2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n823), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n825), .B1(new_n708), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n772), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G396));
  NAND2_X1  g0629(.A1(new_n457), .A2(new_n697), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n468), .A2(new_n471), .A3(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT104), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n700), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n657), .ZN(new_n836));
  INV_X1    g0636(.A(new_n674), .ZN(new_n837));
  AOI21_X1  g0637(.A(KEYINPUT97), .B1(new_n671), .B2(new_n673), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n656), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n836), .B1(new_n839), .B2(new_n753), .ZN(new_n840));
  INV_X1    g0640(.A(new_n677), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n841), .B(new_n680), .C1(new_n837), .C2(new_n838), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n673), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n835), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT105), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n682), .A2(KEYINPUT105), .A3(new_n835), .ZN(new_n847));
  INV_X1    g0647(.A(new_n471), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n833), .B1(new_n848), .B2(new_n697), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n846), .A2(new_n847), .B1(new_n749), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n850), .A2(new_n748), .ZN(new_n851));
  OR2_X1    g0651(.A1(new_n851), .A2(KEYINPUT106), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(KEYINPUT106), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n770), .B1(new_n850), .B2(new_n748), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n774), .A2(new_n821), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT101), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n770), .B1(new_n857), .B2(G77), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT102), .ZN(new_n859));
  INV_X1    g0659(.A(G311), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n255), .B1(new_n782), .B2(new_n860), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n778), .A2(new_n460), .B1(new_n786), .B2(new_n632), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n861), .B(new_n862), .C1(G97), .C2(new_n789), .ZN(new_n863));
  AOI22_X1  g0663(.A1(G294), .A2(new_n799), .B1(new_n801), .B2(G303), .ZN(new_n864));
  AOI22_X1  g0664(.A1(G116), .A2(new_n792), .B1(new_n795), .B2(G283), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  AOI22_X1  g0666(.A1(G143), .A2(new_n799), .B1(new_n792), .B2(G159), .ZN(new_n867));
  INV_X1    g0667(.A(G137), .ZN(new_n868));
  INV_X1    g0668(.A(G150), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n867), .B1(new_n868), .B2(new_n800), .C1(new_n869), .C2(new_n794), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT34), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n786), .ZN(new_n873));
  AOI22_X1  g0673(.A1(G50), .A2(new_n779), .B1(new_n873), .B2(G68), .ZN(new_n874));
  INV_X1    g0674(.A(G132), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n874), .B1(new_n875), .B2(new_n782), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(G58), .B2(new_n789), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n872), .A2(new_n815), .A3(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n870), .A2(new_n871), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n866), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n880), .A2(KEYINPUT103), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(KEYINPUT103), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n774), .ZN(new_n883));
  INV_X1    g0683(.A(new_n849), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n859), .B1(new_n881), .B2(new_n883), .C1(new_n884), .C2(new_n822), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n855), .A2(new_n885), .ZN(G384));
  NOR3_X1   g0686(.A1(new_n303), .A2(new_n207), .A3(new_n499), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n581), .B(KEYINPUT107), .Z(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT35), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n890), .B2(new_n889), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n892), .B(KEYINPUT36), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n219), .B(G77), .C1(new_n292), .C2(new_n201), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n291), .A2(G68), .ZN(new_n895));
  AOI211_X1 g0695(.A(new_n206), .B(G13), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n471), .A2(new_n697), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT105), .B1(new_n682), .B2(new_n835), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n845), .B(new_n834), .C1(new_n676), .C2(new_n681), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n375), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n362), .A2(new_n304), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n354), .B1(new_n361), .B2(new_n201), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n369), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n903), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n382), .B1(new_n907), .B2(new_n695), .ZN(new_n908));
  INV_X1    g0708(.A(new_n389), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT37), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n695), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n387), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT37), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n390), .A2(new_n913), .A3(new_n914), .A4(new_n382), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n907), .A2(new_n695), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n385), .B2(new_n394), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT38), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n916), .A2(new_n918), .A3(KEYINPUT38), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n438), .A2(new_n439), .A3(new_n697), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT108), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n924), .B(new_n925), .ZN(new_n926));
  NOR3_X1   g0726(.A1(new_n685), .A2(new_n926), .A3(new_n686), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n419), .A2(new_n423), .A3(new_n448), .ZN(new_n928));
  INV_X1    g0728(.A(new_n924), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT109), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n926), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n442), .A2(new_n932), .A3(new_n448), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT109), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n928), .A2(new_n929), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n931), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n902), .A2(new_n923), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n394), .A2(new_n695), .ZN(new_n939));
  INV_X1    g0739(.A(new_n913), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n385), .B2(new_n394), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n390), .A2(new_n913), .A3(new_n382), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(KEYINPUT37), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n915), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n920), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n922), .ZN(new_n947));
  NOR3_X1   g0747(.A1(new_n947), .A2(KEYINPUT110), .A3(KEYINPUT39), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT39), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n916), .A2(new_n918), .A3(KEYINPUT38), .ZN(new_n950));
  AOI21_X1  g0750(.A(KEYINPUT38), .B1(new_n916), .B2(new_n918), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n946), .A2(KEYINPUT110), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n948), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n442), .A2(new_n697), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n938), .B(new_n939), .C1(new_n955), .C2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n751), .A2(new_n764), .A3(new_n473), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n690), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n958), .B(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n740), .B1(new_n742), .B2(new_n743), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n723), .B2(new_n738), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n937), .A2(new_n884), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT38), .B1(new_n941), .B2(new_n944), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n950), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(KEYINPUT40), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(KEYINPUT40), .B1(new_n921), .B2(new_n922), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n849), .B1(new_n931), .B2(new_n936), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n968), .A2(new_n963), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n971), .A2(new_n473), .A3(new_n963), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n473), .A2(new_n963), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n967), .A2(new_n973), .A3(new_n970), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n972), .A2(G330), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n961), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n206), .B2(new_n767), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n961), .A2(new_n975), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n897), .B1(new_n977), .B2(new_n978), .ZN(G367));
  INV_X1    g0779(.A(KEYINPUT113), .ZN(new_n980));
  INV_X1    g0780(.A(new_n709), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n712), .A2(new_n710), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n656), .A2(new_n697), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n588), .A2(new_n697), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n601), .A2(new_n606), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n982), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT44), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n712), .A2(new_n710), .A3(new_n986), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT45), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n981), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n991), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT44), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n988), .B(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n993), .A2(new_n995), .A3(new_n709), .ZN(new_n996));
  AND2_X1   g0796(.A1(new_n711), .A2(new_n700), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n704), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n712), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n999), .A2(G330), .A3(new_n708), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n708), .A2(G330), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n998), .A2(new_n1001), .A3(new_n712), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n765), .A2(new_n992), .A3(new_n996), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n765), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n715), .B(KEYINPUT41), .Z(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n769), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n704), .A2(new_n997), .A3(KEYINPUT42), .A4(new_n986), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT42), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n712), .B2(new_n987), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n601), .B1(new_n985), .B2(new_n568), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n700), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n668), .A2(new_n669), .A3(new_n697), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n757), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n673), .B2(new_n1016), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(KEYINPUT43), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1015), .A2(KEYINPUT112), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT112), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n1009), .A2(new_n1011), .B1(new_n700), .B2(new_n1013), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1022), .B(new_n1026), .C1(new_n1015), .C2(new_n1020), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n709), .A2(new_n987), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1027), .B(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n980), .B1(new_n1008), .B2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1027), .B(new_n1028), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1006), .B1(new_n1004), .B2(new_n765), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1032), .B(KEYINPUT113), .C1(new_n1033), .C2(new_n769), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n816), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n824), .B1(new_n210), .B2(new_n453), .C1(new_n1036), .C2(new_n238), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n792), .A2(G283), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n799), .A2(G303), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n527), .B2(new_n794), .C1(new_n860), .C2(new_n800), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n873), .A2(G97), .ZN(new_n1042));
  XOR2_X1   g0842(.A(KEYINPUT114), .B(G317), .Z(new_n1043));
  INV_X1    g0843(.A(new_n789), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1042), .B1(new_n782), .B2(new_n1043), .C1(new_n460), .C2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n778), .A2(new_n499), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT46), .ZN(new_n1047));
  NOR4_X1   g0847(.A1(new_n1041), .A2(new_n815), .A3(new_n1045), .A4(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT115), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G143), .A2(new_n801), .B1(new_n795), .B2(G159), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n291), .B2(new_n791), .C1(new_n869), .C2(new_n798), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1044), .A2(new_n201), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n256), .B1(new_n868), .B2(new_n782), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n778), .A2(new_n292), .B1(new_n786), .B2(new_n202), .ZN(new_n1054));
  NOR4_X1   g0854(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1049), .A2(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT47), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n770), .B(new_n1037), .C1(new_n1057), .C2(new_n775), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1018), .A2(new_n826), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1035), .A2(new_n1061), .ZN(G387));
  INV_X1    g0862(.A(new_n717), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n818), .A2(new_n1063), .B1(new_n460), .B2(new_n714), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n235), .A2(new_n270), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n296), .A2(G50), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT50), .Z(new_n1067));
  NAND3_X1  g0867(.A1(new_n717), .A2(new_n270), .A3(new_n240), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n816), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1064), .B1(new_n1065), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n824), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n770), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n704), .A2(new_n826), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1044), .A2(new_n453), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n799), .B2(G50), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT116), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1042), .B1(new_n202), .B2(new_n778), .C1(new_n869), .C2(new_n782), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G68), .B2(new_n792), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n300), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1079), .A2(new_n795), .B1(new_n801), .B2(G159), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1076), .A2(new_n815), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G303), .A2(new_n792), .B1(new_n795), .B2(G311), .ZN(new_n1082));
  INV_X1    g0882(.A(G322), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n1082), .B1(new_n1083), .B2(new_n800), .C1(new_n798), .C2(new_n1043), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT48), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n1044), .A2(new_n785), .B1(new_n778), .B2(new_n527), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1086), .A2(KEYINPUT49), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n815), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G116), .A2(new_n873), .B1(new_n783), .B2(G326), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(KEYINPUT49), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1081), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1072), .B(new_n1073), .C1(new_n774), .C2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n1003), .B2(new_n769), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n765), .A2(new_n1003), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n715), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n765), .A2(new_n1003), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1096), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(KEYINPUT117), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT117), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1102), .B(new_n1096), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n1103), .ZN(G393));
  OAI21_X1  g0904(.A(new_n824), .B1(new_n400), .B2(new_n210), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n247), .B2(new_n816), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G311), .A2(new_n799), .B1(new_n801), .B2(G317), .ZN(new_n1107));
  XOR2_X1   g0907(.A(new_n1107), .B(KEYINPUT52), .Z(new_n1108));
  OAI21_X1  g0908(.A(new_n255), .B1(new_n786), .B2(new_n460), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n778), .A2(new_n785), .B1(new_n782), .B2(new_n1083), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1109), .B(new_n1110), .C1(G116), .C2(new_n789), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(G294), .A2(new_n792), .B1(new_n795), .B2(G303), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1108), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n869), .A2(new_n800), .B1(new_n798), .B2(new_n808), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT51), .Z(new_n1115));
  OAI22_X1  g0915(.A1(new_n778), .A2(new_n201), .B1(new_n786), .B2(new_n632), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(G143), .B2(new_n783), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n202), .B2(new_n1044), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n291), .A2(new_n794), .B1(new_n791), .B2(new_n296), .ZN(new_n1119));
  OR3_X1    g0919(.A1(new_n1118), .A2(new_n1090), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1113), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n773), .B(new_n1106), .C1(new_n1121), .C2(new_n774), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n986), .B2(new_n826), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n992), .A2(new_n996), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1123), .B1(new_n1124), .B2(new_n768), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1004), .A2(new_n715), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1124), .A2(new_n1097), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(G390));
  AOI21_X1  g0929(.A(new_n898), .B1(new_n763), .B2(new_n835), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n937), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n957), .B(new_n947), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n748), .A2(new_n884), .A3(new_n937), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n956), .B1(new_n902), .B2(new_n937), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT110), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n965), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(KEYINPUT39), .B1(new_n923), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n966), .A2(new_n1135), .A3(new_n949), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1132), .B(new_n1133), .C1(new_n1134), .C2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n947), .A2(new_n957), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n898), .B1(new_n846), .B2(new_n847), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n957), .B1(new_n1144), .B2(new_n1131), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1143), .B1(new_n1145), .B2(new_n955), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n969), .A2(G330), .A3(new_n963), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1140), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n723), .A2(new_n738), .ZN(new_n1149));
  OAI211_X1 g0949(.A(G330), .B(new_n884), .C1(new_n1149), .C2(new_n746), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n1131), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n1147), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n902), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n963), .A2(G330), .A3(new_n884), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n1131), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1133), .A2(new_n1130), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n473), .A2(G330), .A3(new_n963), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n959), .A2(new_n690), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1148), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1159), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1140), .B(new_n1163), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1162), .A2(new_n715), .A3(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n770), .B1(new_n857), .B2(new_n1079), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n499), .A2(new_n798), .B1(new_n800), .B2(new_n785), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G107), .B2(new_n795), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n786), .A2(new_n201), .B1(new_n782), .B2(new_n527), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT118), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n255), .B1(new_n778), .B2(new_n632), .C1(new_n1044), .C2(new_n202), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G97), .B2(new_n792), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1168), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n778), .A2(new_n869), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT53), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n1174), .A2(new_n1175), .B1(new_n1044), .B2(new_n808), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n1175), .B2(new_n1174), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(KEYINPUT54), .B(G143), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(G132), .A2(new_n799), .B1(new_n792), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(G125), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n256), .B1(new_n782), .B2(new_n1181), .C1(new_n291), .C2(new_n786), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(G128), .B2(new_n801), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n795), .A2(G137), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1177), .A2(new_n1180), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1173), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1166), .B1(new_n1186), .B2(new_n774), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n1139), .B2(new_n822), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT119), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1188), .B(new_n1189), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1140), .B(new_n769), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1191));
  AND2_X1   g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1165), .A2(new_n1192), .ZN(G378));
  AND2_X1   g0993(.A1(new_n1164), .A2(new_n1160), .ZN(new_n1194));
  XOR2_X1   g0994(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n306), .A2(new_n912), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT55), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n313), .A2(new_n321), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1198), .B1(new_n313), .B2(new_n321), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1196), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1198), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n322), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n313), .A2(new_n321), .A3(new_n1198), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1203), .A2(new_n1195), .A3(new_n1204), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1201), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n971), .B2(G330), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n721), .B(new_n1206), .C1(new_n967), .C2(new_n970), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n958), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n947), .A2(new_n969), .A3(new_n963), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n937), .A2(new_n884), .A3(new_n963), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(KEYINPUT40), .A2(new_n1211), .B1(new_n1212), .B2(new_n968), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1206), .B1(new_n1213), .B2(new_n721), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n971), .A2(G330), .A3(new_n1207), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1139), .A2(new_n956), .B1(new_n394), .B2(new_n695), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1214), .A2(new_n938), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1210), .A2(new_n1217), .A3(KEYINPUT57), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n715), .B1(new_n1194), .B2(new_n1218), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1210), .A2(new_n1217), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1164), .A2(new_n1160), .ZN(new_n1221));
  AOI21_X1  g1021(.A(KEYINPUT57), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1219), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1210), .A2(new_n1217), .A3(new_n769), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n770), .B1(new_n857), .B2(G50), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n269), .B1(new_n778), .B2(new_n202), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n786), .A2(new_n292), .B1(new_n782), .B2(new_n785), .ZN(new_n1227));
  NOR4_X1   g1027(.A1(new_n815), .A2(new_n1052), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(G97), .A2(new_n795), .B1(new_n799), .B2(G107), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(G116), .A2(new_n801), .B1(new_n792), .B2(new_n641), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1231), .B(KEYINPUT58), .ZN(new_n1232));
  AOI21_X1  g1032(.A(G41), .B1(new_n815), .B2(G33), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n1044), .A2(new_n869), .B1(new_n1178), .B2(new_n778), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(G125), .A2(new_n801), .B1(new_n799), .B2(G128), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n868), .B2(new_n791), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n1234), .B(new_n1236), .C1(G132), .C2(new_n795), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1238), .A2(KEYINPUT59), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n251), .B(new_n269), .C1(new_n786), .C2(new_n808), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G124), .B2(new_n783), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT59), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1241), .B1(new_n1237), .B2(new_n1242), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n1232), .B1(G50), .B2(new_n1233), .C1(new_n1239), .C2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1225), .B1(new_n1244), .B2(new_n774), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1245), .B1(new_n1206), .B2(new_n822), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1224), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1223), .A2(new_n1247), .ZN(G375));
  NAND2_X1  g1048(.A1(new_n1131), .A2(new_n821), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n770), .B1(new_n857), .B2(G68), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(G283), .A2(new_n799), .B1(new_n801), .B2(G294), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(G107), .A2(new_n792), .B1(new_n795), .B2(G116), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n255), .B1(new_n786), .B2(new_n202), .ZN(new_n1253));
  INV_X1    g1053(.A(G303), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n778), .A2(new_n400), .B1(new_n782), .B2(new_n1254), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1074), .A2(new_n1253), .A3(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1251), .A2(new_n1252), .A3(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n815), .B1(new_n292), .B2(new_n786), .ZN(new_n1258));
  XOR2_X1   g1058(.A(new_n1258), .B(KEYINPUT121), .Z(new_n1259));
  AOI22_X1  g1059(.A1(G159), .A2(new_n779), .B1(new_n783), .B2(G128), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n291), .B2(new_n1044), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(new_n795), .B2(new_n1179), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(G132), .A2(new_n801), .B1(new_n792), .B2(G150), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1262), .B(new_n1263), .C1(new_n868), .C2(new_n798), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1257), .B1(new_n1259), .B2(new_n1264), .ZN(new_n1265));
  OR2_X1    g1065(.A1(new_n1265), .A2(KEYINPUT122), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n775), .B1(new_n1265), .B2(KEYINPUT122), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1250), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1157), .A2(new_n769), .B1(new_n1249), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1161), .A2(new_n1007), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1269), .B1(new_n1270), .B2(new_n1271), .ZN(G381));
  INV_X1    g1072(.A(G375), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1060), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1165), .A2(new_n1192), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1101), .A2(new_n828), .A3(new_n1103), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NOR3_X1   g1077(.A1(G390), .A2(G381), .A3(G384), .ZN(new_n1278));
  AND4_X1   g1078(.A1(new_n1274), .A2(new_n1275), .A3(new_n1277), .A4(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1273), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT123), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1280), .B(new_n1281), .ZN(G407));
  NAND2_X1  g1082(.A1(new_n1275), .A2(new_n696), .ZN(new_n1283));
  OAI211_X1 g1083(.A(G407), .B(G213), .C1(G375), .C2(new_n1283), .ZN(G409));
  INV_X1    g1084(.A(KEYINPUT61), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n696), .A2(G213), .ZN(new_n1286));
  OAI211_X1 g1086(.A(G378), .B(new_n1247), .C1(new_n1219), .C2(new_n1222), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1220), .A2(new_n1221), .A3(new_n1007), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1247), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1275), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1286), .B1(new_n1287), .B2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1286), .A2(G2897), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1153), .A2(new_n1156), .A3(new_n1159), .A4(KEYINPUT60), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n715), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1161), .A2(KEYINPUT60), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1296), .B1(new_n1297), .B2(new_n1271), .ZN(new_n1298));
  AOI21_X1  g1098(.A(G384), .B1(new_n1298), .B2(new_n1269), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1271), .B1(KEYINPUT60), .B2(new_n1161), .ZN(new_n1300));
  OAI211_X1 g1100(.A(G384), .B(new_n1269), .C1(new_n1300), .C2(new_n1295), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1293), .B1(new_n1299), .B2(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1269), .B1(new_n1300), .B2(new_n1295), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1304), .A2(new_n855), .A3(new_n885), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1305), .A2(new_n1301), .A3(new_n1292), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1303), .A2(new_n1306), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1285), .B1(new_n1291), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(KEYINPUT127), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT127), .ZN(new_n1310));
  OAI211_X1 g1110(.A(new_n1310), .B(new_n1285), .C1(new_n1291), .C2(new_n1307), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1299), .A2(new_n1302), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1291), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(KEYINPUT62), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT62), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1291), .A2(new_n1315), .A3(new_n1312), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1309), .A2(new_n1311), .A3(new_n1314), .A4(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(KEYINPUT125), .B1(new_n1274), .B2(G390), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n828), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1277), .A2(new_n1319), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1274), .A2(G390), .ZN(new_n1321));
  AOI211_X1 g1121(.A(new_n1060), .B(new_n1128), .C1(new_n1031), .C2(new_n1034), .ZN(new_n1322));
  OAI22_X1  g1122(.A1(new_n1318), .A2(new_n1320), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(G387), .A2(new_n1128), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1320), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1274), .A2(G390), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1324), .A2(new_n1325), .A3(KEYINPUT125), .A4(new_n1326), .ZN(new_n1327));
  AND2_X1   g1127(.A1(new_n1323), .A2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1317), .A2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1291), .A2(KEYINPUT63), .A3(new_n1312), .ZN(new_n1330));
  XNOR2_X1  g1130(.A(new_n1330), .B(KEYINPUT126), .ZN(new_n1331));
  XOR2_X1   g1131(.A(KEYINPUT124), .B(KEYINPUT63), .Z(new_n1332));
  AOI21_X1  g1132(.A(new_n1332), .B1(new_n1291), .B2(new_n1312), .ZN(new_n1333));
  NOR3_X1   g1133(.A1(new_n1308), .A2(new_n1333), .A3(new_n1328), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1331), .A2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1329), .A2(new_n1335), .ZN(G405));
  NAND2_X1  g1136(.A1(G375), .A2(new_n1275), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(new_n1287), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1338), .A2(new_n1312), .ZN(new_n1339));
  OAI211_X1 g1139(.A(new_n1337), .B(new_n1287), .C1(new_n1299), .C2(new_n1302), .ZN(new_n1340));
  AND3_X1   g1140(.A1(new_n1339), .A2(new_n1328), .A3(new_n1340), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1328), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1341), .A2(new_n1342), .ZN(G402));
endmodule


