//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 1 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991;
  AND2_X1   g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT75), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G155gat), .ZN(new_n205));
  INV_X1    g004(.A(G162gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT75), .ZN(new_n208));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  AND2_X1   g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n209), .A2(KEYINPUT2), .ZN(new_n214));
  NAND4_X1  g013(.A1(new_n204), .A2(new_n210), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G141gat), .B(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(KEYINPUT74), .A2(KEYINPUT2), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT74), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT2), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n218), .A2(new_n219), .B1(G155gat), .B2(G162gat), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n216), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT73), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n222), .B1(new_n202), .B2(new_n203), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n207), .A2(KEYINPUT73), .A3(new_n209), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n215), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT3), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n218), .A2(new_n219), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n228), .A2(new_n217), .A3(new_n209), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(new_n213), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n230), .A2(new_n223), .A3(new_n224), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT3), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(new_n232), .A3(new_n215), .ZN(new_n233));
  XNOR2_X1  g032(.A(G113gat), .B(G120gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G127gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n237), .A2(G134gat), .ZN(new_n238));
  INV_X1    g037(.A(G134gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n239), .A2(G127gat), .ZN(new_n240));
  OAI22_X1  g039(.A1(new_n234), .A2(new_n236), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G120gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G113gat), .ZN(new_n243));
  INV_X1    g042(.A(G113gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G120gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G127gat), .B(G134gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(new_n247), .A3(new_n235), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n241), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n227), .A2(new_n233), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G225gat), .A2(G233gat), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n252), .B1(new_n226), .B2(new_n249), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n241), .A2(new_n248), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n254), .A2(KEYINPUT4), .A3(new_n231), .A4(new_n215), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n250), .A2(new_n251), .A3(new_n253), .A4(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT5), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n254), .A2(new_n231), .A3(new_n215), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n226), .A2(new_n249), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n251), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n257), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n256), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT76), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(new_n266), .A3(new_n257), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT76), .B1(new_n256), .B2(KEYINPUT5), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n264), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(G1gat), .B(G29gat), .Z(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT0), .ZN(new_n271));
  XNOR2_X1  g070(.A(G57gat), .B(G85gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT6), .B1(new_n269), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n268), .ZN(new_n275));
  NOR3_X1   g074(.A1(new_n256), .A2(KEYINPUT76), .A3(KEYINPUT5), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n263), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n273), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n277), .A2(KEYINPUT6), .A3(new_n278), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G197gat), .B(G204gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT22), .ZN(new_n285));
  INV_X1    g084(.A(G211gat), .ZN(new_n286));
  INV_X1    g085(.A(G218gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G211gat), .B(G218gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n290), .A2(new_n284), .A3(new_n288), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G226gat), .A2(G233gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT25), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT24), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n299), .A2(G183gat), .A3(G190gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(G183gat), .B(G190gat), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n300), .B1(new_n301), .B2(new_n299), .ZN(new_n302));
  INV_X1    g101(.A(G169gat), .ZN(new_n303));
  INV_X1    g102(.A(G176gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n303), .A2(new_n304), .A3(KEYINPUT23), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT23), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(G169gat), .B2(G176gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n298), .B1(new_n302), .B2(new_n309), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n305), .A2(new_n307), .A3(KEYINPUT25), .A4(new_n308), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT64), .B1(new_n302), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n311), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n299), .A2(G183gat), .A3(G190gat), .ZN(new_n314));
  INV_X1    g113(.A(G183gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G190gat), .ZN(new_n316));
  INV_X1    g115(.A(G190gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G183gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n314), .B1(new_n319), .B2(KEYINPUT24), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT64), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n313), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n310), .A2(new_n312), .A3(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(G169gat), .A2(G176gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n324), .A2(KEYINPUT26), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n308), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n324), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT27), .B(G183gat), .ZN(new_n328));
  AND3_X1   g127(.A1(new_n328), .A2(KEYINPUT28), .A3(new_n317), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT28), .B1(new_n328), .B2(new_n317), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n326), .B(new_n327), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n323), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT29), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n297), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n296), .B1(new_n323), .B2(new_n331), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n295), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G8gat), .B(G36gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(G64gat), .B(G92gat), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n337), .B(new_n338), .Z(new_n339));
  NAND2_X1  g138(.A1(new_n332), .A2(new_n297), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT29), .B1(new_n323), .B2(new_n331), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n340), .B(new_n294), .C1(new_n297), .C2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n336), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT30), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n336), .A2(new_n342), .ZN(new_n346));
  INV_X1    g145(.A(new_n339), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n336), .A2(KEYINPUT30), .A3(new_n342), .A4(new_n339), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n345), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NOR3_X1   g149(.A1(new_n283), .A2(KEYINPUT35), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n323), .A2(new_n254), .A3(new_n331), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT66), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n332), .A2(new_n249), .ZN(new_n355));
  NAND2_X1  g154(.A1(G227gat), .A2(G233gat), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n323), .A2(KEYINPUT66), .A3(new_n254), .A4(new_n331), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n354), .A2(new_n355), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n254), .B1(new_n323), .B2(new_n331), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n361), .B1(new_n353), .B2(new_n352), .ZN(new_n362));
  NAND2_X1  g161(.A1(KEYINPUT69), .A2(KEYINPUT34), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n362), .A2(new_n356), .A3(new_n357), .A4(new_n363), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT32), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n354), .A2(new_n357), .A3(new_n355), .ZN(new_n367));
  INV_X1    g166(.A(new_n356), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT33), .B1(new_n367), .B2(new_n368), .ZN(new_n370));
  XNOR2_X1  g169(.A(G15gat), .B(G43gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(G71gat), .B(G99gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n369), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n367), .A2(new_n368), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT32), .ZN(new_n376));
  INV_X1    g175(.A(new_n373), .ZN(new_n377));
  AND2_X1   g176(.A1(new_n377), .A2(KEYINPUT67), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT33), .B1(new_n377), .B2(KEYINPUT67), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n365), .B1(new_n374), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT33), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n375), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n376), .A2(new_n384), .A3(new_n377), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n369), .B1(new_n378), .B2(new_n379), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n360), .A2(new_n364), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  AND2_X1   g187(.A1(new_n382), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(KEYINPUT31), .B(G50gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(G228gat), .A2(G233gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n294), .A2(new_n333), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT3), .B1(new_n392), .B2(KEYINPUT77), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n392), .A2(KEYINPUT77), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n226), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n294), .B1(new_n233), .B2(new_n333), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n391), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n226), .A2(new_n333), .A3(new_n294), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n400), .A2(new_n227), .A3(new_n391), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n401), .A2(new_n397), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n390), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G78gat), .B(G106gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(G22gat), .ZN(new_n405));
  INV_X1    g204(.A(new_n402), .ZN(new_n406));
  INV_X1    g205(.A(new_n390), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n393), .B1(KEYINPUT77), .B2(new_n392), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n397), .B1(new_n408), .B2(new_n226), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n406), .B(new_n407), .C1(new_n409), .C2(new_n391), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n403), .A2(new_n405), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n405), .B1(new_n403), .B2(new_n410), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n389), .A2(new_n414), .ZN(new_n415));
  OAI22_X1  g214(.A1(new_n374), .A2(new_n381), .B1(KEYINPUT68), .B2(new_n365), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT68), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n385), .A2(new_n417), .A3(new_n386), .A4(new_n387), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT72), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n348), .A2(new_n420), .A3(new_n349), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n345), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n420), .B1(new_n348), .B2(new_n349), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n419), .A2(new_n282), .A3(new_n424), .A4(new_n413), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n351), .A2(new_n415), .B1(KEYINPUT35), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  XOR2_X1   g226(.A(KEYINPUT70), .B(KEYINPUT36), .Z(new_n428));
  NAND3_X1  g227(.A1(new_n382), .A2(new_n428), .A3(new_n388), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT71), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n419), .A2(KEYINPUT36), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT71), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n382), .A2(new_n432), .A3(new_n388), .A4(new_n428), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n430), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT40), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT39), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n231), .A2(new_n232), .A3(new_n215), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n232), .B1(new_n231), .B2(new_n215), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n437), .A2(new_n438), .A3(new_n254), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n253), .A2(new_n255), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n436), .B(new_n261), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n273), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n258), .A2(new_n259), .A3(new_n251), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT39), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n250), .A2(new_n253), .A3(new_n255), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n444), .B1(new_n445), .B2(new_n261), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n435), .B1(new_n442), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT78), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT78), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n449), .B(new_n435), .C1(new_n442), .C2(new_n446), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n261), .B1(new_n439), .B2(new_n440), .ZN(new_n452));
  INV_X1    g251(.A(new_n444), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n454), .A2(KEYINPUT40), .A3(new_n273), .A4(new_n441), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT79), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n441), .A2(new_n273), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n458), .A2(KEYINPUT79), .A3(KEYINPUT40), .A4(new_n454), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n451), .A2(new_n460), .A3(new_n279), .A4(new_n350), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT38), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT37), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n336), .A2(new_n463), .A3(new_n342), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n346), .A2(KEYINPUT37), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n347), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT80), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI211_X1 g268(.A(new_n468), .B(new_n339), .C1(new_n346), .C2(KEYINPUT37), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n462), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n343), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n464), .A2(new_n462), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n339), .B1(new_n346), .B2(KEYINPUT37), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n280), .A2(new_n281), .A3(new_n476), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n413), .B(new_n461), .C1(new_n472), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n282), .A2(new_n424), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n414), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n434), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n427), .A2(new_n481), .ZN(new_n482));
  XOR2_X1   g281(.A(G43gat), .B(G50gat), .Z(new_n483));
  INV_X1    g282(.A(KEYINPUT15), .ZN(new_n484));
  OR2_X1    g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT14), .ZN(new_n486));
  INV_X1    g285(.A(G29gat), .ZN(new_n487));
  INV_X1    g286(.A(G36gat), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT81), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT81), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n491), .A2(new_n486), .A3(new_n487), .A4(new_n488), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT82), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n495), .A2(new_n496), .B1(G29gat), .B2(G36gat), .ZN(new_n497));
  INV_X1    g296(.A(new_n494), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n498), .B1(new_n490), .B2(new_n492), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT82), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n485), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n484), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n502), .B(KEYINPUT83), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n489), .A2(new_n494), .ZN(new_n504));
  NAND2_X1  g303(.A1(G29gat), .A2(G36gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT84), .ZN(new_n506));
  OR2_X1    g305(.A1(new_n505), .A2(KEYINPUT84), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n485), .A2(new_n504), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT85), .B1(new_n501), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n485), .ZN(new_n511));
  INV_X1    g310(.A(new_n500), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n505), .B1(new_n499), .B2(KEYINPUT82), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT85), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n514), .B(new_n515), .C1(new_n503), .C2(new_n508), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G15gat), .B(G22gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT87), .ZN(new_n519));
  XOR2_X1   g318(.A(new_n519), .B(G8gat), .Z(new_n520));
  INV_X1    g319(.A(KEYINPUT16), .ZN(new_n521));
  AOI21_X1  g320(.A(G1gat), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n520), .B(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n517), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n510), .A2(new_n516), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT86), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n510), .A2(new_n516), .A3(KEYINPUT86), .A4(new_n525), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n501), .A2(new_n509), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT17), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n523), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n524), .B1(new_n530), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G229gat), .A2(G233gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT88), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n538), .A2(KEYINPUT18), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n536), .B(KEYINPUT13), .Z(new_n541));
  AND2_X1   g340(.A1(new_n517), .A2(new_n523), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n541), .B1(new_n542), .B2(new_n524), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n535), .B(new_n536), .C1(new_n538), .C2(KEYINPUT18), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n540), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G113gat), .B(G141gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(G197gat), .ZN(new_n547));
  XOR2_X1   g346(.A(KEYINPUT11), .B(G169gat), .Z(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n549), .B(KEYINPUT12), .Z(new_n550));
  NAND2_X1  g349(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n550), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n540), .A2(new_n552), .A3(new_n544), .A4(new_n543), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n482), .A2(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n555), .B(KEYINPUT89), .Z(new_n556));
  NAND3_X1  g355(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT95), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT7), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT96), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n560), .A2(G85gat), .A3(G92gat), .ZN(new_n561));
  MUX2_X1   g360(.A(new_n559), .B(KEYINPUT7), .S(new_n561), .Z(new_n562));
  XNOR2_X1  g361(.A(G99gat), .B(G106gat), .ZN(new_n563));
  INV_X1    g362(.A(G99gat), .ZN(new_n564));
  INV_X1    g363(.A(G106gat), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT8), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(G85gat), .ZN(new_n567));
  INV_X1    g366(.A(G92gat), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT95), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n568), .ZN(new_n570));
  AND3_X1   g369(.A1(new_n566), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n562), .A2(new_n563), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n563), .B1(new_n562), .B2(new_n571), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n557), .B1(new_n517), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n574), .B1(new_n531), .B2(KEYINPUT17), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n576), .B1(new_n530), .B2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G190gat), .B(G218gat), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(new_n580), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G134gat), .B(G162gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT94), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n585), .B(new_n586), .Z(new_n587));
  NOR2_X1   g386(.A1(new_n578), .A2(new_n580), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT97), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n583), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n581), .A2(new_n589), .A3(new_n582), .A4(new_n587), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT21), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT90), .ZN(new_n595));
  XNOR2_X1  g394(.A(G57gat), .B(G64gat), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AND2_X1   g397(.A1(G71gat), .A2(G78gat), .ZN(new_n599));
  NOR2_X1   g398(.A1(G71gat), .A2(G78gat), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  OAI221_X1 g401(.A(new_n595), .B1(new_n599), .B2(new_n600), .C1(new_n596), .C2(new_n597), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT92), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n523), .B1(new_n594), .B2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT93), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT91), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(G155gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n608), .B(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n604), .A2(KEYINPUT21), .ZN(new_n613));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(new_n237), .ZN(new_n616));
  XOR2_X1   g415(.A(G183gat), .B(G211gat), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n612), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n612), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n593), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT98), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n604), .B1(new_n572), .B2(new_n573), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n562), .A2(new_n571), .ZN(new_n625));
  INV_X1    g424(.A(new_n563), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n604), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n562), .A2(new_n563), .A3(new_n571), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(KEYINPUT10), .B1(new_n624), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n627), .A2(KEYINPUT10), .A3(new_n629), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n606), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G230gat), .A2(G233gat), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n623), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  OAI211_X1 g436(.A(KEYINPUT98), .B(new_n635), .C1(new_n631), .C2(new_n633), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G120gat), .B(G148gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(G176gat), .B(G204gat), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n640), .B(new_n641), .Z(new_n642));
  NAND2_X1  g441(.A1(new_n624), .A2(new_n630), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n639), .B(new_n642), .C1(new_n635), .C2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n642), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n635), .B(KEYINPUT99), .Z(new_n646));
  NOR2_X1   g445(.A1(new_n634), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n643), .A2(new_n635), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n622), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n556), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n283), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n350), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n658), .A2(G8gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(KEYINPUT16), .B(G8gat), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT42), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(KEYINPUT42), .B2(new_n661), .ZN(G1325gat));
  OAI21_X1  g462(.A(G15gat), .B1(new_n654), .B2(new_n434), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n389), .A2(G15gat), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n664), .B1(new_n654), .B2(new_n665), .ZN(G1326gat));
  NOR2_X1   g465(.A1(new_n654), .A2(new_n413), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT43), .B(G22gat), .Z(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  AND4_X1   g468(.A1(new_n556), .A2(new_n593), .A3(new_n621), .A4(new_n651), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n670), .A2(new_n487), .A3(new_n283), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT45), .ZN(new_n672));
  AND4_X1   g471(.A1(KEYINPUT101), .A2(new_n434), .A3(new_n478), .A4(new_n480), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n464), .B1(new_n475), .B2(KEYINPUT80), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT38), .B1(new_n674), .B2(new_n470), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n675), .A2(new_n281), .A3(new_n280), .A4(new_n476), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n461), .A2(new_n413), .ZN(new_n677));
  AOI22_X1  g476(.A1(new_n676), .A2(new_n677), .B1(new_n479), .B2(new_n414), .ZN(new_n678));
  AOI21_X1  g477(.A(KEYINPUT101), .B1(new_n678), .B2(new_n434), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n427), .B1(new_n673), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT102), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT101), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n481), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n678), .A2(KEYINPUT101), .A3(new_n434), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n426), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n591), .A2(new_n592), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n688), .A2(KEYINPUT44), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n681), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n482), .A2(new_n593), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT44), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n554), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n650), .B(KEYINPUT100), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n621), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n694), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n693), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(G29gat), .B1(new_n699), .B2(new_n282), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n672), .A2(new_n700), .ZN(G1328gat));
  NAND3_X1  g500(.A1(new_n670), .A2(new_n488), .A3(new_n350), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT46), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n703), .A2(KEYINPUT103), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n703), .A2(KEYINPUT103), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n702), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n350), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n699), .A2(new_n707), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n708), .A2(KEYINPUT104), .ZN(new_n709));
  OAI21_X1  g508(.A(G36gat), .B1(new_n708), .B2(KEYINPUT104), .ZN(new_n710));
  OAI221_X1 g509(.A(new_n706), .B1(new_n704), .B2(new_n702), .C1(new_n709), .C2(new_n710), .ZN(G1329gat));
  INV_X1    g510(.A(G43gat), .ZN(new_n712));
  INV_X1    g511(.A(new_n389), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n670), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT47), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n699), .A2(KEYINPUT105), .A3(new_n434), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n699), .A2(new_n434), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n719));
  OAI21_X1  g518(.A(G43gat), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n716), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n718), .A2(new_n712), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n715), .B1(new_n714), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(G1330gat));
  NOR2_X1   g523(.A1(new_n413), .A2(G50gat), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n693), .A2(new_n414), .A3(new_n698), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n670), .A2(new_n725), .B1(G50gat), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g527(.A1(new_n685), .A2(new_n686), .ZN(new_n729));
  AOI211_X1 g528(.A(KEYINPUT102), .B(new_n426), .C1(new_n683), .C2(new_n684), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR4_X1   g530(.A1(new_n593), .A2(new_n554), .A3(new_n621), .A4(new_n695), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n733), .A2(new_n282), .ZN(new_n734));
  XOR2_X1   g533(.A(KEYINPUT106), .B(G57gat), .Z(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1332gat));
  INV_X1    g535(.A(new_n733), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n707), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT107), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n740), .B(new_n741), .Z(G1333gat));
  INV_X1    g541(.A(G71gat), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n733), .A2(new_n743), .A3(new_n434), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT108), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n743), .B1(new_n733), .B2(new_n389), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g547(.A1(new_n737), .A2(new_n414), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G78gat), .ZN(G1335gat));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(new_n685), .B2(new_n688), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n680), .A2(KEYINPUT110), .A3(new_n593), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n554), .A2(new_n697), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT109), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n752), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n752), .A2(new_n753), .A3(KEYINPUT51), .A4(new_n755), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n760), .A2(new_n567), .A3(new_n283), .A4(new_n650), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n755), .A2(new_n650), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n762), .B1(new_n690), .B2(new_n692), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(G85gat), .B1(new_n764), .B2(new_n282), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n761), .A2(new_n765), .ZN(G1336gat));
  AOI21_X1  g565(.A(new_n568), .B1(new_n763), .B2(new_n350), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n695), .A2(G92gat), .A3(new_n707), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n769), .B1(new_n758), .B2(new_n759), .ZN(new_n770));
  OAI21_X1  g569(.A(KEYINPUT52), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT111), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n773), .B(KEYINPUT52), .C1(new_n767), .C2(new_n770), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n762), .ZN(new_n776));
  INV_X1    g575(.A(new_n689), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n729), .A2(new_n730), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n692), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n350), .B(new_n776), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G92gat), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n754), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n683), .A2(new_n684), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n688), .B1(new_n784), .B2(new_n427), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n783), .B1(new_n785), .B2(KEYINPUT110), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT51), .B1(new_n786), .B2(new_n752), .ZN(new_n787));
  AND4_X1   g586(.A1(KEYINPUT51), .A2(new_n752), .A3(new_n753), .A4(new_n755), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n768), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n781), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT112), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n781), .A2(new_n789), .A3(new_n793), .A4(new_n790), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n775), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT113), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n775), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(G1337gat));
  NAND4_X1  g599(.A1(new_n760), .A2(new_n564), .A3(new_n713), .A4(new_n650), .ZN(new_n801));
  OAI21_X1  g600(.A(G99gat), .B1(new_n764), .B2(new_n434), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(G1338gat));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n804));
  OAI21_X1  g603(.A(G106gat), .B1(new_n764), .B2(new_n413), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n760), .A2(new_n565), .A3(new_n414), .A4(new_n696), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n805), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n807), .B(new_n809), .ZN(G1339gat));
  NOR2_X1   g609(.A1(new_n652), .A2(new_n554), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  XNOR2_X1  g611(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n642), .B1(new_n647), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n816), .B1(new_n634), .B2(new_n646), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT10), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n643), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n604), .B(KEYINPUT92), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(new_n574), .A3(KEYINPUT10), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT98), .B1(new_n822), .B2(new_n635), .ZN(new_n823));
  INV_X1    g622(.A(new_n638), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n817), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT115), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI211_X1 g626(.A(KEYINPUT115), .B(new_n817), .C1(new_n823), .C2(new_n824), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n815), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n644), .B1(new_n829), .B2(KEYINPUT55), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n831));
  AOI211_X1 g630(.A(new_n831), .B(new_n815), .C1(new_n827), .C2(new_n828), .ZN(new_n832));
  OAI21_X1  g631(.A(KEYINPUT117), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n834), .B1(new_n535), .B2(new_n536), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n542), .A2(new_n524), .ZN(new_n836));
  INV_X1    g635(.A(new_n541), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n536), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n533), .B1(new_n528), .B2(new_n529), .ZN(new_n840));
  OAI211_X1 g639(.A(KEYINPUT118), .B(new_n839), .C1(new_n840), .C2(new_n524), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n835), .A2(new_n838), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n549), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n843), .A2(new_n553), .ZN(new_n844));
  INV_X1    g643(.A(new_n828), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT115), .B1(new_n639), .B2(new_n817), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n814), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n831), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n829), .A2(KEYINPUT55), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n848), .A2(new_n849), .A3(new_n850), .A4(new_n644), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n833), .A2(new_n593), .A3(new_n844), .A4(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AND4_X1   g653(.A1(new_n553), .A2(new_n591), .A3(new_n843), .A4(new_n592), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n855), .A2(KEYINPUT119), .A3(new_n833), .A4(new_n851), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n833), .A2(new_n554), .A3(new_n851), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n844), .A2(new_n650), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI22_X1  g658(.A1(new_n854), .A2(new_n856), .B1(new_n859), .B2(new_n688), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n812), .B1(new_n860), .B2(new_n697), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n861), .A2(new_n415), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n282), .A2(new_n350), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(G113gat), .B1(new_n864), .B2(new_n694), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n419), .A2(new_n413), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n861), .A2(new_n283), .A3(new_n707), .A4(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(new_n244), .A3(new_n554), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g670(.A(new_n871), .B(KEYINPUT120), .Z(G1340gat));
  NOR3_X1   g671(.A1(new_n864), .A2(new_n242), .A3(new_n695), .ZN(new_n873));
  AOI21_X1  g672(.A(G120gat), .B1(new_n869), .B2(new_n650), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(G1341gat));
  OAI21_X1  g674(.A(G127gat), .B1(new_n864), .B2(new_n621), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n869), .A2(new_n237), .A3(new_n697), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1342gat));
  NAND3_X1  g677(.A1(new_n869), .A2(new_n239), .A3(new_n593), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n879), .A2(KEYINPUT56), .ZN(new_n880));
  OAI21_X1  g679(.A(G134gat), .B1(new_n864), .B2(new_n688), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(KEYINPUT56), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(G1343gat));
  AND2_X1   g682(.A1(new_n434), .A2(new_n863), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT57), .B1(new_n861), .B2(new_n414), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n414), .A2(KEYINPUT57), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n854), .A2(new_n856), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n848), .A2(new_n849), .A3(new_n644), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n858), .B1(new_n694), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n688), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n621), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n886), .B1(new_n892), .B2(new_n812), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n554), .B(new_n884), .C1(new_n885), .C2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(G141gat), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n434), .A2(new_n414), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n896), .A2(new_n707), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n861), .A2(new_n283), .A3(new_n897), .ZN(new_n898));
  OR2_X1    g697(.A1(new_n694), .A2(G141gat), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n895), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(KEYINPUT122), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n904), .B1(new_n894), .B2(G141gat), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT58), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT122), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n895), .A2(new_n908), .A3(new_n901), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n903), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n908), .B1(new_n895), .B2(new_n901), .ZN(new_n911));
  AOI211_X1 g710(.A(KEYINPUT122), .B(new_n900), .C1(new_n894), .C2(G141gat), .ZN(new_n912));
  OAI22_X1  g711(.A1(new_n911), .A2(new_n912), .B1(new_n906), .B2(new_n905), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n910), .A2(new_n913), .ZN(G1344gat));
  INV_X1    g713(.A(KEYINPUT124), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n811), .B(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n855), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n890), .B1(new_n917), .B2(new_n888), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n621), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n413), .B1(new_n920), .B2(KEYINPUT125), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT125), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n916), .A2(new_n922), .A3(new_n919), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT57), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  AND3_X1   g723(.A1(new_n861), .A2(KEYINPUT57), .A3(new_n414), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n884), .A2(new_n650), .ZN(new_n927));
  OAI211_X1 g726(.A(KEYINPUT59), .B(G148gat), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n884), .B1(new_n885), .B2(new_n893), .ZN(new_n929));
  OAI21_X1  g728(.A(G148gat), .B1(new_n929), .B2(new_n651), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT59), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n898), .A2(G148gat), .A3(new_n651), .ZN(new_n933));
  XOR2_X1   g732(.A(new_n933), .B(KEYINPUT123), .Z(new_n934));
  NAND3_X1  g733(.A1(new_n928), .A2(new_n932), .A3(new_n934), .ZN(G1345gat));
  OAI21_X1  g734(.A(G155gat), .B1(new_n929), .B2(new_n621), .ZN(new_n936));
  INV_X1    g735(.A(new_n898), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n937), .A2(new_n205), .A3(new_n697), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1346gat));
  OAI21_X1  g738(.A(G162gat), .B1(new_n929), .B2(new_n688), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n937), .A2(new_n206), .A3(new_n593), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1347gat));
  NOR2_X1   g741(.A1(new_n283), .A2(new_n707), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n862), .A2(new_n943), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n944), .A2(new_n303), .A3(new_n694), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n861), .A2(new_n282), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n946), .A2(KEYINPUT126), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n707), .B1(new_n946), .B2(KEYINPUT126), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n949), .A2(new_n867), .A3(new_n554), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n945), .B1(new_n950), .B2(new_n303), .ZN(G1348gat));
  OAI21_X1  g750(.A(G176gat), .B1(new_n944), .B2(new_n695), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n949), .A2(new_n867), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n650), .A2(new_n304), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(G1349gat));
  NAND4_X1  g754(.A1(new_n949), .A2(new_n328), .A3(new_n867), .A4(new_n697), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n862), .A2(new_n697), .A3(new_n943), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n315), .B1(new_n957), .B2(KEYINPUT127), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n958), .B1(KEYINPUT127), .B2(new_n957), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(KEYINPUT60), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT60), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n956), .A2(new_n959), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n961), .A2(new_n963), .ZN(G1350gat));
  OAI21_X1  g763(.A(G190gat), .B1(new_n944), .B2(new_n688), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n965), .A2(KEYINPUT61), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n965), .A2(KEYINPUT61), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n593), .A2(new_n317), .ZN(new_n968));
  OAI22_X1  g767(.A1(new_n966), .A2(new_n967), .B1(new_n953), .B2(new_n968), .ZN(G1351gat));
  AND2_X1   g768(.A1(new_n949), .A2(new_n896), .ZN(new_n970));
  AOI21_X1  g769(.A(G197gat), .B1(new_n970), .B2(new_n554), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n434), .A2(new_n943), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n926), .A2(new_n972), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n554), .A2(G197gat), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n971), .B1(new_n973), .B2(new_n974), .ZN(G1352gat));
  NOR2_X1   g774(.A1(new_n651), .A2(G204gat), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n970), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(KEYINPUT62), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT62), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n970), .A2(new_n979), .A3(new_n976), .ZN(new_n980));
  INV_X1    g779(.A(new_n972), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n981), .B1(new_n924), .B2(new_n925), .ZN(new_n982));
  OAI21_X1  g781(.A(G204gat), .B1(new_n982), .B2(new_n695), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n978), .A2(new_n980), .A3(new_n983), .ZN(G1353gat));
  NAND3_X1  g783(.A1(new_n970), .A2(new_n286), .A3(new_n697), .ZN(new_n985));
  OAI211_X1 g784(.A(new_n697), .B(new_n981), .C1(new_n924), .C2(new_n925), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n986), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT63), .B1(new_n986), .B2(G211gat), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(G1354gat));
  NAND3_X1  g788(.A1(new_n970), .A2(new_n287), .A3(new_n593), .ZN(new_n990));
  OAI21_X1  g789(.A(G218gat), .B1(new_n982), .B2(new_n688), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(G1355gat));
endmodule


