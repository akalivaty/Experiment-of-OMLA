//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1302, new_n1303, new_n1304;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n211), .B(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(KEYINPUT65), .B(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G107), .A2(G264), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n209), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  AND2_X1   g0024(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR3_X1   g0027(.A1(new_n226), .A2(new_n207), .A3(new_n227), .ZN(new_n228));
  NOR4_X1   g0028(.A1(new_n213), .A2(new_n224), .A3(new_n225), .A4(new_n228), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT67), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G58), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  XNOR2_X1  g0046(.A(KEYINPUT3), .B(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n247), .A2(G222), .A3(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G77), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n247), .A2(G1698), .ZN(new_n251));
  INV_X1    g0051(.A(G223), .ZN(new_n252));
  OAI221_X1 g0052(.A(new_n249), .B1(new_n250), .B2(new_n247), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G1), .A3(G13), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT68), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT68), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G41), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  OAI211_X1 g0062(.A(KEYINPUT69), .B(new_n206), .C1(new_n262), .C2(G45), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT69), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n206), .A2(G45), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT68), .B(G41), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n264), .B(new_n265), .C1(new_n266), .C2(G1), .ZN(new_n267));
  INV_X1    g0067(.A(G274), .ZN(new_n268));
  INV_X1    g0068(.A(new_n227), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n268), .B1(new_n269), .B2(new_n254), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n263), .A2(new_n267), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G45), .ZN(new_n272));
  AOI21_X1  g0072(.A(G1), .B1(new_n258), .B2(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n256), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G226), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n257), .A2(new_n271), .A3(new_n275), .ZN(new_n276));
  OR2_X1    g0076(.A1(new_n276), .A2(G179), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n227), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G150), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n207), .A2(G33), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT70), .ZN(new_n283));
  XNOR2_X1  g0083(.A(new_n282), .B(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n281), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G58), .A2(G68), .ZN(new_n287));
  INV_X1    g0087(.A(G50), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n207), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT71), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n279), .B1(new_n286), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G13), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(G1), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G20), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(new_n279), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n288), .B1(new_n206), .B2(G20), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n296), .A2(new_n297), .B1(new_n288), .B2(new_n295), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n291), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n276), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n277), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n299), .B(KEYINPUT9), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n276), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  OR2_X1    g0107(.A1(new_n307), .A2(KEYINPUT76), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n276), .A2(G200), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT75), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n307), .A2(KEYINPUT76), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n308), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT10), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT74), .ZN(new_n314));
  OR2_X1    g0114(.A1(new_n304), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n304), .A2(new_n314), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT10), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n306), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n315), .A2(new_n310), .A3(new_n316), .A4(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n303), .B1(new_n313), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n296), .ZN(new_n321));
  INV_X1    g0121(.A(new_n285), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n206), .A2(G20), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n321), .A2(new_n324), .B1(new_n294), .B2(new_n322), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT7), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(new_n247), .B2(G20), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT3), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n328), .A2(G33), .ZN(new_n329));
  INV_X1    g0129(.A(G33), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(KEYINPUT3), .ZN(new_n331));
  OAI211_X1 g0131(.A(KEYINPUT7), .B(new_n207), .C1(new_n329), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G68), .ZN(new_n334));
  INV_X1    g0134(.A(G58), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n335), .A2(new_n215), .ZN(new_n336));
  OAI21_X1  g0136(.A(G20), .B1(new_n336), .B2(new_n287), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n280), .A2(G159), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n334), .A2(KEYINPUT16), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT16), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n215), .B1(new_n327), .B2(new_n332), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n342), .B1(new_n343), .B2(new_n339), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n341), .A2(new_n344), .A3(new_n279), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT78), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n341), .A2(new_n344), .A3(KEYINPUT78), .A4(new_n279), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n325), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(G33), .A2(G87), .ZN(new_n350));
  INV_X1    g0150(.A(G226), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n247), .A2(new_n248), .ZN(new_n352));
  OAI221_X1 g0152(.A(new_n350), .B1(new_n251), .B2(new_n351), .C1(new_n252), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n256), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n274), .A2(G232), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(new_n355), .A3(new_n271), .ZN(new_n356));
  INV_X1    g0156(.A(G200), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n271), .A2(new_n355), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT79), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n271), .A2(KEYINPUT79), .A3(new_n355), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n361), .A2(new_n305), .A3(new_n354), .A4(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n349), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT17), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n347), .A2(new_n348), .ZN(new_n368));
  INV_X1    g0168(.A(new_n325), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n356), .A2(new_n300), .ZN(new_n371));
  INV_X1    g0171(.A(G179), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n361), .A2(new_n372), .A3(new_n354), .A4(new_n362), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT18), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n370), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT18), .B1(new_n349), .B2(new_n374), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n349), .A2(KEYINPUT17), .A3(new_n364), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n367), .A2(new_n377), .A3(new_n378), .A4(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  OAI22_X1  g0181(.A1(new_n251), .A2(new_n214), .B1(new_n203), .B2(new_n247), .ZN(new_n382));
  AND3_X1   g0182(.A1(new_n247), .A2(G232), .A3(new_n248), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n256), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n274), .A2(G244), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(new_n271), .A3(new_n385), .ZN(new_n386));
  OR2_X1    g0186(.A1(new_n386), .A2(KEYINPUT72), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(KEYINPUT72), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G190), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n296), .A2(G77), .A3(new_n323), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT73), .B1(new_n295), .B2(new_n250), .ZN(new_n392));
  AND3_X1   g0192(.A1(new_n295), .A2(KEYINPUT73), .A3(new_n250), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n279), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n322), .A2(new_n280), .B1(G20), .B2(G77), .ZN(new_n396));
  XNOR2_X1  g0196(.A(KEYINPUT15), .B(G87), .ZN(new_n397));
  OR2_X1    g0197(.A1(new_n397), .A2(new_n282), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n395), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n394), .A2(new_n399), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n390), .B(new_n400), .C1(new_n357), .C2(new_n389), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n400), .B1(new_n389), .B2(new_n372), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n387), .A2(new_n300), .A3(new_n388), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n247), .A2(G232), .A3(G1698), .ZN(new_n407));
  NAND2_X1  g0207(.A1(G33), .A2(G97), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n407), .B(new_n408), .C1(new_n352), .C2(new_n351), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n256), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n274), .A2(G238), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n410), .A2(KEYINPUT13), .A3(new_n271), .A4(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n412), .A2(KEYINPUT77), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n410), .A2(new_n271), .A3(new_n411), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT13), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n415), .B1(KEYINPUT77), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n305), .B1(new_n414), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n415), .A2(new_n416), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n419), .A2(G200), .A3(new_n412), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n280), .A2(G50), .B1(G20), .B2(new_n215), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(new_n284), .B2(new_n250), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n422), .A2(KEYINPUT11), .A3(new_n279), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n296), .A2(G68), .A3(new_n323), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT12), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n295), .B2(new_n215), .ZN(new_n426));
  NOR3_X1   g0226(.A1(new_n294), .A2(KEYINPUT12), .A3(G68), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n423), .B(new_n424), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT11), .B1(new_n422), .B2(new_n279), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n420), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n418), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n417), .ZN(new_n433));
  OAI21_X1  g0233(.A(G179), .B1(new_n433), .B2(new_n413), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n419), .A2(G169), .A3(new_n412), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT14), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT14), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n419), .A2(new_n437), .A3(G169), .A4(new_n412), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n434), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n430), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n432), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n320), .A2(new_n381), .A3(new_n406), .A4(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n206), .A2(G33), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n395), .A2(new_n294), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(G116), .ZN(new_n446));
  XNOR2_X1  g0246(.A(KEYINPUT83), .B(G116), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  OAI22_X1  g0248(.A1(new_n445), .A2(new_n446), .B1(new_n294), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n447), .A2(G20), .ZN(new_n451));
  AOI21_X1  g0251(.A(G20), .B1(G33), .B2(G283), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n330), .A2(G97), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n452), .A2(new_n453), .B1(new_n278), .B2(new_n227), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT20), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n451), .A2(KEYINPUT20), .A3(new_n454), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n450), .B(KEYINPUT87), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT87), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n456), .A2(new_n455), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n458), .B1(new_n459), .B2(new_n449), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT5), .B1(new_n259), .B2(new_n261), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT5), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n206), .B(G45), .C1(new_n463), .C2(G41), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(new_n256), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G270), .ZN(new_n467));
  INV_X1    g0267(.A(new_n464), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n270), .B(new_n468), .C1(KEYINPUT5), .C2(new_n266), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n247), .A2(G264), .A3(G1698), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n330), .A2(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n328), .A2(G33), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G303), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G257), .ZN(new_n477));
  OAI21_X1  g0277(.A(KEYINPUT85), .B1(new_n352), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT85), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n247), .A2(new_n479), .A3(G257), .A4(new_n248), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n476), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n256), .B1(new_n481), .B2(KEYINPUT86), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT86), .ZN(new_n483));
  AOI211_X1 g0283(.A(new_n483), .B(new_n476), .C1(new_n480), .C2(new_n478), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n470), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n461), .A2(new_n485), .A3(new_n372), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n300), .B1(new_n457), .B2(new_n460), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n485), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT21), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT21), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n487), .A2(new_n485), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n486), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(G250), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n493), .B1(new_n272), .B2(G1), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n206), .A2(new_n268), .A3(G45), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n255), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT83), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(G116), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n446), .A2(KEYINPUT83), .ZN(new_n500));
  OAI21_X1  g0300(.A(G33), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n472), .A2(new_n473), .A3(G238), .A4(new_n248), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n472), .A2(new_n473), .A3(G244), .A4(G1698), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n497), .B1(new_n504), .B2(new_n256), .ZN(new_n505));
  OR2_X1    g0305(.A1(new_n505), .A2(new_n357), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n247), .A2(new_n207), .A3(G68), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT19), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n207), .B1(new_n408), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(G87), .B2(new_n204), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n508), .B1(new_n282), .B2(new_n202), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n507), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n512), .A2(new_n279), .B1(new_n295), .B2(new_n397), .ZN(new_n513));
  INV_X1    g0313(.A(new_n445), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G87), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n505), .A2(G190), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n506), .A2(new_n513), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT84), .ZN(new_n518));
  INV_X1    g0318(.A(new_n397), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n518), .B1(new_n514), .B2(new_n519), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n445), .A2(KEYINPUT84), .A3(new_n397), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n513), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI211_X1 g0322(.A(new_n372), .B(new_n497), .C1(new_n504), .C2(new_n256), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n504), .A2(new_n256), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n300), .B1(new_n524), .B2(new_n496), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n522), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n517), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n457), .A2(new_n460), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n485), .B2(G200), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n305), .B2(new_n485), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n492), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n295), .A2(new_n203), .ZN(new_n532));
  NOR2_X1   g0332(.A1(KEYINPUT90), .A2(KEYINPUT25), .ZN(new_n533));
  OR2_X1    g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g0334(.A1(KEYINPUT90), .A2(KEYINPUT25), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(new_n532), .B2(new_n533), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n534), .A2(new_n536), .B1(G107), .B2(new_n514), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n472), .A2(new_n473), .A3(new_n207), .A4(G87), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT22), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT22), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n247), .A2(new_n541), .A3(new_n207), .A4(G87), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n446), .A2(KEYINPUT83), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n498), .A2(G116), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n330), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT23), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n207), .B2(G107), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n203), .A2(KEYINPUT23), .A3(G20), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n546), .A2(new_n207), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT88), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n543), .A2(KEYINPUT88), .A3(new_n550), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(KEYINPUT24), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT88), .B1(new_n543), .B2(new_n550), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT24), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n395), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT89), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n555), .A2(KEYINPUT89), .A3(new_n558), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n538), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n466), .A2(G264), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n477), .A2(G1698), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(G250), .B2(G1698), .ZN(new_n566));
  INV_X1    g0366(.A(G294), .ZN(new_n567));
  OAI22_X1  g0367(.A1(new_n566), .A2(new_n474), .B1(new_n330), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n256), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n564), .A2(new_n469), .A3(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n570), .A2(new_n305), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n571), .B1(G200), .B2(new_n570), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n563), .A2(new_n572), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n555), .A2(KEYINPUT89), .A3(new_n558), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT89), .B1(new_n555), .B2(new_n558), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n537), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n570), .A2(new_n300), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(G179), .B2(new_n570), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n573), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n203), .A2(G97), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT80), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n584), .A2(KEYINPUT6), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT6), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n586), .A2(KEYINPUT80), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n583), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(KEYINPUT80), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n584), .A2(KEYINPUT6), .ZN(new_n590));
  NAND2_X1  g0390(.A1(G97), .A2(G107), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n204), .A2(new_n589), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n588), .A2(new_n592), .A3(G20), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n280), .A2(G77), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n203), .B1(new_n327), .B2(new_n332), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n279), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n294), .A2(G97), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n514), .B2(G97), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n472), .A2(new_n473), .A3(G244), .A4(new_n248), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT4), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n247), .A2(KEYINPUT4), .A3(G244), .A4(new_n248), .ZN(new_n604));
  NAND2_X1  g0404(.A1(G33), .A2(G283), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n247), .A2(G250), .A3(G1698), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n603), .A2(new_n604), .A3(new_n605), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n256), .ZN(new_n608));
  OAI211_X1 g0408(.A(G257), .B(new_n255), .C1(new_n462), .C2(new_n464), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n609), .A2(new_n469), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n600), .B1(G200), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(new_n305), .B2(new_n611), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n608), .A2(new_n610), .A3(KEYINPUT81), .A4(new_n372), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n600), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n608), .A2(new_n372), .A3(new_n610), .ZN(new_n616));
  AOI21_X1  g0416(.A(G169), .B1(new_n608), .B2(new_n610), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT81), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n613), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g0421(.A(new_n621), .B(KEYINPUT82), .ZN(new_n622));
  AND4_X1   g0422(.A1(new_n443), .A2(new_n531), .A3(new_n582), .A4(new_n622), .ZN(G372));
  NAND2_X1  g0423(.A1(new_n377), .A2(new_n378), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n439), .A2(new_n440), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(new_n404), .B2(new_n432), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n367), .A2(new_n379), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n624), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n319), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(KEYINPUT10), .B2(new_n312), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n302), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n563), .A2(KEYINPUT92), .A3(new_n578), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT92), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n634), .B1(new_n576), .B2(new_n579), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n492), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n516), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n513), .A2(new_n515), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n505), .A2(new_n357), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT91), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n525), .B2(new_n523), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n524), .A2(G179), .A3(new_n496), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n643), .B(KEYINPUT91), .C1(new_n300), .C2(new_n505), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n640), .B1(new_n645), .B2(new_n522), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n646), .A2(new_n613), .A3(new_n620), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n647), .A2(new_n573), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n600), .A2(new_n614), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n609), .A2(new_n469), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n650), .B1(new_n256), .B2(new_n607), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT81), .B1(new_n651), .B2(G169), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n649), .B1(new_n616), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n645), .A2(new_n522), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n653), .A2(new_n654), .A3(new_n655), .A4(new_n517), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n517), .A2(new_n526), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT26), .B1(new_n620), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n656), .A2(new_n654), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(KEYINPUT93), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n615), .A2(new_n619), .A3(new_n526), .A4(new_n517), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n661), .A2(KEYINPUT26), .B1(new_n522), .B2(new_n645), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT93), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(new_n663), .A3(new_n656), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n636), .A2(new_n648), .B1(new_n660), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n632), .B1(new_n442), .B2(new_n665), .ZN(G369));
  INV_X1    g0466(.A(G330), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n293), .A2(new_n207), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(G213), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(G343), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n492), .B(new_n530), .C1(new_n461), .C2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n485), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n676), .A2(G179), .A3(new_n528), .ZN(new_n677));
  INV_X1    g0477(.A(new_n491), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n490), .B1(new_n487), .B2(new_n485), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n680), .A2(new_n528), .A3(new_n673), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n667), .B1(new_n675), .B2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n563), .A2(new_n674), .ZN(new_n683));
  OAI22_X1  g0483(.A1(new_n581), .A2(new_n683), .B1(new_n580), .B2(new_n674), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n580), .A2(KEYINPUT92), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n576), .A2(new_n634), .A3(new_n579), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(new_n687), .A3(new_n674), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n680), .A2(new_n573), .A3(new_n580), .A4(new_n674), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n685), .A2(new_n691), .ZN(G399));
  INV_X1    g0492(.A(new_n210), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(new_n262), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n204), .A2(G87), .A3(G116), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G1), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n226), .B2(new_n695), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  OR3_X1    g0499(.A1(new_n665), .A2(KEYINPUT29), .A3(new_n673), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n531), .A2(new_n622), .A3(new_n582), .A4(new_n674), .ZN(new_n701));
  AND4_X1   g0501(.A1(new_n523), .A2(new_n651), .A3(new_n564), .A4(new_n569), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n676), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT30), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n676), .A2(new_n702), .A3(KEYINPUT30), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n570), .A2(new_n372), .A3(new_n611), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n505), .B(KEYINPUT94), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(new_n485), .A3(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n705), .A2(new_n706), .A3(new_n709), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n710), .A2(KEYINPUT31), .A3(new_n673), .ZN(new_n711));
  AOI21_X1  g0511(.A(KEYINPUT31), .B1(new_n710), .B2(new_n673), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n701), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n561), .A2(new_n562), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n578), .B1(new_n716), .B2(new_n537), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n647), .B(new_n573), .C1(new_n680), .C2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n655), .B1(new_n646), .B2(new_n653), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n654), .B1(new_n661), .B2(KEYINPUT26), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n673), .B1(new_n718), .B2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT29), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n700), .A2(new_n715), .A3(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n699), .B1(new_n726), .B2(G1), .ZN(G364));
  NOR2_X1   g0527(.A1(new_n292), .A2(G20), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n206), .B1(new_n728), .B2(G45), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n694), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n682), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n675), .A2(new_n667), .A3(new_n681), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G13), .A2(G33), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G20), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n675), .A2(new_n681), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n210), .A2(G355), .A3(new_n247), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n693), .A2(new_n247), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(G45), .B2(new_n226), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n245), .A2(new_n272), .ZN(new_n742));
  OAI221_X1 g0542(.A(new_n739), .B1(G116), .B2(new_n210), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n227), .B1(G20), .B2(new_n300), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n737), .A2(new_n744), .ZN(new_n745));
  AOI211_X1 g0545(.A(new_n694), .B(new_n730), .C1(new_n743), .C2(new_n745), .ZN(new_n746));
  XOR2_X1   g0546(.A(new_n746), .B(KEYINPUT95), .Z(new_n747));
  INV_X1    g0547(.A(new_n744), .ZN(new_n748));
  NOR4_X1   g0548(.A1(new_n207), .A2(new_n372), .A3(new_n305), .A4(G200), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n305), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n750), .A2(new_n335), .B1(new_n288), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n207), .A2(G190), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n756), .A2(new_n372), .A3(G200), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n757), .A2(KEYINPUT96), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(KEYINPUT96), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n754), .B1(new_n761), .B2(G77), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n762), .B(KEYINPUT97), .Z(new_n763));
  NOR2_X1   g0563(.A1(G179), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n755), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G159), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT32), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n372), .A2(G200), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT98), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n771), .A2(new_n207), .A3(new_n305), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G87), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n771), .A2(new_n756), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G107), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n207), .B1(new_n764), .B2(G190), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n474), .B1(new_n777), .B2(G97), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n773), .A2(new_n775), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n751), .A2(G190), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n768), .B(new_n779), .C1(G68), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n763), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n766), .A2(G329), .ZN(new_n783));
  INV_X1    g0583(.A(new_n757), .ZN(new_n784));
  INV_X1    g0584(.A(G311), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n247), .B(new_n786), .C1(G322), .C2(new_n749), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n776), .A2(new_n567), .ZN(new_n788));
  INV_X1    g0588(.A(new_n780), .ZN(new_n789));
  OR2_X1    g0589(.A1(KEYINPUT33), .A2(G317), .ZN(new_n790));
  NAND2_X1  g0590(.A1(KEYINPUT33), .A2(G317), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n788), .B(new_n792), .C1(G326), .C2(new_n752), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n774), .A2(G283), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n772), .A2(G303), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n787), .A2(new_n793), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n782), .A2(new_n796), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n738), .B(new_n747), .C1(new_n748), .C2(new_n797), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n734), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(G396));
  NOR2_X1   g0600(.A1(new_n405), .A2(new_n673), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(KEYINPUT101), .B1(new_n665), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n680), .B1(new_n686), .B2(new_n687), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n647), .A2(new_n573), .ZN(new_n805));
  AND3_X1   g0605(.A1(new_n662), .A2(new_n663), .A3(new_n656), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n663), .B1(new_n662), .B2(new_n656), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n804), .A2(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT101), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n808), .A2(new_n809), .A3(new_n801), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n803), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n401), .B1(new_n400), .B2(new_n674), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n404), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n404), .A2(new_n673), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(new_n808), .B2(new_n674), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n812), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n731), .B1(new_n821), .B2(new_n715), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n715), .B2(new_n821), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n748), .A2(new_n736), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n731), .B1(G77), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n247), .B1(new_n772), .B2(G107), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT99), .Z(new_n827));
  INV_X1    g0627(.A(G283), .ZN(new_n828));
  INV_X1    g0628(.A(G303), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n789), .A2(new_n828), .B1(new_n753), .B2(new_n829), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n750), .A2(new_n567), .B1(new_n765), .B2(new_n785), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n830), .B(new_n831), .C1(G97), .C2(new_n777), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n761), .A2(new_n448), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n774), .A2(G87), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n827), .A2(new_n832), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n749), .A2(G143), .B1(G137), .B2(new_n752), .ZN(new_n836));
  INV_X1    g0636(.A(G150), .ZN(new_n837));
  INV_X1    g0637(.A(G159), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n836), .B1(new_n837), .B2(new_n789), .C1(new_n760), .C2(new_n838), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT34), .Z(new_n840));
  NAND2_X1  g0640(.A1(new_n774), .A2(G68), .ZN(new_n841));
  INV_X1    g0641(.A(G132), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n247), .B1(new_n765), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G58), .B2(new_n777), .ZN(new_n844));
  INV_X1    g0644(.A(new_n772), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n841), .B(new_n844), .C1(new_n845), .C2(new_n288), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT100), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n835), .B1(new_n840), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n825), .B1(new_n848), .B2(new_n744), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n818), .B2(new_n736), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n823), .A2(new_n850), .ZN(G384));
  NOR3_X1   g0651(.A1(new_n227), .A2(new_n207), .A3(new_n446), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n588), .A2(new_n592), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT35), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n854), .B2(new_n853), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT36), .Z(new_n857));
  OAI21_X1  g0657(.A(G77), .B1(new_n335), .B2(new_n215), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n858), .A2(new_n226), .B1(G50), .B2(new_n215), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n859), .A2(G1), .A3(new_n292), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT102), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n625), .A2(new_n673), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT104), .ZN(new_n864));
  INV_X1    g0664(.A(new_n671), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n370), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT104), .B1(new_n349), .B2(new_n671), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT37), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n370), .A2(new_n375), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n868), .A2(new_n869), .A3(new_n870), .A4(new_n365), .ZN(new_n871));
  INV_X1    g0671(.A(new_n365), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n345), .A2(new_n369), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n374), .B2(new_n671), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT37), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n873), .A2(new_n671), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n380), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n876), .A2(KEYINPUT38), .A3(new_n878), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n881), .A2(KEYINPUT39), .A3(new_n882), .ZN(new_n883));
  AOI221_X4 g0683(.A(new_n880), .B1(new_n380), .B2(new_n877), .C1(new_n871), .C2(new_n875), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n866), .A2(new_n867), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n870), .A2(new_n365), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT37), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n871), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT105), .B1(new_n381), .B2(new_n868), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT105), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n380), .A2(new_n885), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n884), .B1(new_n892), .B2(new_n880), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n863), .B(new_n883), .C1(new_n893), .C2(KEYINPUT39), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n665), .A2(KEYINPUT101), .A3(new_n802), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n809), .B1(new_n808), .B2(new_n801), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n816), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n881), .A2(new_n882), .ZN(new_n898));
  INV_X1    g0698(.A(new_n432), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n440), .A2(new_n673), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n625), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT103), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n441), .A2(KEYINPUT103), .A3(new_n900), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n432), .A2(new_n439), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n906), .A2(new_n900), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n897), .A2(new_n898), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n624), .A2(new_n671), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n894), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n700), .A2(new_n724), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n631), .B1(new_n913), .B2(new_n443), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n912), .B(new_n914), .Z(new_n915));
  NAND3_X1  g0715(.A1(new_n909), .A2(new_n714), .A3(new_n818), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT40), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n892), .A2(new_n880), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n882), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n881), .A2(new_n882), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n917), .B1(new_n922), .B2(new_n916), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n443), .A2(new_n714), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n926), .A2(G330), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n915), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n206), .B2(new_n728), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n915), .A2(new_n928), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n862), .B1(new_n930), .B2(new_n931), .ZN(G367));
  NAND2_X1  g0732(.A1(new_n638), .A2(new_n673), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n646), .A2(new_n933), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n934), .A2(KEYINPUT106), .B1(new_n654), .B2(new_n933), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(KEYINPUT106), .B2(new_n934), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT43), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n936), .B(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n600), .A2(new_n673), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n613), .A2(new_n620), .A3(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n940), .A2(KEYINPUT107), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(KEYINPUT107), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(KEYINPUT108), .B1(new_n620), .B2(new_n674), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT108), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n653), .A2(new_n945), .A3(new_n673), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n680), .A2(new_n674), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n948), .A2(KEYINPUT42), .A3(new_n582), .A4(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT42), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n941), .A2(new_n942), .B1(new_n944), .B2(new_n946), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n952), .B1(new_n953), .B2(new_n689), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n620), .B1(new_n953), .B2(new_n580), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n674), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n938), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT109), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n951), .A2(new_n954), .B1(new_n956), .B2(new_n674), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n936), .A2(new_n937), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n958), .A2(new_n959), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n685), .A2(new_n953), .ZN(new_n964));
  OAI21_X1  g0764(.A(KEYINPUT109), .B1(new_n960), .B2(new_n938), .ZN(new_n965));
  AND3_X1   g0765(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n964), .B1(new_n963), .B2(new_n965), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n694), .B(KEYINPUT41), .Z(new_n969));
  INV_X1    g0769(.A(KEYINPUT110), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n948), .A2(new_n970), .A3(new_n688), .A4(new_n689), .ZN(new_n971));
  OAI21_X1  g0771(.A(KEYINPUT110), .B1(new_n953), .B2(new_n690), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT45), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n953), .A2(new_n690), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT44), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n976), .B(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n971), .A2(new_n972), .A3(KEYINPUT45), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n975), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n685), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n682), .A2(KEYINPUT111), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n689), .B1(new_n684), .B2(new_n950), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT111), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n986), .B(new_n667), .C1(new_n675), .C2(new_n681), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n984), .B1(new_n983), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n989), .A2(new_n725), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n975), .A2(new_n978), .A3(new_n685), .A4(new_n979), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n982), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n969), .B1(new_n992), .B2(new_n726), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n968), .B1(new_n993), .B2(new_n730), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT112), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n968), .B(KEYINPUT112), .C1(new_n993), .C2(new_n730), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n936), .A2(new_n737), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT46), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n1000), .A2(new_n446), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n761), .A2(G283), .B1(new_n772), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(G317), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n474), .B1(new_n765), .B2(new_n1003), .C1(new_n750), .C2(new_n829), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(G97), .B2(new_n774), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1000), .B1(new_n845), .B2(new_n447), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n753), .A2(new_n785), .B1(new_n776), .B2(new_n203), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(G294), .B2(new_n780), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1002), .A2(new_n1005), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n761), .A2(G50), .B1(new_n774), .B2(G77), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n776), .A2(new_n215), .ZN(new_n1011));
  INV_X1    g0811(.A(G143), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n753), .A2(new_n1012), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1011), .B(new_n1013), .C1(G159), .C2(new_n780), .ZN(new_n1014));
  INV_X1    g0814(.A(G137), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n247), .B1(new_n765), .B2(new_n1015), .C1(new_n750), .C2(new_n837), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G58), .B2(new_n772), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1010), .A2(new_n1014), .A3(new_n1017), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n1009), .A2(new_n1018), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1019), .A2(KEYINPUT47), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(KEYINPUT47), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1020), .A2(new_n744), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n740), .A2(new_n237), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1023), .B(new_n745), .C1(new_n210), .C2(new_n397), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n731), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT113), .Z(new_n1026));
  NAND3_X1  g0826(.A1(new_n999), .A2(new_n1022), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n998), .A2(new_n1027), .ZN(G387));
  INV_X1    g0828(.A(new_n989), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n737), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n684), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n696), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1032), .A2(new_n210), .A3(new_n247), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(G107), .B2(new_n210), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n234), .A2(G45), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n740), .ZN(new_n1036));
  AOI211_X1 g0836(.A(G45), .B(new_n1032), .C1(G68), .C2(G77), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n285), .A2(G50), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1038), .B(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1036), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1034), .B1(new_n1035), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n745), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n731), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n774), .A2(new_n448), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n247), .B1(new_n766), .B2(G326), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n845), .A2(new_n567), .B1(new_n828), .B2(new_n776), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n750), .A2(new_n1003), .B1(new_n785), .B2(new_n789), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(G322), .B2(new_n752), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n829), .B2(new_n760), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT48), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1047), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n1051), .B2(new_n1050), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT49), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1045), .B(new_n1046), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n777), .A2(new_n519), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n789), .B2(new_n285), .C1(new_n838), .C2(new_n753), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n772), .A2(G77), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n774), .A2(G97), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n474), .B1(new_n766), .B2(G150), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n757), .A2(G68), .B1(new_n749), .B2(G50), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n1055), .A2(new_n1056), .B1(new_n1058), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1044), .B1(new_n1064), .B2(new_n744), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n1029), .A2(new_n730), .B1(new_n1031), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n694), .B1(new_n989), .B2(new_n725), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT115), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n1067), .A2(new_n1068), .B1(new_n726), .B2(new_n1029), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1066), .B1(new_n1069), .B2(new_n1070), .ZN(G393));
  INV_X1    g0871(.A(KEYINPUT116), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n992), .A2(new_n694), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n990), .B1(new_n982), .B2(new_n991), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n982), .A2(new_n730), .A3(new_n991), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n242), .A2(new_n1036), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n745), .B1(new_n202), .B2(new_n210), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n731), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n750), .A2(new_n838), .B1(new_n837), .B2(new_n753), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT51), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n776), .A2(new_n250), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n247), .B1(new_n765), .B2(new_n1012), .C1(new_n789), .C2(new_n288), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n1081), .B2(new_n1080), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n834), .B1(new_n845), .B2(new_n215), .C1(new_n760), .C2(new_n285), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n749), .A2(G311), .B1(G317), .B2(new_n752), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT52), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n474), .B1(new_n784), .B2(new_n567), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G322), .B2(new_n766), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n777), .A2(new_n448), .B1(G303), .B2(new_n780), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n772), .A2(G283), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1091), .A2(new_n775), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n1086), .A2(new_n1087), .B1(new_n1089), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1079), .B1(new_n1095), .B2(new_n744), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n948), .B2(new_n1030), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1076), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1072), .B1(new_n1075), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1098), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1100), .B(KEYINPUT116), .C1(new_n1074), .C2(new_n1073), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1099), .A2(new_n1101), .ZN(G390));
  INV_X1    g0902(.A(new_n863), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n815), .B1(new_n803), .B2(new_n810), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n907), .B1(new_n903), .B2(new_n904), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1103), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n883), .B1(new_n893), .B2(KEYINPUT39), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n815), .B1(new_n722), .B2(new_n814), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1103), .B1(new_n1109), .B2(new_n1105), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n893), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n667), .B1(new_n701), .B2(new_n713), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1112), .A2(new_n818), .A3(new_n909), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT117), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1111), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1108), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1117), .B1(new_n1108), .B2(new_n1116), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1105), .B1(new_n715), .B2(new_n817), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1104), .B1(new_n1121), .B2(new_n1113), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1121), .A2(new_n1113), .A3(new_n1109), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n443), .A2(new_n1112), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n914), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1120), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1127), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1130), .A2(new_n694), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1107), .A2(new_n735), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n731), .B1(new_n322), .B2(new_n824), .ZN(new_n1135));
  XOR2_X1   g0935(.A(KEYINPUT54), .B(G143), .Z(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT118), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n760), .A2(new_n1137), .B1(new_n1015), .B2(new_n789), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1138), .B(KEYINPUT119), .Z(new_n1139));
  OR3_X1    g0939(.A1(new_n845), .A2(KEYINPUT53), .A3(new_n837), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n774), .A2(G50), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n474), .B1(new_n766), .B2(G125), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n842), .B2(new_n750), .ZN(new_n1143));
  INV_X1    g0943(.A(G128), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n753), .A2(new_n1144), .B1(new_n776), .B2(new_n838), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(KEYINPUT53), .B1(new_n845), .B2(new_n837), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1140), .A2(new_n1141), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n750), .A2(new_n446), .B1(new_n765), .B2(new_n567), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n789), .A2(new_n203), .B1(new_n753), .B2(new_n828), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n1149), .A2(new_n1083), .A3(new_n1150), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1151), .B(new_n841), .C1(new_n202), .C2(new_n760), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n773), .A2(new_n474), .ZN(new_n1153));
  XOR2_X1   g0953(.A(new_n1153), .B(KEYINPUT120), .Z(new_n1154));
  OAI22_X1  g0954(.A1(new_n1139), .A2(new_n1148), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1135), .B1(new_n1155), .B2(new_n744), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1134), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n1120), .B2(new_n729), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1133), .A2(new_n1159), .ZN(G378));
  OAI21_X1  g0960(.A(new_n731), .B1(G50), .B2(new_n824), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n474), .B(new_n266), .C1(new_n784), .C2(new_n397), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n750), .A2(new_n203), .B1(new_n765), .B2(new_n828), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n753), .A2(new_n446), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1011), .B(new_n1165), .C1(G97), .C2(new_n780), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n774), .A2(G58), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1164), .A2(new_n1059), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT58), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n288), .B1(G33), .B2(G41), .C1(new_n262), .C2(new_n247), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n784), .A2(new_n1015), .B1(new_n1144), .B2(new_n750), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G132), .B2(new_n780), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n777), .A2(G150), .B1(G125), .B2(new_n752), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1172), .B(new_n1173), .C1(new_n845), .C2(new_n1137), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(KEYINPUT59), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n774), .A2(G159), .ZN(new_n1176));
  AOI211_X1 g0976(.A(G33), .B(G41), .C1(new_n766), .C2(G124), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1174), .A2(KEYINPUT59), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1169), .B(new_n1170), .C1(new_n1178), .C2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT121), .ZN(new_n1181));
  OR2_X1    g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n748), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1161), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n299), .A2(new_n865), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n320), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1185), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n630), .B2(new_n303), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1186), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1184), .B1(new_n1194), .B2(new_n736), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n921), .A2(new_n923), .A3(G330), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n911), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1105), .B1(new_n811), .B2(new_n816), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1198), .B1(new_n1199), .B2(new_n898), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1194), .B1(new_n1200), .B2(new_n894), .ZN(new_n1201));
  AND4_X1   g1001(.A1(new_n894), .A2(new_n910), .A3(new_n911), .A4(new_n1194), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1197), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1194), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n912), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1200), .A2(new_n894), .A3(new_n1194), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1197), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1203), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1196), .B1(new_n1209), .B2(new_n730), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1132), .A2(new_n1128), .B1(new_n1203), .B2(new_n1208), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n694), .B1(new_n1211), .B2(KEYINPUT57), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1132), .A2(new_n1128), .ZN(new_n1213));
  AND3_X1   g1013(.A1(new_n1213), .A2(KEYINPUT57), .A3(new_n1209), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1210), .B1(new_n1212), .B2(new_n1214), .ZN(G375));
  NOR2_X1   g1015(.A1(new_n1131), .A2(new_n969), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1125), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n1127), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n731), .B1(G68), .B2(new_n824), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n474), .B1(new_n765), .B2(new_n829), .C1(new_n750), .C2(new_n828), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G77), .B2(new_n774), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1222), .B1(new_n202), .B2(new_n845), .C1(new_n203), .C2(new_n760), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1057), .B1(new_n789), .B2(new_n447), .C1(new_n567), .C2(new_n753), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n474), .B1(new_n757), .B2(G150), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(G128), .A2(new_n766), .B1(new_n749), .B2(G137), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n777), .A2(G50), .B1(G132), .B2(new_n752), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1167), .B1(new_n1137), .B2(new_n789), .C1(new_n845), .C2(new_n838), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n1223), .A2(new_n1224), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1220), .B1(new_n1230), .B2(new_n744), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n909), .B2(new_n736), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n729), .B(KEYINPUT122), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1232), .B1(new_n1217), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1219), .A2(new_n1235), .ZN(G381));
  OAI211_X1 g1036(.A(new_n799), .B(new_n1066), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1237));
  OR4_X1    g1037(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1237), .ZN(new_n1238));
  OR4_X1    g1038(.A1(G387), .A2(new_n1238), .A3(G378), .A4(G375), .ZN(G407));
  AOI21_X1  g1039(.A(new_n695), .B1(new_n1120), .B2(new_n1129), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1158), .B1(new_n1132), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n672), .A2(G213), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1241), .A2(new_n1243), .ZN(new_n1244));
  OAI211_X1 g1044(.A(G407), .B(G213), .C1(G375), .C2(new_n1244), .ZN(G409));
  INV_X1    g1045(.A(KEYINPUT61), .ZN(new_n1246));
  INV_X1    g1046(.A(G390), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(G387), .A2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n998), .A2(new_n1027), .A3(G390), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(G393), .A2(G396), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT125), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n1250), .A2(new_n1251), .A3(new_n1237), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1251), .B1(new_n1250), .B2(new_n1237), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1248), .A2(new_n1249), .A3(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1253), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1246), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  OAI211_X1 g1058(.A(G378), .B(new_n1210), .C1(new_n1212), .C2(new_n1214), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1213), .A2(new_n1209), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1260), .A2(new_n969), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1209), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1195), .B1(new_n1262), .B2(new_n1233), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1241), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1243), .B1(new_n1259), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT60), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1218), .B1(new_n1131), .B2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1217), .A2(KEYINPUT60), .A3(new_n1127), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1267), .A2(new_n694), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1235), .ZN(new_n1270));
  INV_X1    g1070(.A(G384), .ZN(new_n1271));
  OR2_X1    g1071(.A1(new_n1271), .A2(KEYINPUT124), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(KEYINPUT124), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1270), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1269), .A2(KEYINPUT124), .A3(new_n1271), .A4(new_n1235), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT63), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1258), .B1(new_n1265), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1259), .A2(new_n1264), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT123), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1259), .A2(new_n1264), .A3(KEYINPUT123), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1283), .A2(new_n1242), .A3(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1243), .A2(G2897), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1276), .A2(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1274), .A2(G2897), .A3(new_n1243), .A4(new_n1275), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1285), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1283), .A2(new_n1242), .A3(new_n1276), .A4(new_n1284), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1278), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1280), .A2(new_n1289), .A3(new_n1291), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1293), .B1(new_n1294), .B2(new_n1265), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT62), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1290), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1265), .A2(KEYINPUT62), .A3(new_n1276), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1295), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  OR2_X1    g1099(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1292), .B1(new_n1299), .B2(new_n1300), .ZN(G405));
  NAND2_X1  g1101(.A1(G375), .A2(new_n1241), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1259), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(new_n1303), .B(new_n1277), .ZN(new_n1304));
  XNOR2_X1  g1104(.A(new_n1304), .B(new_n1300), .ZN(G402));
endmodule


