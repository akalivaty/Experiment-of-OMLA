//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT75), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G204gat), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n204), .B1(KEYINPUT22), .B2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G211gat), .B(G218gat), .Z(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G162gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G155gat), .ZN(new_n212));
  INV_X1    g011(.A(G155gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G162gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT78), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n212), .A2(new_n214), .A3(KEYINPUT78), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT79), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(new_n211), .ZN(new_n221));
  NAND2_X1  g020(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n213), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT2), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT80), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(G141gat), .B(G148gat), .Z(new_n226));
  INV_X1    g025(.A(KEYINPUT80), .ZN(new_n227));
  AND2_X1   g026(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n227), .B(KEYINPUT2), .C1(new_n230), .C2(new_n213), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n219), .A2(new_n225), .A3(new_n226), .A4(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n226), .A2(new_n224), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(new_n215), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT29), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n210), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n232), .A2(KEYINPUT81), .A3(new_n235), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT81), .B1(new_n232), .B2(new_n235), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n209), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n208), .B(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n233), .B1(new_n245), .B2(KEYINPUT29), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n239), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  AND2_X1   g046(.A1(G228gat), .A2(G233gat), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n235), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n249), .ZN(new_n252));
  OAI22_X1  g051(.A1(new_n247), .A2(new_n249), .B1(new_n252), .B2(new_n239), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(G22gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(G78gat), .B(G106gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(KEYINPUT31), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n256), .B(G50gat), .Z(new_n257));
  INV_X1    g056(.A(KEYINPUT85), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n254), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n257), .B(KEYINPUT85), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n260), .B1(new_n254), .B2(new_n261), .ZN(new_n262));
  AND2_X1   g061(.A1(G227gat), .A2(G233gat), .ZN(new_n263));
  INV_X1    g062(.A(G113gat), .ZN(new_n264));
  INV_X1    g063(.A(G120gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT1), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n267), .B1(G113gat), .B2(G120gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n272), .A2(G127gat), .ZN(new_n273));
  INV_X1    g072(.A(G127gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n274), .A2(KEYINPUT69), .ZN(new_n275));
  OAI21_X1  g074(.A(G134gat), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(G127gat), .A2(G134gat), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n271), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(G134gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n274), .A2(KEYINPUT69), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n272), .A2(G127gat), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NOR3_X1   g082(.A1(new_n283), .A2(KEYINPUT70), .A3(new_n277), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n270), .B1(new_n279), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT70), .B1(new_n283), .B2(new_n277), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT69), .B(G127gat), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n271), .B(new_n278), .C1(new_n289), .C2(new_n280), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(KEYINPUT71), .A3(new_n270), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  XOR2_X1   g092(.A(KEYINPUT72), .B(G120gat), .Z(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT73), .B(G113gat), .ZN(new_n295));
  OAI22_X1  g094(.A1(new_n294), .A2(new_n264), .B1(new_n295), .B2(new_n265), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n274), .A2(new_n280), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n296), .B(new_n267), .C1(new_n277), .C2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT67), .ZN(new_n299));
  NAND2_X1  g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT65), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT65), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n302), .A2(G169gat), .A3(G176gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G169gat), .ZN(new_n305));
  INV_X1    g104(.A(G176gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT23), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT23), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(G169gat), .B2(G176gat), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n304), .A2(KEYINPUT25), .A3(new_n307), .A4(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n311), .B1(G183gat), .B2(G190gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(G183gat), .A2(G190gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT66), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT24), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n312), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n299), .B1(new_n310), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n314), .A2(new_n315), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT24), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(new_n320), .A3(new_n313), .ZN(new_n321));
  NOR2_X1   g120(.A1(G183gat), .A2(G190gat), .ZN(new_n322));
  AND2_X1   g121(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n322), .B1(new_n323), .B2(G190gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n307), .A2(new_n309), .A3(KEYINPUT25), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n325), .A2(KEYINPUT67), .A3(new_n326), .A4(new_n304), .ZN(new_n327));
  OR2_X1    g126(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n328), .A2(KEYINPUT23), .A3(new_n305), .A4(new_n329), .ZN(new_n330));
  AND2_X1   g129(.A1(G169gat), .A2(G176gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n305), .A2(new_n306), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n331), .B1(new_n332), .B2(new_n308), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n330), .B(new_n333), .C1(new_n312), .C2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT25), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n318), .A2(new_n327), .A3(new_n337), .ZN(new_n338));
  OR3_X1    g137(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(new_n340), .A3(new_n300), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(new_n314), .ZN(new_n342));
  NAND2_X1  g141(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n343));
  AOI21_X1  g142(.A(G190gat), .B1(new_n343), .B2(KEYINPUT27), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n344), .B1(KEYINPUT27), .B2(new_n343), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT28), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT27), .B(G183gat), .ZN(new_n348));
  INV_X1    g147(.A(G190gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(KEYINPUT28), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n342), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n338), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n293), .A2(new_n298), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT71), .B1(new_n291), .B2(new_n270), .ZN(new_n355));
  AOI211_X1 g154(.A(new_n286), .B(new_n269), .C1(new_n288), .C2(new_n290), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n298), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n325), .A2(new_n304), .A3(new_n326), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n358), .A2(new_n299), .B1(new_n335), .B2(new_n336), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n351), .B1(new_n359), .B2(new_n327), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n263), .B1(new_n354), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n354), .A2(new_n361), .A3(new_n263), .ZN(new_n364));
  XOR2_X1   g163(.A(G71gat), .B(G99gat), .Z(new_n365));
  XNOR2_X1  g164(.A(G15gat), .B(G43gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT33), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n364), .A2(KEYINPUT32), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT74), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT74), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n364), .A2(new_n371), .A3(KEYINPUT32), .A4(new_n368), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT34), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n364), .A2(KEYINPUT32), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT33), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n364), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n375), .A2(new_n377), .A3(new_n367), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n373), .A2(new_n374), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n374), .B1(new_n373), .B2(new_n378), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n363), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n373), .A2(new_n378), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT34), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n373), .A2(new_n374), .A3(new_n378), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n362), .A3(new_n384), .ZN(new_n385));
  AND3_X1   g184(.A1(new_n381), .A2(new_n385), .A3(KEYINPUT90), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT90), .B1(new_n381), .B2(new_n385), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n262), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G8gat), .B(G36gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(G64gat), .ZN(new_n390));
  INV_X1    g189(.A(G92gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G226gat), .ZN(new_n393));
  INV_X1    g192(.A(G233gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n353), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT29), .B1(new_n338), .B2(new_n352), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n396), .B(new_n210), .C1(new_n395), .C2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n395), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n360), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT76), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n401), .B1(new_n397), .B2(new_n395), .ZN(new_n402));
  OAI211_X1 g201(.A(KEYINPUT76), .B(new_n399), .C1(new_n360), .C2(KEYINPUT29), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n400), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n392), .B(new_n398), .C1(new_n404), .C2(new_n210), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(KEYINPUT77), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT30), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n398), .B1(new_n404), .B2(new_n210), .ZN(new_n409));
  INV_X1    g208(.A(new_n392), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n398), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n353), .A2(new_n238), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT76), .B1(new_n413), .B2(new_n399), .ZN(new_n414));
  NOR3_X1   g213(.A1(new_n397), .A2(new_n401), .A3(new_n395), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n396), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n412), .B1(new_n416), .B2(new_n245), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n417), .A2(KEYINPUT30), .A3(new_n392), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n408), .A2(new_n411), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  XOR2_X1   g219(.A(KEYINPUT84), .B(KEYINPUT0), .Z(new_n421));
  XNOR2_X1  g220(.A(G1gat), .B(G29gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G57gat), .B(G85gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  NAND4_X1  g224(.A1(new_n293), .A2(new_n235), .A3(new_n232), .A4(new_n298), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT4), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n236), .B1(new_n293), .B2(new_n298), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT81), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n250), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n431), .A2(KEYINPUT3), .A3(new_n240), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT82), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n429), .A2(KEYINPUT82), .A3(new_n432), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n428), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT5), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n426), .A2(new_n427), .ZN(new_n439));
  NAND2_X1  g238(.A1(G225gat), .A2(G233gat), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n437), .A2(new_n438), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  OR2_X1    g240(.A1(new_n426), .A2(new_n427), .ZN(new_n442));
  INV_X1    g241(.A(new_n440), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n426), .B1(new_n427), .B2(new_n443), .ZN(new_n444));
  AND4_X1   g243(.A1(KEYINPUT82), .A2(new_n432), .A3(new_n237), .A4(new_n357), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT82), .B1(new_n429), .B2(new_n432), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n442), .B(new_n444), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n243), .A2(new_n357), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n426), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n438), .B1(new_n449), .B2(new_n443), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n447), .A2(KEYINPUT83), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT83), .B1(new_n447), .B2(new_n450), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n425), .B(new_n441), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n447), .A2(new_n450), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT83), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n447), .A2(KEYINPUT83), .A3(new_n450), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n425), .B1(new_n460), .B2(new_n441), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n441), .B1(new_n451), .B2(new_n452), .ZN(new_n463));
  INV_X1    g262(.A(new_n425), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n463), .A2(KEYINPUT6), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n420), .B1(new_n462), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n202), .B1(new_n388), .B2(new_n467), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n379), .A2(new_n380), .A3(new_n363), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n362), .B1(new_n383), .B2(new_n384), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n262), .A2(new_n471), .A3(KEYINPUT35), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n463), .A2(new_n464), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n473), .A2(new_n454), .A3(new_n453), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n419), .B1(new_n474), .B2(new_n465), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n402), .A2(new_n403), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n245), .B1(new_n477), .B2(new_n396), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n396), .B(new_n245), .C1(new_n395), .C2(new_n397), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT37), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT88), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n479), .A2(KEYINPUT37), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT88), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n482), .B(new_n483), .C1(new_n245), .C2(new_n404), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT37), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n486), .B(new_n398), .C1(new_n404), .C2(new_n210), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n392), .A2(KEYINPUT38), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n406), .ZN(new_n491));
  INV_X1    g290(.A(new_n487), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n392), .B1(new_n409), .B2(KEYINPUT37), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n492), .B1(new_n493), .B2(KEYINPUT89), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n410), .B1(new_n417), .B2(new_n486), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT89), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n491), .B1(KEYINPUT38), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n474), .A2(new_n499), .A3(new_n465), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n437), .A2(new_n439), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n443), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT39), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n448), .A2(new_n426), .A3(new_n440), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT86), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n448), .A2(KEYINPUT86), .A3(new_n426), .A4(new_n440), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT87), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT87), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n506), .A2(new_n510), .A3(new_n507), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n502), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n440), .B1(new_n437), .B2(new_n439), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n464), .B1(new_n513), .B2(new_n503), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT40), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n512), .A2(KEYINPUT40), .A3(new_n514), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n517), .A2(new_n419), .A3(new_n473), .A4(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n500), .A2(new_n262), .A3(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n381), .A2(new_n385), .A3(KEYINPUT36), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT36), .B1(new_n381), .B2(new_n385), .ZN(new_n524));
  OAI22_X1  g323(.A1(new_n475), .A2(new_n262), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n468), .B(new_n476), .C1(new_n521), .C2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(G64gat), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n527), .A2(G57gat), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n527), .A2(G57gat), .ZN(new_n529));
  INV_X1    g328(.A(G71gat), .ZN(new_n530));
  INV_X1    g329(.A(G78gat), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI22_X1  g331(.A1(new_n528), .A2(new_n529), .B1(new_n532), .B2(KEYINPUT9), .ZN(new_n533));
  XOR2_X1   g332(.A(G71gat), .B(G78gat), .Z(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n533), .B(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n536), .A2(KEYINPUT21), .ZN(new_n537));
  XNOR2_X1  g336(.A(G127gat), .B(G155gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(new_n205), .ZN(new_n540));
  XOR2_X1   g339(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n541));
  NAND2_X1  g340(.A1(G231gat), .A2(G233gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n540), .B(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(G8gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(G15gat), .B(G22gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT16), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n546), .B1(new_n547), .B2(G1gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT93), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n545), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n548), .B1(G1gat), .B2(new_n546), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n552), .B1(KEYINPUT21), .B2(new_n536), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  OR2_X1    g353(.A1(new_n544), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n544), .A2(new_n554), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT95), .B(G183gat), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g361(.A1(G232gat), .A2(G233gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n563), .A2(KEYINPUT41), .ZN(new_n564));
  XNOR2_X1  g363(.A(G134gat), .B(G162gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n566), .B(KEYINPUT97), .Z(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  OR3_X1    g367(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n569), .A2(KEYINPUT91), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n571));
  NOR3_X1   g370(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT91), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G43gat), .B(G50gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT15), .ZN(new_n577));
  NAND2_X1  g376(.A1(G29gat), .A2(G36gat), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(G43gat), .B(G50gat), .Z(new_n580));
  INV_X1    g379(.A(KEYINPUT15), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n575), .A2(new_n579), .A3(KEYINPUT92), .A4(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT92), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n582), .A2(new_n578), .A3(new_n577), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n570), .A2(new_n574), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n569), .A2(new_n571), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n577), .B1(new_n589), .B2(new_n578), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G85gat), .A2(G92gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT7), .ZN(new_n594));
  NAND2_X1  g393(.A1(G99gat), .A2(G106gat), .ZN(new_n595));
  INV_X1    g394(.A(G85gat), .ZN(new_n596));
  AOI22_X1  g395(.A1(KEYINPUT8), .A2(new_n595), .B1(new_n596), .B2(new_n391), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G99gat), .B(G106gat), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT96), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n600), .B(KEYINPUT96), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n598), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  AOI22_X1  g405(.A1(new_n592), .A2(new_n606), .B1(KEYINPUT41), .B2(new_n563), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n590), .B1(new_n583), .B2(new_n587), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n603), .B(new_n605), .C1(new_n608), .C2(KEYINPUT17), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n608), .A2(KEYINPUT17), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G190gat), .B(G218gat), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n568), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n566), .A2(KEYINPUT97), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n613), .A2(new_n614), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G230gat), .A2(G233gat), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n599), .A2(new_n602), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n604), .A2(new_n598), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n536), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n533), .B(new_n534), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n624), .A2(new_n603), .A3(new_n605), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT10), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n623), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT98), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT98), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n623), .A2(new_n625), .A3(new_n629), .A4(new_n626), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT99), .B1(new_n623), .B2(new_n626), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT99), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n606), .A2(new_n633), .A3(KEYINPUT10), .A4(new_n536), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n620), .B1(new_n631), .B2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G176gat), .B(G204gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(KEYINPUT101), .B(G148gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT100), .B(G120gat), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n639), .B(new_n640), .Z(new_n641));
  AND2_X1   g440(.A1(new_n623), .A2(new_n625), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n636), .B(new_n641), .C1(new_n620), .C2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n641), .ZN(new_n644));
  AOI22_X1  g443(.A1(new_n628), .A2(new_n630), .B1(new_n632), .B2(new_n634), .ZN(new_n645));
  INV_X1    g444(.A(new_n620), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n642), .A2(new_n620), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n644), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n643), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n562), .A2(new_n619), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n592), .A2(new_n552), .ZN(new_n653));
  NAND2_X1  g452(.A1(G229gat), .A2(G233gat), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n550), .B(new_n551), .Z(new_n655));
  OAI21_X1  g454(.A(new_n655), .B1(new_n608), .B2(KEYINPUT17), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n653), .B(new_n654), .C1(new_n610), .C2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT18), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G113gat), .B(G141gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT11), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(new_n305), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G197gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT12), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n659), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n655), .A2(new_n608), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n653), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n654), .B(KEYINPUT13), .Z(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n669), .B1(new_n657), .B2(new_n658), .ZN(new_n670));
  OR3_X1    g469(.A1(new_n665), .A2(KEYINPUT94), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT94), .B1(new_n665), .B2(new_n670), .ZN(new_n672));
  INV_X1    g471(.A(new_n659), .ZN(new_n673));
  OR2_X1    g472(.A1(new_n673), .A2(new_n670), .ZN(new_n674));
  INV_X1    g473(.A(new_n664), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n671), .A2(new_n672), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n652), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n526), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n474), .A2(new_n465), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g481(.A1(new_n547), .A2(new_n545), .ZN(new_n683));
  NAND2_X1  g482(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n678), .A2(new_n419), .A3(new_n683), .A4(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT42), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n678), .ZN(new_n688));
  OAI21_X1  g487(.A(G8gat), .B1(new_n688), .B2(new_n420), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n685), .A2(new_n686), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n687), .A2(new_n689), .A3(new_n690), .ZN(G1325gat));
  INV_X1    g490(.A(new_n524), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT102), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n692), .A2(new_n693), .A3(new_n522), .ZN(new_n694));
  OAI21_X1  g493(.A(KEYINPUT102), .B1(new_n523), .B2(new_n524), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(G15gat), .B1(new_n688), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT90), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n699), .B1(new_n469), .B2(new_n470), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n381), .A2(new_n385), .A3(KEYINPUT90), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n703), .A2(G15gat), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n698), .B1(new_n688), .B2(new_n704), .ZN(G1326gat));
  INV_X1    g504(.A(new_n262), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n678), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(KEYINPUT43), .B(G22gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1327gat));
  INV_X1    g508(.A(new_n562), .ZN(new_n710));
  INV_X1    g509(.A(new_n676), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(new_n711), .A3(new_n651), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n619), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n526), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(G29gat), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n714), .A2(new_n715), .A3(new_n680), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT45), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n618), .A2(KEYINPUT44), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n526), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n712), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n702), .A2(new_n475), .A3(new_n262), .ZN(new_n721));
  AOI22_X1  g520(.A1(new_n721), .A2(new_n202), .B1(new_n475), .B2(new_n472), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n467), .A2(new_n706), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n723), .A2(new_n520), .A3(new_n694), .A4(new_n695), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n619), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n719), .B(new_n720), .C1(new_n725), .C2(KEYINPUT44), .ZN(new_n726));
  OAI21_X1  g525(.A(G29gat), .B1(new_n726), .B2(new_n679), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n717), .A2(new_n727), .ZN(G1328gat));
  INV_X1    g527(.A(G36gat), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n729), .A3(new_n419), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n730), .B(KEYINPUT46), .Z(new_n731));
  OAI21_X1  g530(.A(G36gat), .B1(new_n726), .B2(new_n420), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(G1329gat));
  OAI21_X1  g532(.A(G43gat), .B1(new_n726), .B2(new_n697), .ZN(new_n734));
  INV_X1    g533(.A(G43gat), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n714), .A2(new_n735), .A3(new_n702), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n737), .B(KEYINPUT47), .Z(G1330gat));
  NOR2_X1   g537(.A1(new_n262), .A2(G50gat), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n526), .A2(new_n713), .A3(new_n739), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n740), .A2(KEYINPUT103), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT48), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n740), .B2(KEYINPUT103), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(G50gat), .B1(new_n726), .B2(new_n262), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n742), .B1(new_n745), .B2(new_n740), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT104), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT104), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n745), .A2(new_n740), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n750), .B(new_n746), .C1(new_n751), .C2(new_n742), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n749), .A2(new_n752), .ZN(G1331gat));
  NAND2_X1  g552(.A1(new_n722), .A2(new_n724), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n562), .A2(new_n676), .A3(new_n619), .A4(new_n650), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n679), .ZN(new_n758));
  XOR2_X1   g557(.A(new_n758), .B(G57gat), .Z(G1332gat));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n757), .B(KEYINPUT105), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n419), .B(KEYINPUT106), .Z(new_n762));
  INV_X1    g561(.A(KEYINPUT49), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n763), .B2(new_n527), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT107), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n760), .B1(new_n761), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n761), .A2(new_n760), .A3(new_n765), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n767), .A2(new_n763), .A3(new_n527), .A4(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n768), .ZN(new_n770));
  OAI22_X1  g569(.A1(new_n770), .A2(new_n766), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(G1333gat));
  AOI21_X1  g571(.A(new_n530), .B1(new_n761), .B2(new_n696), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n754), .A2(new_n530), .A3(new_n702), .A4(new_n756), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  OR3_X1    g575(.A1(new_n773), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n774), .B1(new_n773), .B2(new_n776), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(G1334gat));
  NAND2_X1  g578(.A1(new_n761), .A2(new_n706), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g580(.A1(new_n562), .A2(new_n711), .A3(new_n651), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n719), .B(new_n782), .C1(new_n725), .C2(KEYINPUT44), .ZN(new_n783));
  OAI21_X1  g582(.A(G85gat), .B1(new_n783), .B2(new_n679), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n562), .A2(new_n711), .ZN(new_n785));
  AND4_X1   g584(.A1(KEYINPUT51), .A2(new_n754), .A3(new_n618), .A4(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT51), .B1(new_n725), .B2(new_n785), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n650), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n680), .A2(new_n596), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n784), .B1(new_n788), .B2(new_n789), .ZN(G1336gat));
  OAI21_X1  g589(.A(G92gat), .B1(new_n783), .B2(new_n420), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT109), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n762), .A2(new_n391), .A3(new_n650), .ZN(new_n794));
  XOR2_X1   g593(.A(new_n794), .B(KEYINPUT110), .Z(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(new_n786), .B2(new_n787), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI211_X1 g597(.A(KEYINPUT109), .B(G92gat), .C1(new_n783), .C2(new_n420), .ZN(new_n799));
  OAI211_X1 g598(.A(KEYINPUT111), .B(new_n795), .C1(new_n786), .C2(new_n787), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n793), .A2(new_n798), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT52), .ZN(new_n802));
  INV_X1    g601(.A(new_n762), .ZN(new_n803));
  OAI21_X1  g602(.A(G92gat), .B1(new_n783), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n804), .A2(new_n796), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n802), .A2(new_n806), .ZN(G1337gat));
  OAI21_X1  g606(.A(G99gat), .B1(new_n783), .B2(new_n697), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n703), .A2(G99gat), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n808), .B1(new_n788), .B2(new_n809), .ZN(G1338gat));
  OAI21_X1  g609(.A(G106gat), .B1(new_n783), .B2(new_n262), .ZN(new_n811));
  NAND2_X1  g610(.A1(KEYINPUT112), .A2(KEYINPUT53), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n262), .A2(G106gat), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n811), .B(new_n812), .C1(new_n788), .C2(new_n813), .ZN(new_n814));
  OR2_X1    g613(.A1(KEYINPUT112), .A2(KEYINPUT53), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n814), .B(new_n815), .ZN(G1339gat));
  NOR2_X1   g615(.A1(new_n652), .A2(new_n711), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n610), .A2(new_n656), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n654), .B1(new_n818), .B2(new_n653), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n667), .A2(new_n668), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n663), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n672), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n665), .A2(new_n670), .A3(KEYINPUT94), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n650), .B(new_n821), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n641), .B1(new_n647), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n645), .A2(new_n646), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n636), .A2(KEYINPUT54), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n828), .A3(KEYINPUT55), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(new_n643), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n826), .A2(new_n828), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n824), .B1(new_n834), .B2(new_n676), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n619), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n830), .A2(new_n618), .A3(new_n833), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n562), .B1(new_n836), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n817), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n842), .A2(new_n679), .ZN(new_n843));
  INV_X1    g642(.A(new_n388), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(new_n844), .A3(new_n803), .ZN(new_n845));
  OAI21_X1  g644(.A(G113gat), .B1(new_n845), .B2(new_n676), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n262), .A2(new_n471), .ZN(new_n847));
  NOR4_X1   g646(.A1(new_n842), .A2(new_n679), .A3(new_n847), .A4(new_n762), .ZN(new_n848));
  INV_X1    g647(.A(new_n295), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n849), .A3(new_n711), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n846), .A2(new_n850), .ZN(G1340gat));
  OAI21_X1  g650(.A(G120gat), .B1(new_n845), .B2(new_n651), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n651), .A2(new_n294), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(KEYINPUT113), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n848), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n852), .A2(new_n855), .ZN(G1341gat));
  NOR3_X1   g655(.A1(new_n845), .A2(new_n289), .A3(new_n710), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT114), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n858), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n848), .A2(KEYINPUT115), .A3(new_n562), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT115), .B1(new_n848), .B2(new_n562), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n862), .A2(new_n273), .A3(new_n275), .ZN(new_n863));
  AOI22_X1  g662(.A1(new_n859), .A2(new_n860), .B1(new_n861), .B2(new_n863), .ZN(G1342gat));
  NOR3_X1   g663(.A1(new_n419), .A2(new_n619), .A3(G134gat), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n843), .A2(new_n471), .A3(new_n262), .A4(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n867));
  OR3_X1    g666(.A1(new_n866), .A2(new_n867), .A3(KEYINPUT56), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n867), .B1(new_n866), .B2(KEYINPUT56), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n843), .A2(new_n844), .A3(new_n618), .A4(new_n803), .ZN(new_n871));
  AOI22_X1  g670(.A1(G134gat), .A2(new_n871), .B1(new_n866), .B2(KEYINPUT56), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT117), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n870), .A2(new_n875), .A3(new_n872), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(G1343gat));
  NOR4_X1   g676(.A1(new_n842), .A2(new_n679), .A3(new_n262), .A4(new_n696), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n676), .A2(G141gat), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n878), .A2(new_n803), .A3(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n880), .B(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(G141gat), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884));
  INV_X1    g683(.A(new_n817), .ZN(new_n885));
  XNOR2_X1  g684(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n831), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n643), .A3(new_n829), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n824), .B1(new_n888), .B2(new_n676), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n618), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n824), .B(KEYINPUT119), .C1(new_n888), .C2(new_n676), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n839), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n885), .B1(new_n562), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n884), .B1(new_n894), .B2(new_n706), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n884), .B(new_n706), .C1(new_n817), .C2(new_n841), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n696), .A2(new_n762), .A3(new_n679), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n883), .B1(new_n899), .B2(new_n711), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT58), .B1(new_n882), .B2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT58), .B1(new_n880), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n903), .B1(new_n902), .B2(new_n880), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n901), .B1(new_n900), .B2(new_n904), .ZN(G1344gat));
  INV_X1    g704(.A(new_n878), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n906), .A2(new_n762), .ZN(new_n907));
  INV_X1    g706(.A(G148gat), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n907), .A2(new_n908), .A3(new_n650), .ZN(new_n909));
  XNOR2_X1  g708(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n710), .B1(new_n893), .B2(KEYINPUT123), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT123), .ZN(new_n912));
  AOI211_X1 g711(.A(new_n912), .B(new_n839), .C1(new_n891), .C2(new_n892), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n885), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n262), .A2(KEYINPUT57), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT57), .B1(new_n842), .B2(new_n262), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n916), .A2(new_n650), .A3(new_n897), .A4(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n910), .B1(new_n918), .B2(G148gat), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n908), .A2(KEYINPUT59), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n920), .B1(new_n899), .B2(new_n650), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n909), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n909), .B(KEYINPUT124), .C1(new_n919), .C2(new_n921), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1345gat));
  AOI21_X1  g725(.A(G155gat), .B1(new_n907), .B2(new_n562), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n562), .A2(G155gat), .ZN(new_n928));
  XOR2_X1   g727(.A(new_n928), .B(KEYINPUT125), .Z(new_n929));
  AOI21_X1  g728(.A(new_n927), .B1(new_n899), .B2(new_n929), .ZN(G1346gat));
  NOR3_X1   g729(.A1(new_n895), .A2(new_n898), .A3(new_n619), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n420), .A2(new_n230), .A3(new_n618), .ZN(new_n932));
  OAI22_X1  g731(.A1(new_n931), .A2(new_n230), .B1(new_n906), .B2(new_n932), .ZN(new_n933));
  XOR2_X1   g732(.A(new_n933), .B(KEYINPUT126), .Z(G1347gat));
  INV_X1    g733(.A(new_n842), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n679), .A2(new_n419), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT127), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n935), .A2(new_n844), .A3(new_n937), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n938), .A2(new_n305), .A3(new_n676), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n842), .A2(new_n680), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n803), .A2(new_n847), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(new_n711), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n939), .B1(new_n944), .B2(new_n305), .ZN(G1348gat));
  AOI21_X1  g744(.A(G176gat), .B1(new_n943), .B2(new_n650), .ZN(new_n946));
  INV_X1    g745(.A(new_n938), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n651), .B1(new_n328), .B2(new_n329), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(G1349gat));
  OAI21_X1  g748(.A(G183gat), .B1(new_n938), .B2(new_n710), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n562), .A2(new_n348), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n950), .B1(new_n942), .B2(new_n951), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g752(.A(G190gat), .B1(new_n938), .B2(new_n619), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT61), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n943), .A2(new_n349), .A3(new_n618), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1351gat));
  AND4_X1   g756(.A1(new_n706), .A2(new_n940), .A3(new_n697), .A4(new_n762), .ZN(new_n958));
  AOI21_X1  g757(.A(G197gat), .B1(new_n958), .B2(new_n711), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n937), .A2(new_n697), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n916), .A2(new_n917), .A3(new_n961), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n711), .A2(G197gat), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(G1352gat));
  NOR2_X1   g763(.A1(new_n651), .A2(G204gat), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n958), .A2(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n967));
  OR2_X1    g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n916), .A2(new_n650), .A3(new_n917), .A4(new_n961), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(G204gat), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n966), .A2(new_n967), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(G1353gat));
  NAND3_X1  g771(.A1(new_n958), .A2(new_n205), .A3(new_n562), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n962), .A2(new_n562), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n974), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT63), .B1(new_n974), .B2(G211gat), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(G1354gat));
  AOI21_X1  g776(.A(G218gat), .B1(new_n958), .B2(new_n618), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n619), .A2(new_n206), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n978), .B1(new_n962), .B2(new_n979), .ZN(G1355gat));
endmodule


