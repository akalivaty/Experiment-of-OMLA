//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 0 1 1 0 0 0 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT77), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G221), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT78), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G469), .ZN(new_n194));
  NOR2_X1   g008(.A1(KEYINPUT84), .A2(KEYINPUT12), .ZN(new_n195));
  INV_X1    g009(.A(G101), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT79), .ZN(new_n197));
  INV_X1    g011(.A(G104), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT79), .A2(G104), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(G107), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n202));
  INV_X1    g016(.A(G107), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(G104), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(G107), .B1(new_n199), .B2(new_n200), .ZN(new_n207));
  NOR3_X1   g021(.A1(new_n207), .A2(KEYINPUT80), .A3(new_n202), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT80), .ZN(new_n209));
  INV_X1    g023(.A(new_n200), .ZN(new_n210));
  NOR2_X1   g024(.A1(KEYINPUT79), .A2(G104), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n203), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n209), .B1(new_n212), .B2(KEYINPUT3), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n196), .B(new_n206), .C1(new_n208), .C2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G143), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT65), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G143), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n218), .A3(G146), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G143), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n219), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n217), .A2(G143), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n215), .A2(KEYINPUT65), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n220), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n222), .B1(new_n227), .B2(KEYINPUT1), .ZN(new_n228));
  INV_X1    g042(.A(new_n221), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT65), .B(G143), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n229), .B1(new_n230), .B2(G146), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n224), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n198), .A2(G107), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n196), .B1(new_n212), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n214), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n220), .A2(G143), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n216), .A2(new_n218), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n237), .B1(new_n238), .B2(new_n220), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n222), .B1(new_n221), .B2(KEYINPUT1), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n224), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n241), .B1(new_n214), .B2(new_n235), .ZN(new_n242));
  OAI211_X1 g056(.A(KEYINPUT83), .B(new_n195), .C1(new_n236), .C2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n214), .A2(new_n232), .A3(new_n235), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT80), .B1(new_n207), .B2(new_n202), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n212), .A2(new_n209), .A3(KEYINPUT3), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n205), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n234), .B1(new_n247), .B2(new_n196), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n244), .B(KEYINPUT84), .C1(new_n248), .C2(new_n241), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n243), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT11), .ZN(new_n251));
  INV_X1    g065(.A(G134), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n251), .B1(new_n252), .B2(G137), .ZN(new_n253));
  INV_X1    g067(.A(G137), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(KEYINPUT11), .A3(G134), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n252), .A2(G137), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT67), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n253), .A2(new_n255), .A3(KEYINPUT67), .A4(new_n256), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT11), .B1(new_n254), .B2(G134), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n254), .A2(G134), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G131), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n264), .A2(KEYINPUT66), .A3(new_n265), .A4(new_n255), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n253), .A2(new_n255), .A3(new_n265), .A4(new_n256), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT66), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n261), .A2(G131), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  OAI211_X1 g085(.A(KEYINPUT83), .B(new_n271), .C1(new_n236), .C2(new_n242), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n250), .A2(new_n271), .B1(KEYINPUT12), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT81), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT4), .B1(new_n247), .B2(new_n196), .ZN(new_n275));
  AOI211_X1 g089(.A(G101), .B(new_n205), .C1(new_n245), .C2(new_n246), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n206), .B1(new_n208), .B2(new_n213), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT4), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n278), .A2(new_n279), .A3(G101), .ZN(new_n280));
  INV_X1    g094(.A(new_n237), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n227), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(KEYINPUT0), .A2(G128), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(KEYINPUT64), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT64), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n285), .B1(KEYINPUT0), .B2(G128), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n284), .B1(new_n283), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n283), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n282), .A2(new_n287), .B1(new_n231), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n280), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n274), .B1(new_n277), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n278), .A2(G101), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(KEYINPUT4), .A3(new_n214), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n293), .A2(KEYINPUT81), .A3(new_n289), .A4(new_n280), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT10), .B1(new_n248), .B2(new_n232), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n214), .A2(KEYINPUT82), .A3(new_n235), .ZN(new_n297));
  AOI21_X1  g111(.A(KEYINPUT82), .B1(new_n214), .B2(new_n235), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n241), .A2(KEYINPUT10), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n296), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n295), .A2(new_n301), .A3(new_n270), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n273), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G953), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT71), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT71), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G953), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G227), .ZN(new_n309));
  XNOR2_X1  g123(.A(G110), .B(G140), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n309), .B(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n303), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n295), .A2(new_n301), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n271), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(new_n311), .A3(new_n302), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n194), .B1(new_n317), .B2(new_n189), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n295), .A2(new_n270), .A3(new_n301), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n270), .B1(new_n295), .B2(new_n301), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n312), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n273), .A2(new_n302), .A3(new_n311), .ZN(new_n322));
  AOI211_X1 g136(.A(G469), .B(G902), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n193), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(G214), .B1(G237), .B2(G902), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT82), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n326), .B1(new_n276), .B2(new_n234), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n214), .A2(KEYINPUT82), .A3(new_n235), .ZN(new_n328));
  AND3_X1   g142(.A1(KEYINPUT69), .A2(KEYINPUT2), .A3(G113), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT69), .B1(KEYINPUT2), .B2(G113), .ZN(new_n330));
  OAI22_X1  g144(.A1(new_n329), .A2(new_n330), .B1(KEYINPUT2), .B2(G113), .ZN(new_n331));
  XNOR2_X1  g145(.A(G116), .B(G119), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(KEYINPUT5), .ZN(new_n335));
  INV_X1    g149(.A(G116), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n336), .A2(KEYINPUT5), .A3(G119), .ZN(new_n337));
  INV_X1    g151(.A(G113), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n334), .B1(new_n335), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n327), .A2(new_n328), .A3(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n331), .B(new_n332), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n343), .B(new_n280), .C1(new_n275), .C2(new_n276), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT6), .ZN(new_n346));
  XNOR2_X1  g160(.A(G110), .B(G122), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n345), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT86), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n347), .B1(new_n341), .B2(new_n344), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT86), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n352), .A3(new_n346), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n341), .A2(new_n344), .A3(new_n347), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT85), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n341), .A2(KEYINPUT85), .A3(new_n344), .A4(new_n347), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n351), .A2(new_n346), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n289), .A2(G125), .ZN(new_n362));
  INV_X1    g176(.A(G125), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n241), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G224), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(G953), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n365), .B1(new_n367), .B2(G953), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n354), .A2(new_n361), .A3(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(G210), .B1(G237), .B2(G902), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT7), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n366), .B1(new_n374), .B2(new_n368), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n375), .B1(new_n374), .B2(new_n370), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n347), .B(KEYINPUT8), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n248), .B(new_n340), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(G902), .B1(new_n379), .B2(new_n359), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n372), .A2(new_n373), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n373), .B1(new_n372), .B2(new_n380), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n325), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n324), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT92), .ZN(new_n385));
  NOR2_X1   g199(.A1(G475), .A2(G902), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT90), .ZN(new_n388));
  INV_X1    g202(.A(G237), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n305), .A2(new_n307), .A3(G214), .A4(new_n389), .ZN(new_n390));
  OR2_X1    g204(.A1(new_n390), .A2(new_n215), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n390), .A2(KEYINPUT87), .A3(new_n230), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT87), .B1(new_n390), .B2(new_n230), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n388), .B1(new_n394), .B2(G131), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(G131), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n390), .A2(new_n230), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT87), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n390), .A2(KEYINPUT87), .A3(new_n230), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n401), .A2(KEYINPUT90), .A3(new_n265), .A4(new_n391), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n395), .A2(new_n396), .A3(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(G125), .B(G140), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT16), .ZN(new_n405));
  OR3_X1    g219(.A1(new_n363), .A2(KEYINPUT16), .A3(G140), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(G146), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n404), .B(KEYINPUT19), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n408), .B1(new_n220), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n403), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n404), .B(G146), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n265), .B1(new_n401), .B2(new_n391), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n412), .B1(new_n413), .B2(KEYINPUT18), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT89), .ZN(new_n415));
  NAND2_X1  g229(.A1(KEYINPUT18), .A2(G131), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n391), .B(new_n416), .C1(new_n392), .C2(new_n393), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT88), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n401), .A2(KEYINPUT88), .A3(new_n391), .A4(new_n416), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n414), .A2(new_n415), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n415), .B1(new_n414), .B2(new_n421), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n411), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(G113), .B(G122), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT91), .B(G104), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n425), .B(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n427), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT17), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n395), .A2(new_n430), .A3(new_n402), .A4(new_n396), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n405), .A2(new_n406), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n220), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n407), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n434), .B1(new_n413), .B2(KEYINPUT17), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n429), .B(new_n436), .C1(new_n422), .C2(new_n423), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n387), .B1(new_n428), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT20), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n385), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n437), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n419), .A2(new_n420), .ZN(new_n442));
  INV_X1    g256(.A(new_n412), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT18), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n443), .B1(new_n396), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(KEYINPUT89), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n414), .A2(new_n415), .A3(new_n421), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n429), .B1(new_n448), .B2(new_n411), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n386), .B1(new_n441), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(KEYINPUT92), .A3(KEYINPUT20), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n446), .A2(new_n447), .B1(new_n403), .B2(new_n410), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n437), .B1(new_n452), .B2(new_n429), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(new_n439), .A3(new_n386), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n440), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G952), .ZN(new_n456));
  AOI211_X1 g270(.A(G953), .B(new_n456), .C1(G234), .C2(G237), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  AOI211_X1 g272(.A(new_n189), .B(new_n308), .C1(G234), .C2(G237), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT21), .B(G898), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n458), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n429), .B1(new_n448), .B2(new_n436), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n189), .B1(new_n441), .B2(new_n464), .ZN(new_n465));
  XOR2_X1   g279(.A(KEYINPUT93), .B(G475), .Z(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(G116), .B(G122), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(new_n203), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n215), .A2(G128), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n470), .B1(new_n230), .B2(G128), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n252), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n471), .A2(KEYINPUT13), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n230), .A2(G128), .ZN(new_n474));
  OAI21_X1  g288(.A(G134), .B1(new_n474), .B2(KEYINPUT13), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n469), .B(new_n472), .C1(new_n473), .C2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n336), .A2(G122), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n336), .A2(G122), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n477), .B1(new_n478), .B2(KEYINPUT14), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n479), .B1(KEYINPUT14), .B2(new_n477), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(G107), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT94), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n468), .A2(new_n203), .ZN(new_n483));
  INV_X1    g297(.A(new_n472), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n471), .A2(new_n252), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n476), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n188), .A2(G217), .A3(new_n304), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n488), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n189), .ZN(new_n492));
  INV_X1    g306(.A(G478), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(KEYINPUT15), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n492), .B(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n455), .A2(new_n463), .A3(new_n467), .A4(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G119), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n499), .A2(G128), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(KEYINPUT74), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(G128), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT23), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT73), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n500), .A2(new_n504), .A3(KEYINPUT23), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n222), .A2(G119), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT23), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT73), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n501), .A2(new_n503), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(G110), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n506), .A2(new_n502), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT24), .B(G110), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XOR2_X1   g328(.A(new_n514), .B(KEYINPUT75), .Z(new_n515));
  NAND2_X1  g329(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n408), .B1(new_n220), .B2(new_n404), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI221_X1 g332(.A(new_n434), .B1(new_n512), .B2(new_n513), .C1(new_n510), .C2(new_n509), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n308), .A2(G221), .A3(G234), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT22), .B(G137), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n521), .B(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n523), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n518), .A2(new_n519), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G217), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n528), .B1(G234), .B2(new_n189), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n529), .A2(G902), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT25), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n518), .A2(new_n519), .A3(new_n525), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n525), .B1(new_n518), .B2(new_n519), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n532), .B(new_n189), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n529), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n532), .B1(new_n527), .B2(new_n189), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n531), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(KEYINPUT76), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n266), .A2(new_n269), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT68), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n254), .A2(G134), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n256), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n541), .B1(new_n543), .B2(G131), .ZN(new_n544));
  AOI211_X1 g358(.A(KEYINPUT68), .B(new_n265), .C1(new_n542), .C2(new_n256), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n540), .A2(new_n241), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n282), .A2(new_n287), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n231), .A2(new_n288), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n547), .B(new_n342), .C1(new_n270), .C2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT70), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n267), .B(KEYINPUT66), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n265), .B1(new_n259), .B2(new_n260), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n289), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n556), .A2(KEYINPUT70), .A3(new_n342), .A4(new_n547), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n308), .A2(G210), .A3(new_n389), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(KEYINPUT27), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT26), .B(G101), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n560), .B(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT30), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n556), .A2(new_n563), .A3(new_n547), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n563), .B1(new_n556), .B2(new_n547), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n343), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n558), .A2(new_n562), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT31), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT31), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n558), .A2(new_n569), .A3(new_n566), .A4(new_n562), .ZN(new_n570));
  INV_X1    g384(.A(new_n551), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(KEYINPUT28), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n547), .B1(new_n270), .B2(new_n550), .ZN(new_n573));
  AOI21_X1  g387(.A(KEYINPUT72), .B1(new_n573), .B2(new_n343), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT72), .ZN(new_n575));
  AOI211_X1 g389(.A(new_n575), .B(new_n342), .C1(new_n556), .C2(new_n547), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n558), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n572), .B1(new_n577), .B2(KEYINPUT28), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n568), .B(new_n570), .C1(new_n578), .C2(new_n562), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT32), .ZN(new_n580));
  INV_X1    g394(.A(G472), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n579), .A2(new_n580), .A3(new_n581), .A4(new_n189), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n568), .A2(new_n570), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n576), .A2(new_n574), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n553), .A2(new_n557), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT28), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n572), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n562), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n581), .B(new_n189), .C1(new_n583), .C2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(KEYINPUT32), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n582), .A2(new_n590), .ZN(new_n591));
  OR2_X1    g405(.A1(new_n564), .A2(new_n565), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n585), .B1(new_n592), .B2(new_n343), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(new_n562), .ZN(new_n594));
  AOI211_X1 g408(.A(KEYINPUT29), .B(new_n594), .C1(new_n578), .C2(new_n562), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n573), .A2(new_n343), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT28), .B1(new_n585), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n587), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n562), .A2(KEYINPUT29), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n189), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(G472), .B1(new_n595), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n539), .B1(new_n591), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n384), .A2(new_n498), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  OAI211_X1 g419(.A(new_n325), .B(new_n463), .C1(new_n381), .C2(new_n382), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT76), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n538), .B(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n189), .B1(new_n583), .B2(new_n588), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(G472), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n609), .A2(new_n589), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n324), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n491), .A2(KEYINPUT33), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n489), .A2(new_n615), .A3(new_n490), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n189), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(G478), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n491), .A2(new_n493), .A3(new_n189), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n455), .B2(new_n467), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n607), .A2(new_n612), .A3(new_n613), .A4(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT34), .B(G104), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G6));
  AOI21_X1  g439(.A(new_n439), .B1(new_n453), .B2(new_n386), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n454), .B1(new_n626), .B2(KEYINPUT92), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n438), .A2(new_n385), .A3(new_n439), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n467), .B(new_n495), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT95), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n607), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n609), .A2(new_n589), .A3(new_n611), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(new_n324), .ZN(new_n634));
  OAI21_X1  g448(.A(KEYINPUT95), .B1(new_n606), .B2(new_n629), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n632), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT35), .B(G107), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G9));
  OR2_X1    g452(.A1(new_n536), .A2(new_n537), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n525), .A2(KEYINPUT36), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n520), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n530), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n611), .A2(new_n589), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(KEYINPUT96), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT96), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n611), .A2(new_n646), .A3(new_n589), .A4(new_n643), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n384), .A3(new_n498), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT37), .B(G110), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT97), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n649), .B(new_n651), .ZN(G12));
  NOR2_X1   g466(.A1(new_n460), .A2(G900), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n457), .B(KEYINPUT98), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n629), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n643), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n591), .B2(new_n602), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n384), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G128), .ZN(G30));
  INV_X1    g474(.A(new_n567), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n562), .B1(new_n558), .B2(new_n596), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n189), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(G472), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n664), .B(KEYINPUT99), .Z(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n591), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n325), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n667), .A2(new_n668), .A3(new_n643), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n372), .A2(new_n380), .ZN(new_n670));
  INV_X1    g484(.A(new_n373), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n372), .A2(new_n373), .A3(new_n380), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT38), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n467), .B1(new_n627), .B2(new_n628), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n496), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n669), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n655), .B(KEYINPUT39), .Z(new_n680));
  NAND2_X1  g494(.A1(new_n613), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT40), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(new_n230), .ZN(G45));
  AOI211_X1 g498(.A(new_n655), .B(new_n621), .C1(new_n467), .C2(new_n455), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n384), .A3(new_n658), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  AOI21_X1  g501(.A(new_n311), .B1(new_n315), .B2(new_n302), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n273), .A2(new_n311), .A3(new_n302), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n189), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(KEYINPUT100), .A2(G469), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n321), .A2(new_n322), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n189), .A3(new_n691), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n693), .A2(new_n695), .A3(new_n193), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT101), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n621), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n676), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n700), .A2(new_n606), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n698), .A2(new_n603), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT102), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT41), .B(G113), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G15));
  NAND4_X1  g519(.A1(new_n698), .A2(new_n632), .A3(new_n603), .A4(new_n635), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G116), .ZN(G18));
  NOR2_X1   g521(.A1(new_n676), .A2(new_n495), .ZN(new_n708));
  INV_X1    g522(.A(new_n696), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n658), .A2(new_n708), .A3(new_n607), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G119), .ZN(G21));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n611), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n610), .A2(KEYINPUT105), .A3(G472), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n581), .A2(new_n189), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT103), .ZN(new_n717));
  INV_X1    g531(.A(new_n562), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n599), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n568), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n570), .B1(new_n720), .B2(new_n721), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n717), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n538), .B(KEYINPUT106), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n715), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n668), .B1(new_n672), .B2(new_n673), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n729), .A2(new_n676), .A3(new_n495), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n698), .A2(new_n728), .A3(new_n463), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  INV_X1    g546(.A(new_n655), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n676), .A2(new_n699), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT107), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n383), .A2(new_n696), .A3(new_n657), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT107), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n622), .A2(new_n737), .A3(new_n733), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n723), .A2(new_n724), .ZN(new_n739));
  AOI22_X1  g553(.A1(new_n739), .A2(new_n717), .B1(new_n713), .B2(new_n714), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n735), .A2(new_n736), .A3(new_n738), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G125), .ZN(G27));
  AND4_X1   g556(.A1(new_n737), .A2(new_n676), .A3(new_n699), .A4(new_n733), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n737), .B1(new_n622), .B2(new_n733), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n672), .A2(new_n325), .A3(new_n673), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n324), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n591), .A2(new_n602), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n748), .A2(new_n726), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n745), .A2(KEYINPUT42), .A3(new_n747), .A4(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT42), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n735), .A2(new_n603), .A3(new_n738), .A4(new_n747), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n751), .B1(new_n752), .B2(KEYINPUT108), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n747), .A2(new_n603), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n754), .B1(new_n745), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n750), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI211_X1 g573(.A(KEYINPUT109), .B(new_n750), .C1(new_n753), .C2(new_n756), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G131), .ZN(G33));
  AND3_X1   g576(.A1(new_n747), .A2(new_n656), .A3(new_n603), .ZN(new_n763));
  XOR2_X1   g577(.A(KEYINPUT110), .B(G134), .Z(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(G36));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT43), .ZN(new_n767));
  AOI211_X1 g581(.A(new_n621), .B(new_n676), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n768), .B1(new_n766), .B2(new_n767), .ZN(new_n769));
  OAI211_X1 g583(.A(KEYINPUT111), .B(KEYINPUT43), .C1(new_n676), .C2(new_n621), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n657), .B1(new_n589), .B2(new_n611), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(KEYINPUT44), .A3(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n317), .B(KEYINPUT45), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(G469), .ZN(new_n778));
  NAND2_X1  g592(.A1(G469), .A2(G902), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(KEYINPUT46), .A3(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n323), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT46), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n782), .B(G469), .C1(new_n777), .C2(G902), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n193), .A3(new_n680), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(new_n746), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n773), .A2(new_n776), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G137), .ZN(G39));
  NOR4_X1   g602(.A1(new_n734), .A2(new_n748), .A3(new_n609), .A4(new_n746), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n784), .A2(KEYINPUT47), .A3(new_n193), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT47), .B1(new_n784), .B2(new_n193), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  NOR3_X1   g607(.A1(new_n666), .A2(new_n539), .A3(new_n458), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n746), .A2(new_n696), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n796), .A2(KEYINPUT117), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(KEYINPUT117), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n797), .A2(new_n677), .A3(new_n621), .A4(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n771), .A2(new_n654), .A3(new_n795), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n740), .A2(new_n643), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n790), .A2(new_n791), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n693), .A2(new_n695), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n803), .B1(new_n193), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n771), .A2(new_n654), .A3(new_n728), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n746), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n802), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n675), .A2(new_n325), .A3(new_n696), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(KEYINPUT50), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n808), .A2(new_n812), .A3(KEYINPUT51), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n797), .A2(new_n622), .A3(new_n798), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n456), .A2(G953), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n709), .A2(new_n729), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n814), .B(new_n815), .C1(new_n806), .C2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n749), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n800), .A2(new_n818), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n819), .A2(KEYINPUT48), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(KEYINPUT48), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n817), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n813), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT51), .B1(new_n808), .B2(new_n812), .ZN(new_n824));
  OR2_X1    g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n731), .A2(new_n706), .A3(new_n702), .A4(new_n710), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n497), .A2(new_n324), .A3(new_n383), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n603), .A2(new_n827), .B1(new_n701), .B2(new_n634), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT112), .B1(new_n607), .B2(new_n630), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT112), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n606), .A2(new_n629), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n634), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n828), .A2(new_n832), .A3(new_n649), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n747), .A2(new_n643), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n735), .A2(new_n740), .A3(new_n738), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n708), .A2(new_n748), .A3(new_n733), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n826), .A2(new_n833), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n763), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n759), .A2(new_n838), .A3(new_n760), .A4(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n643), .A2(new_n655), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT113), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n730), .A2(new_n613), .A3(new_n666), .A4(new_n843), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n384), .B(new_n658), .C1(new_n685), .C2(new_n656), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n741), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n741), .A2(new_n844), .A3(new_n845), .A4(KEYINPUT52), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OR2_X1    g666(.A1(new_n840), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT114), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n848), .A2(KEYINPUT114), .A3(new_n849), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT53), .B1(new_n840), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n853), .A2(new_n858), .A3(KEYINPUT54), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n851), .B1(new_n840), .B2(new_n857), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n839), .A2(new_n828), .A3(new_n832), .A4(new_n649), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n862), .A2(KEYINPUT115), .A3(new_n837), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT115), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n649), .A2(new_n604), .A3(new_n623), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n612), .A2(new_n613), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n607), .A2(new_n630), .A3(KEYINPUT112), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n830), .B1(new_n606), .B2(new_n629), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n865), .A2(new_n869), .A3(new_n763), .ZN(new_n870));
  INV_X1    g684(.A(new_n837), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n864), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n863), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n851), .B1(new_n848), .B2(new_n849), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT116), .ZN(new_n875));
  INV_X1    g689(.A(new_n826), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n757), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n875), .B1(new_n757), .B2(new_n876), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n873), .B(new_n874), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n860), .A2(new_n861), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n859), .A2(new_n880), .ZN(new_n881));
  OAI22_X1  g695(.A1(new_n825), .A2(new_n881), .B1(G952), .B2(G953), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n675), .A2(new_n676), .A3(new_n621), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n804), .B(KEYINPUT49), .Z(new_n884));
  AND3_X1   g698(.A1(new_n726), .A2(new_n193), .A3(new_n325), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n883), .A2(new_n667), .A3(new_n884), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n882), .A2(new_n886), .ZN(G75));
  NOR2_X1   g701(.A1(new_n308), .A2(G952), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n189), .B1(new_n860), .B2(new_n879), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT56), .B1(new_n890), .B2(G210), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n354), .A2(new_n361), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT118), .Z(new_n893));
  XNOR2_X1  g707(.A(new_n371), .B(KEYINPUT55), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n893), .B(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n889), .B1(new_n891), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT56), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n890), .A2(G210), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n898), .B1(new_n899), .B2(KEYINPUT119), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n899), .A2(KEYINPUT119), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n896), .B1(new_n900), .B2(new_n901), .ZN(G51));
  AOI211_X1 g716(.A(KEYINPUT120), .B(new_n861), .C1(new_n860), .C2(new_n879), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n861), .B1(new_n860), .B2(new_n879), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT120), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n880), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n903), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n779), .B(KEYINPUT57), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n694), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n890), .A2(G469), .A3(new_n777), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n888), .B1(new_n910), .B2(new_n911), .ZN(G54));
  NAND2_X1  g726(.A1(KEYINPUT58), .A2(G475), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT121), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n890), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n889), .B1(new_n915), .B2(new_n453), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n453), .B2(new_n915), .ZN(G60));
  NAND2_X1  g731(.A1(G478), .A2(G902), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT59), .Z(new_n919));
  AOI21_X1  g733(.A(new_n919), .B1(new_n859), .B2(new_n880), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n889), .B1(new_n920), .B2(new_n617), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT122), .ZN(new_n922));
  INV_X1    g736(.A(new_n617), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n923), .A2(new_n919), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n922), .B1(new_n908), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n904), .B1(new_n906), .B2(new_n880), .ZN(new_n927));
  OAI211_X1 g741(.A(KEYINPUT122), .B(new_n924), .C1(new_n927), .C2(new_n903), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n921), .B1(new_n926), .B2(new_n928), .ZN(G63));
  NAND2_X1  g743(.A1(new_n860), .A2(new_n879), .ZN(new_n930));
  OAI21_X1  g744(.A(KEYINPUT60), .B1(new_n528), .B2(new_n189), .ZN(new_n931));
  OR3_X1    g745(.A1(new_n528), .A2(new_n189), .A3(KEYINPUT60), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n527), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n930), .A2(new_n641), .A3(new_n931), .A4(new_n932), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n935), .A2(new_n889), .A3(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(G66));
  OAI21_X1  g753(.A(G953), .B1(new_n461), .B2(new_n367), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n826), .A2(new_n833), .ZN(new_n941));
  INV_X1    g755(.A(new_n308), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n893), .B1(G898), .B2(new_n308), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(G69));
  OAI211_X1 g759(.A(new_n755), .B(new_n680), .C1(new_n622), .C2(new_n630), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n787), .A2(new_n792), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n741), .A2(new_n845), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n683), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT62), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT123), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n947), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n951), .B1(new_n947), .B2(new_n950), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n592), .B(new_n409), .Z(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n749), .A2(new_n730), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n785), .A2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n948), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n787), .A2(KEYINPUT124), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT124), .B1(new_n787), .B2(new_n960), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n792), .B(new_n959), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n761), .A2(new_n839), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n956), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n308), .B1(new_n957), .B2(new_n966), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n956), .A2(G227), .ZN(new_n968));
  OAI21_X1  g782(.A(G900), .B1(new_n956), .B2(G227), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n942), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n967), .A2(new_n970), .ZN(G72));
  NOR2_X1   g785(.A1(new_n593), .A2(new_n718), .ZN(new_n972));
  INV_X1    g786(.A(new_n941), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n952), .A2(new_n953), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(G472), .A2(G902), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT63), .Z(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT125), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n972), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n594), .A2(new_n661), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n853), .A2(new_n858), .A3(new_n976), .A4(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n978), .A2(new_n889), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n593), .A2(new_n718), .ZN(new_n982));
  INV_X1    g796(.A(new_n977), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n964), .A2(new_n941), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n983), .B1(new_n963), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(KEYINPUT126), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT126), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n987), .B(new_n983), .C1(new_n963), .C2(new_n984), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n982), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n981), .A2(new_n989), .ZN(G57));
endmodule


