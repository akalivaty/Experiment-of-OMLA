//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070;
  XNOR2_X1  g000(.A(G125), .B(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT16), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NOR3_X1   g003(.A1(new_n189), .A2(KEYINPUT16), .A3(G140), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n188), .A2(G146), .A3(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G140), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G125), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n189), .A2(G140), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n198));
  INV_X1    g012(.A(G119), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G128), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT23), .A3(G119), .ZN(new_n202));
  INV_X1    g016(.A(G110), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(G128), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n200), .A2(new_n202), .A3(new_n203), .A4(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT74), .ZN(new_n206));
  XOR2_X1   g020(.A(KEYINPUT24), .B(G110), .Z(new_n207));
  XNOR2_X1  g021(.A(G119), .B(G128), .ZN(new_n208));
  OAI22_X1  g022(.A1(new_n205), .A2(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AND2_X1   g023(.A1(new_n205), .A2(new_n206), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n192), .B(new_n197), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n200), .A2(new_n204), .A3(new_n202), .ZN(new_n212));
  AOI22_X1  g026(.A1(G110), .A2(new_n212), .B1(new_n207), .B2(new_n208), .ZN(new_n213));
  AOI211_X1 g027(.A(new_n196), .B(new_n190), .C1(KEYINPUT16), .C2(new_n187), .ZN(new_n214));
  AOI21_X1  g028(.A(G146), .B1(new_n188), .B2(new_n191), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT22), .B(G137), .ZN(new_n218));
  INV_X1    g032(.A(G953), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(G221), .A3(G234), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n218), .B(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n211), .A2(new_n216), .A3(new_n221), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g039(.A(KEYINPUT71), .B(G902), .Z(new_n226));
  OAI21_X1  g040(.A(KEYINPUT25), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT25), .ZN(new_n228));
  INV_X1    g042(.A(new_n226), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n223), .A2(new_n228), .A3(new_n229), .A4(new_n224), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT72), .B(G217), .ZN(new_n231));
  INV_X1    g045(.A(G234), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n231), .B1(new_n226), .B2(new_n232), .ZN(new_n233));
  XOR2_X1   g047(.A(new_n233), .B(KEYINPUT73), .Z(new_n234));
  AND2_X1   g048(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n225), .A2(KEYINPUT75), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT75), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n223), .A2(new_n237), .A3(new_n224), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n234), .A2(G902), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n227), .A2(new_n235), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G116), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT67), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G116), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n244), .A2(new_n246), .A3(G119), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n243), .A2(G119), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G113), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT2), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT2), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G113), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n247), .A2(new_n249), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n254), .B1(new_n247), .B2(new_n249), .ZN(new_n256));
  OR2_X1    g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G137), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT66), .A3(G134), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT66), .ZN(new_n260));
  INV_X1    g074(.A(G134), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n260), .B1(new_n261), .B2(G137), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n258), .A2(G134), .ZN(new_n263));
  OAI211_X1 g077(.A(G131), .B(new_n259), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT11), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n265), .B1(new_n261), .B2(G137), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n258), .A2(KEYINPUT11), .A3(G134), .ZN(new_n267));
  INV_X1    g081(.A(G131), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n261), .A2(G137), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n266), .A2(new_n267), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n196), .A2(G143), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n201), .B1(new_n272), .B2(KEYINPUT1), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT65), .B1(new_n196), .B2(G143), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT65), .ZN(new_n275));
  INV_X1    g089(.A(G143), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n276), .A3(G146), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(KEYINPUT64), .A2(G143), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(KEYINPUT64), .A2(G143), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n196), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n273), .B1(new_n278), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT64), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n276), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(G146), .A3(new_n279), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n272), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n271), .B1(new_n283), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n266), .A2(new_n267), .A3(new_n269), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(G131), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n270), .ZN(new_n293));
  AND2_X1   g107(.A1(KEYINPUT0), .A2(G128), .ZN(new_n294));
  NOR2_X1   g108(.A1(KEYINPUT0), .A2(G128), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(G146), .B1(new_n285), .B2(new_n279), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n274), .A2(new_n277), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n286), .A2(new_n272), .A3(new_n294), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n293), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT30), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n290), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n302), .B1(new_n290), .B2(new_n301), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n257), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT31), .ZN(new_n306));
  INV_X1    g120(.A(G237), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(new_n219), .A3(G210), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n308), .B(KEYINPUT27), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT26), .B(G101), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n309), .B(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n255), .A2(new_n256), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n290), .A2(new_n301), .A3(new_n312), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n305), .A2(new_n306), .A3(new_n311), .A4(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT28), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n293), .A2(new_n299), .A3(new_n300), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n264), .A2(new_n270), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n272), .A2(KEYINPUT1), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G128), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n319), .B1(new_n297), .B2(new_n298), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n317), .B1(new_n288), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n257), .B1(new_n316), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n315), .B1(new_n322), .B2(new_n313), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT69), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n313), .A2(new_n324), .A3(new_n315), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n324), .B1(new_n313), .B2(new_n315), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n314), .B1(new_n327), .B2(new_n311), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n305), .A2(new_n311), .A3(new_n313), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT31), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT68), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n329), .A2(KEYINPUT68), .A3(KEYINPUT31), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n328), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(G472), .A2(G902), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(KEYINPUT32), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT30), .B1(new_n316), .B2(new_n321), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n290), .A2(new_n301), .A3(new_n302), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n312), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n311), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n290), .A2(new_n301), .A3(new_n312), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n312), .B1(new_n290), .B2(new_n301), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT28), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n313), .A2(new_n315), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT69), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n313), .A2(new_n324), .A3(new_n315), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n345), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n343), .A2(new_n306), .B1(new_n349), .B2(new_n341), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n329), .A2(KEYINPUT68), .A3(KEYINPUT31), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT68), .B1(new_n329), .B2(KEYINPUT31), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT32), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(new_n335), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n337), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n311), .B1(new_n305), .B2(new_n313), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n357), .A2(KEYINPUT29), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n345), .A2(new_n347), .A3(new_n311), .A4(new_n348), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n226), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT29), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n362), .A2(KEYINPUT70), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT70), .ZN(new_n364));
  NOR3_X1   g178(.A1(new_n359), .A2(new_n364), .A3(new_n361), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n360), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G472), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n242), .B1(new_n356), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(G210), .B1(G237), .B2(G902), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n369), .B(KEYINPUT82), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT76), .ZN(new_n371));
  XNOR2_X1  g185(.A(G104), .B(G107), .ZN(new_n372));
  INV_X1    g186(.A(G101), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G104), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT3), .B1(new_n375), .B2(G107), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT3), .ZN(new_n377));
  INV_X1    g191(.A(G107), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(G104), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n375), .A2(G107), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n376), .A2(new_n379), .A3(new_n373), .A4(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n375), .A2(G107), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n378), .A2(G104), .ZN(new_n383));
  OAI211_X1 g197(.A(KEYINPUT76), .B(G101), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n374), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(KEYINPUT67), .B(G116), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n248), .B1(new_n386), .B2(G119), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n254), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n247), .A2(KEYINPUT5), .A3(new_n249), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT5), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n250), .B1(new_n248), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n385), .A2(new_n388), .A3(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(G110), .B(G122), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n376), .A2(new_n379), .A3(new_n380), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G101), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n396), .A2(KEYINPUT4), .A3(new_n381), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT4), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n395), .A2(new_n398), .A3(G101), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(new_n255), .B2(new_n256), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n393), .B(new_n394), .C1(new_n397), .C2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(KEYINPUT79), .B(G224), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n219), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT7), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n320), .A2(new_n189), .A3(new_n288), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n189), .B1(new_n299), .B2(new_n300), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT80), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n394), .B(KEYINPUT8), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n389), .A2(new_n391), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n374), .A2(new_n381), .A3(new_n384), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n410), .A2(new_n411), .A3(new_n255), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n374), .A2(new_n384), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n413), .A2(new_n381), .B1(new_n392), .B2(new_n388), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n409), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n406), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n320), .A2(new_n189), .A3(new_n288), .ZN(new_n417));
  INV_X1    g231(.A(new_n404), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT80), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n420), .B(new_n404), .C1(new_n405), .C2(new_n406), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n408), .A2(new_n415), .A3(new_n419), .A4(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n401), .B1(new_n422), .B2(KEYINPUT81), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT81), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n418), .B1(new_n416), .B2(new_n417), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n411), .B1(new_n410), .B2(new_n255), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n393), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n425), .A2(new_n420), .B1(new_n427), .B2(new_n409), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n405), .A2(new_n406), .A3(new_n404), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(KEYINPUT80), .B2(new_n407), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n424), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n423), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n394), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n400), .A2(new_n397), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n433), .B1(new_n434), .B2(new_n412), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(KEYINPUT6), .A3(new_n401), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n219), .B(new_n402), .C1(new_n405), .C2(new_n406), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n416), .A2(new_n417), .A3(new_n403), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT6), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n440), .B(new_n433), .C1(new_n434), .C2(new_n412), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n436), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G902), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n370), .B1(new_n432), .B2(new_n444), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n442), .A2(new_n443), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n422), .A2(KEYINPUT81), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n428), .A2(new_n430), .A3(new_n424), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n448), .A3(new_n401), .ZN(new_n449));
  INV_X1    g263(.A(new_n370), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n446), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n445), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(G110), .B(G140), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n219), .A2(G227), .ZN(new_n454));
  XOR2_X1   g268(.A(new_n453), .B(new_n454), .Z(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n286), .A2(new_n272), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT1), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT64), .B(G143), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n458), .B1(new_n459), .B2(new_n196), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n457), .B1(new_n460), .B2(new_n201), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT77), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n286), .A2(new_n462), .A3(new_n272), .A4(new_n287), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n288), .A2(KEYINPUT77), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n461), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n385), .ZN(new_n466));
  XOR2_X1   g280(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n293), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n299), .A2(new_n399), .A3(new_n300), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n396), .A2(KEYINPUT4), .A3(new_n381), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT10), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n473), .B1(new_n320), .B2(new_n288), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n471), .A2(new_n472), .B1(new_n474), .B2(new_n385), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n468), .A2(new_n469), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n411), .A2(new_n288), .A3(new_n320), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n466), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(KEYINPUT12), .B1(new_n478), .B2(new_n293), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT12), .ZN(new_n480));
  AOI211_X1 g294(.A(new_n480), .B(new_n469), .C1(new_n466), .C2(new_n477), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n456), .B(new_n476), .C1(new_n479), .C2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n469), .B1(new_n468), .B2(new_n475), .ZN(new_n483));
  INV_X1    g297(.A(new_n467), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n484), .B1(new_n465), .B2(new_n385), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT10), .B1(new_n283), .B2(new_n289), .ZN(new_n486));
  OAI22_X1  g300(.A1(new_n486), .A2(new_n411), .B1(new_n397), .B2(new_n470), .ZN(new_n487));
  NOR3_X1   g301(.A1(new_n485), .A2(new_n487), .A3(new_n293), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n455), .B1(new_n483), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n482), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G469), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n229), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n491), .A2(new_n443), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n293), .B1(new_n485), .B2(new_n487), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n476), .A2(new_n495), .A3(new_n456), .ZN(new_n496));
  OAI21_X1  g310(.A(G128), .B1(new_n297), .B2(new_n458), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n497), .A2(new_n457), .B1(new_n288), .B2(KEYINPUT77), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n411), .B1(new_n498), .B2(new_n463), .ZN(new_n499));
  INV_X1    g313(.A(new_n477), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n293), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n480), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n478), .A2(KEYINPUT12), .A3(new_n293), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n485), .A2(new_n487), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n502), .A2(new_n503), .B1(new_n504), .B2(new_n469), .ZN(new_n505));
  OAI211_X1 g319(.A(G469), .B(new_n496), .C1(new_n505), .C2(new_n456), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n492), .A2(new_n494), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(G214), .B1(G237), .B2(G902), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT9), .B(G234), .ZN(new_n509));
  OAI21_X1  g323(.A(G221), .B1(new_n509), .B2(G902), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n452), .A2(new_n507), .A3(new_n508), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(KEYINPUT18), .A2(G131), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n307), .A2(new_n219), .A3(G214), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n285), .A3(new_n279), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n307), .A2(new_n219), .A3(G143), .A4(G214), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n515), .A2(KEYINPUT83), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(KEYINPUT83), .B1(new_n515), .B2(new_n516), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n513), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(G214), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n520), .A2(G237), .A3(G953), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n512), .B(new_n516), .C1(new_n459), .C2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT85), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT85), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n515), .A2(new_n524), .A3(new_n512), .A4(new_n516), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n197), .A2(KEYINPUT84), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n194), .A2(new_n195), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(G146), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n528), .A2(KEYINPUT84), .A3(G146), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n519), .A2(new_n526), .A3(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n214), .A2(new_n215), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n516), .B1(new_n459), .B2(new_n521), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(G131), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT17), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n515), .A2(new_n268), .A3(new_n516), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n535), .A2(KEYINPUT17), .A3(G131), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n534), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(G113), .B(G122), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(G104), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(KEYINPUT88), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n533), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n543), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n533), .A2(new_n541), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT89), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n533), .A2(new_n541), .A3(KEYINPUT89), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n546), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(G475), .B1(new_n552), .B2(G902), .ZN(new_n553));
  NOR2_X1   g367(.A1(G475), .A2(G902), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(KEYINPUT86), .A2(KEYINPUT19), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n194), .A2(new_n195), .A3(new_n556), .ZN(new_n557));
  XOR2_X1   g371(.A(KEYINPUT86), .B(KEYINPUT19), .Z(new_n558));
  OAI211_X1 g372(.A(new_n196), .B(new_n557), .C1(new_n558), .C2(new_n187), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n559), .A2(new_n192), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n536), .A2(new_n538), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n533), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT87), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n533), .A2(KEYINPUT87), .A3(new_n562), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n543), .A3(new_n566), .ZN(new_n567));
  AOI211_X1 g381(.A(KEYINPUT20), .B(new_n555), .C1(new_n567), .C2(new_n545), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT20), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n523), .A2(new_n525), .B1(new_n530), .B2(new_n531), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n570), .A2(new_n519), .B1(new_n560), .B2(new_n561), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n543), .B1(new_n571), .B2(KEYINPUT87), .ZN(new_n572));
  INV_X1    g386(.A(new_n566), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n545), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n569), .B1(new_n574), .B2(new_n554), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n553), .B1(new_n568), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT90), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n276), .A2(G128), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n580), .B1(new_n459), .B2(new_n201), .ZN(new_n581));
  OAI21_X1  g395(.A(G134), .B1(new_n579), .B2(KEYINPUT13), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n581), .B(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT91), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n244), .A2(new_n246), .A3(G122), .ZN(new_n585));
  INV_X1    g399(.A(G122), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(G116), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n584), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n585), .A2(new_n584), .A3(new_n587), .ZN(new_n590));
  AOI21_X1  g404(.A(G107), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n590), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n592), .A2(new_n588), .A3(new_n378), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n583), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n581), .B(G134), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n378), .B1(new_n592), .B2(new_n588), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT92), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT14), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n587), .A2(new_n598), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n585), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n597), .B1(new_n585), .B2(new_n599), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n585), .A2(KEYINPUT14), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n595), .B(new_n596), .C1(new_n603), .C2(new_n378), .ZN(new_n604));
  INV_X1    g418(.A(new_n509), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(new_n219), .A3(new_n231), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n594), .A2(new_n604), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n607), .B1(new_n594), .B2(new_n604), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n229), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(G478), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(KEYINPUT15), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n594), .A2(new_n604), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n606), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n226), .B1(new_n616), .B2(new_n608), .ZN(new_n617));
  INV_X1    g431(.A(new_n613), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n219), .A2(G952), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(G234), .B2(G237), .ZN(new_n622));
  AOI211_X1 g436(.A(new_n219), .B(new_n229), .C1(G234), .C2(G237), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT21), .B(G898), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n553), .B(KEYINPUT90), .C1(new_n568), .C2(new_n575), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n578), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n511), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n368), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G101), .ZN(G3));
  OAI21_X1  g445(.A(KEYINPUT33), .B1(new_n609), .B2(new_n610), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT33), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n616), .A2(new_n633), .A3(new_n608), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n226), .A2(new_n612), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n635), .A2(new_n636), .B1(new_n612), .B2(new_n611), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n627), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n547), .B1(new_n563), .B2(new_n564), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n546), .B1(new_n640), .B2(new_n566), .ZN(new_n641));
  OAI21_X1  g455(.A(KEYINPUT20), .B1(new_n641), .B2(new_n555), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n574), .A2(new_n569), .A3(new_n554), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT90), .B1(new_n644), .B2(new_n553), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n638), .B1(new_n639), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n625), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n432), .A2(new_n444), .A3(new_n370), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n450), .B1(new_n446), .B2(new_n449), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n647), .B(new_n508), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n506), .A2(new_n494), .ZN(new_n653));
  AOI211_X1 g467(.A(G469), .B(new_n226), .C1(new_n482), .C2(new_n489), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n241), .B(new_n510), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n334), .A2(new_n336), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n353), .A2(KEYINPUT93), .A3(new_n229), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(G472), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n332), .A2(new_n333), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n226), .B1(new_n661), .B2(new_n350), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(KEYINPUT93), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n656), .B(new_n658), .C1(new_n660), .C2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n652), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT34), .B(G104), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G6));
  INV_X1    g481(.A(new_n664), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT94), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n642), .A2(new_n643), .A3(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n669), .B1(new_n642), .B2(new_n643), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n553), .B(new_n620), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n650), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n668), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT35), .B(G107), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G9));
  INV_X1    g491(.A(G472), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n678), .B1(new_n662), .B2(KEYINPUT93), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n353), .A2(new_n229), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT93), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n657), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  OR3_X1    g497(.A1(new_n217), .A2(KEYINPUT36), .A3(new_n222), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n217), .B1(KEYINPUT36), .B2(new_n222), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n684), .A2(new_n240), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n686), .B1(new_n235), .B2(new_n227), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n683), .A2(new_n629), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT37), .B(G110), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT95), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n689), .B(new_n691), .ZN(G12));
  XOR2_X1   g506(.A(new_n622), .B(KEYINPUT96), .Z(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(G900), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n694), .B1(new_n695), .B2(new_n623), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n673), .A2(new_n696), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n353), .A2(new_n354), .A3(new_n335), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n354), .B1(new_n353), .B2(new_n335), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n367), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n508), .B1(new_n648), .B2(new_n649), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n510), .B1(new_n653), .B2(new_n654), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n697), .A2(new_n700), .A3(new_n703), .A4(new_n688), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G128), .ZN(G30));
  XOR2_X1   g519(.A(new_n696), .B(KEYINPUT39), .Z(new_n706));
  NAND3_X1  g520(.A1(new_n507), .A2(new_n510), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT40), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT97), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT38), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n452), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n445), .A2(KEYINPUT38), .A3(new_n451), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n639), .A2(new_n645), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n305), .A2(new_n313), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n311), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n342), .A2(new_n344), .ZN(new_n720));
  AOI21_X1  g534(.A(G902), .B1(new_n720), .B2(new_n341), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n678), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n723), .B1(new_n698), .B2(new_n699), .ZN(new_n724));
  INV_X1    g538(.A(new_n620), .ZN(new_n725));
  INV_X1    g539(.A(new_n508), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n725), .A2(new_n688), .A3(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n715), .A2(new_n717), .A3(new_n724), .A4(new_n727), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n710), .A2(new_n711), .A3(new_n728), .ZN(new_n729));
  XOR2_X1   g543(.A(new_n729), .B(new_n459), .Z(G45));
  AOI211_X1 g544(.A(new_n637), .B(new_n696), .C1(new_n578), .C2(new_n627), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n731), .A2(new_n700), .A3(new_n703), .A4(new_n688), .ZN(new_n732));
  XOR2_X1   g546(.A(KEYINPUT98), .B(G146), .Z(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G48));
  NOR2_X1   g548(.A1(new_n488), .A2(new_n455), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n502), .A2(new_n503), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n476), .A2(new_n495), .ZN(new_n737));
  AOI22_X1  g551(.A1(new_n735), .A2(new_n736), .B1(new_n737), .B2(new_n455), .ZN(new_n738));
  OAI21_X1  g552(.A(G469), .B1(new_n738), .B2(new_n226), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n739), .A2(new_n510), .A3(new_n492), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n651), .A2(new_n700), .A3(new_n241), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(KEYINPUT41), .B(G113), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G15));
  NAND4_X1  g557(.A1(new_n674), .A2(new_n700), .A3(new_n241), .A4(new_n740), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT99), .B(G116), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G18));
  INV_X1    g560(.A(new_n628), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n739), .A2(new_n492), .A3(new_n510), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n701), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n700), .A2(new_n747), .A3(new_n749), .A4(new_n688), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G119), .ZN(G21));
  NAND2_X1  g565(.A1(new_n349), .A2(new_n341), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n330), .A3(new_n314), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n335), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT100), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT100), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n753), .A2(new_n756), .A3(new_n335), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n678), .B1(new_n353), .B2(new_n229), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n758), .A2(new_n759), .A3(new_n242), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n726), .B1(new_n445), .B2(new_n451), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n725), .B1(new_n578), .B2(new_n627), .ZN(new_n762));
  AND4_X1   g576(.A1(new_n647), .A2(new_n739), .A3(new_n510), .A4(new_n492), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n760), .A2(new_n761), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G122), .ZN(G24));
  NOR3_X1   g579(.A1(new_n758), .A2(new_n759), .A3(new_n687), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n731), .A3(new_n749), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G125), .ZN(G27));
  INV_X1    g582(.A(KEYINPUT42), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n445), .A2(new_n508), .A3(new_n451), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT101), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n770), .B1(new_n702), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n507), .A2(KEYINPUT101), .A3(new_n510), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n700), .A2(new_n772), .A3(new_n241), .A4(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n731), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n769), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n702), .A2(new_n771), .ZN(new_n777));
  INV_X1    g591(.A(new_n770), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n778), .A3(new_n773), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n780), .A2(new_n368), .A3(KEYINPUT42), .A4(new_n731), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n776), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G131), .ZN(G33));
  NAND3_X1  g597(.A1(new_n780), .A2(new_n368), .A3(new_n697), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G134), .ZN(G36));
  OAI21_X1  g599(.A(new_n496), .B1(new_n505), .B2(new_n456), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n491), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI211_X1 g602(.A(KEYINPUT45), .B(new_n496), .C1(new_n505), .C2(new_n456), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n493), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n492), .B1(new_n790), .B2(KEYINPUT46), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n788), .A2(new_n789), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n792), .A2(KEYINPUT46), .A3(new_n494), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n510), .B(new_n706), .C1(new_n791), .C2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n578), .A2(new_n627), .A3(new_n638), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT43), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n578), .A2(new_n638), .A3(KEYINPUT43), .A4(new_n627), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n682), .A2(G472), .A3(new_n659), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n658), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n799), .A2(new_n801), .A3(new_n688), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT44), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n794), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n804), .B(new_n778), .C1(new_n803), .C2(new_n802), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G137), .ZN(G39));
  OAI21_X1  g620(.A(new_n510), .B1(new_n791), .B2(new_n793), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT47), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI211_X1 g623(.A(KEYINPUT47), .B(new_n510), .C1(new_n791), .C2(new_n793), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n700), .A2(new_n241), .A3(new_n770), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(new_n731), .A3(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G140), .ZN(G42));
  AOI21_X1  g628(.A(new_n722), .B1(new_n337), .B2(new_n355), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n241), .A2(new_n622), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n770), .A2(new_n748), .A3(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n646), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n621), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n740), .A2(new_n761), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n693), .B1(new_n797), .B2(new_n798), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n760), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n778), .A2(new_n740), .ZN(new_n824));
  AOI211_X1 g638(.A(new_n693), .B(new_n824), .C1(new_n797), .C2(new_n798), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n368), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n826), .A2(KEYINPUT48), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(KEYINPUT48), .ZN(new_n828));
  OAI221_X1 g642(.A(new_n820), .B1(new_n821), .B2(new_n823), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n739), .A2(new_n492), .A3(new_n726), .A4(new_n510), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n830), .B1(new_n713), .B2(new_n714), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n799), .A2(new_n694), .A3(new_n760), .A4(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT50), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n822), .A2(KEYINPUT50), .A3(new_n760), .A4(new_n831), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AND4_X1   g650(.A1(new_n716), .A2(new_n815), .A3(new_n817), .A4(new_n637), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n837), .B1(new_n825), .B2(new_n766), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT108), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n836), .A2(new_n838), .A3(KEYINPUT108), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT107), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n843), .B1(new_n823), .B2(new_n770), .ZN(new_n844));
  INV_X1    g658(.A(new_n510), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n739), .A2(new_n492), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n809), .A2(new_n810), .A3(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n822), .A2(KEYINPUT107), .A3(new_n760), .A4(new_n778), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n844), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n841), .A2(new_n842), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n829), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT109), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n836), .A2(new_n853), .A3(new_n838), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n853), .B1(new_n836), .B2(new_n838), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT110), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n847), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n809), .A2(KEYINPUT110), .A3(new_n810), .A4(new_n846), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n858), .A2(new_n859), .A3(new_n844), .A4(new_n848), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT51), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT111), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n856), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n860), .A2(KEYINPUT51), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n839), .A2(KEYINPUT109), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n836), .A2(new_n838), .A3(new_n853), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT111), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n852), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT112), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n872));
  AND4_X1   g686(.A1(new_n741), .A2(new_n744), .A3(new_n750), .A4(new_n764), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n872), .B1(new_n873), .B2(KEYINPUT105), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n578), .A2(new_n627), .A3(new_n620), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n650), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n876), .A2(new_n658), .A3(new_n800), .A4(new_n656), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n689), .A2(KEYINPUT102), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT102), .B1(new_n689), .B2(new_n877), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n630), .B1(new_n652), .B2(new_n664), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n741), .A2(new_n744), .A3(new_n750), .A4(new_n764), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT105), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n874), .A2(new_n881), .A3(new_n782), .A4(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT103), .ZN(new_n886));
  INV_X1    g700(.A(new_n696), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n614), .A2(new_n619), .A3(new_n887), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n888), .A2(new_n687), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n702), .A2(new_n770), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n672), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n670), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n892), .A2(new_n553), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n890), .A2(new_n893), .A3(new_n700), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n766), .A2(new_n731), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n894), .B1(new_n895), .B2(new_n779), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n700), .A2(new_n241), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n892), .A2(new_n553), .A3(new_n620), .A4(new_n887), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n897), .A2(new_n779), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n886), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n687), .A2(new_n887), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n724), .A2(new_n703), .A3(new_n762), .A4(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n704), .A2(new_n732), .A3(new_n767), .A4(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT52), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n780), .A2(new_n731), .A3(new_n766), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n784), .A2(new_n906), .A3(KEYINPUT103), .A4(new_n894), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n687), .B1(new_n356), .B2(new_n367), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n908), .B(new_n703), .C1(new_n697), .C2(new_n731), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT52), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n909), .A2(new_n910), .A3(new_n767), .A4(new_n903), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n900), .A2(new_n905), .A3(new_n907), .A4(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(KEYINPUT106), .B1(new_n885), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT54), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n878), .A2(new_n880), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n747), .A2(new_n703), .A3(new_n688), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n716), .A2(new_n647), .A3(new_n620), .A4(new_n761), .ZN(new_n917));
  OAI22_X1  g731(.A1(new_n916), .A2(new_n801), .B1(new_n664), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT102), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n915), .A2(new_n782), .A3(new_n920), .A4(new_n873), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n872), .B1(new_n921), .B2(new_n912), .ZN(new_n922));
  AND4_X1   g736(.A1(new_n905), .A2(new_n900), .A3(new_n911), .A4(new_n907), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n716), .A2(new_n725), .A3(new_n701), .ZN(new_n924));
  INV_X1    g738(.A(new_n759), .ZN(new_n925));
  INV_X1    g739(.A(new_n757), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n756), .B1(new_n753), .B2(new_n335), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AND4_X1   g742(.A1(new_n241), .A2(new_n925), .A3(new_n928), .A4(new_n763), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n821), .A2(new_n628), .ZN(new_n930));
  AOI22_X1  g744(.A1(new_n924), .A2(new_n929), .B1(new_n908), .B2(new_n930), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n931), .A2(KEYINPUT105), .A3(new_n741), .A4(new_n744), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n884), .A2(new_n932), .A3(KEYINPUT53), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT106), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n689), .A2(new_n877), .A3(KEYINPUT102), .ZN(new_n935));
  AOI22_X1  g749(.A1(new_n668), .A2(new_n651), .B1(new_n368), .B2(new_n629), .ZN(new_n936));
  AND4_X1   g750(.A1(new_n782), .A2(new_n920), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n923), .A2(new_n933), .A3(new_n934), .A4(new_n937), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n913), .A2(new_n914), .A3(new_n922), .A4(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n782), .A2(new_n920), .A3(new_n935), .A4(new_n936), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n940), .A2(new_n882), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n905), .A2(KEYINPUT104), .A3(new_n911), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n872), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n941), .A2(new_n923), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n943), .B1(new_n941), .B2(new_n923), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT54), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n939), .A2(new_n946), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n852), .B(KEYINPUT112), .C1(new_n863), .C2(new_n868), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n871), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(KEYINPUT113), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT113), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n871), .A2(new_n947), .A3(new_n951), .A4(new_n948), .ZN(new_n952));
  OR2_X1    g766(.A1(G952), .A2(G953), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n950), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n739), .A2(new_n492), .ZN(new_n955));
  OR2_X1    g769(.A1(new_n955), .A2(KEYINPUT49), .ZN(new_n956));
  NOR4_X1   g770(.A1(new_n242), .A2(new_n637), .A3(new_n726), .A4(new_n845), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n955), .A2(KEYINPUT49), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  OR4_X1    g773(.A1(new_n717), .A2(new_n959), .A3(new_n715), .A4(new_n724), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n954), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT114), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n954), .A2(KEYINPUT114), .A3(new_n960), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(G75));
  NOR2_X1   g779(.A1(new_n219), .A2(G952), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n913), .A2(new_n922), .A3(new_n938), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n226), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(KEYINPUT56), .B1(new_n970), .B2(new_n370), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n436), .A2(new_n441), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(new_n439), .Z(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT55), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n967), .B1(new_n971), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n971), .B2(new_n975), .ZN(G51));
  NAND2_X1  g791(.A1(new_n968), .A2(KEYINPUT54), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n939), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n493), .B(KEYINPUT115), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT57), .Z(new_n981));
  AOI21_X1  g795(.A(new_n738), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  OR2_X1    g796(.A1(new_n982), .A2(KEYINPUT116), .ZN(new_n983));
  INV_X1    g797(.A(new_n792), .ZN(new_n984));
  AOI22_X1  g798(.A1(new_n982), .A2(KEYINPUT116), .B1(new_n984), .B2(new_n970), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n966), .B1(new_n983), .B2(new_n985), .ZN(G54));
  AND2_X1   g800(.A1(KEYINPUT58), .A2(G475), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n970), .A2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n989), .A2(KEYINPUT117), .A3(new_n574), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n967), .B1(new_n989), .B2(new_n574), .ZN(new_n991));
  AOI21_X1  g805(.A(KEYINPUT117), .B1(new_n989), .B2(new_n574), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(G60));
  NAND2_X1  g807(.A1(G478), .A2(G902), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT59), .Z(new_n995));
  NOR2_X1   g809(.A1(new_n947), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n996), .A2(new_n635), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n995), .B1(new_n632), .B2(new_n634), .ZN(new_n998));
  AOI211_X1 g812(.A(new_n966), .B(new_n997), .C1(new_n979), .C2(new_n998), .ZN(G63));
  NAND2_X1  g813(.A1(G217), .A2(G902), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(KEYINPUT118), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(KEYINPUT60), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n938), .A2(new_n922), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n884), .A2(new_n932), .A3(KEYINPUT53), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n1004), .A2(new_n940), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n934), .B1(new_n1005), .B2(new_n923), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1002), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(new_n239), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  AND2_X1   g823(.A1(new_n684), .A2(new_n685), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n968), .A2(new_n1010), .A3(new_n1002), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n1009), .A2(KEYINPUT61), .A3(new_n967), .A4(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT120), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n966), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n1015), .A2(KEYINPUT120), .A3(KEYINPUT61), .A4(new_n1011), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  AOI211_X1 g831(.A(KEYINPUT119), .B(KEYINPUT61), .C1(new_n1015), .C2(new_n1011), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT119), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1015), .A2(new_n1011), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT61), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1019), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1017), .B1(new_n1018), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT121), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI211_X1 g839(.A(new_n1017), .B(KEYINPUT121), .C1(new_n1018), .C2(new_n1022), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1025), .A2(new_n1026), .ZN(G66));
  INV_X1    g841(.A(new_n624), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n219), .B1(new_n1028), .B2(new_n402), .ZN(new_n1029));
  XOR2_X1   g843(.A(new_n1029), .B(KEYINPUT122), .Z(new_n1030));
  NAND2_X1  g844(.A1(new_n881), .A2(new_n873), .ZN(new_n1031));
  INV_X1    g845(.A(new_n1031), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1030), .B1(new_n1032), .B2(G953), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n972), .B1(G898), .B2(new_n219), .ZN(new_n1034));
  XNOR2_X1  g848(.A(new_n1033), .B(new_n1034), .ZN(G69));
  NAND2_X1  g849(.A1(new_n338), .A2(new_n339), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n557), .B1(new_n558), .B2(new_n187), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1037), .B(KEYINPUT123), .Z(new_n1038));
  XNOR2_X1  g852(.A(new_n1036), .B(new_n1038), .ZN(new_n1039));
  INV_X1    g853(.A(new_n782), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n805), .A2(new_n813), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n909), .A2(new_n767), .ZN(new_n1042));
  XNOR2_X1  g856(.A(new_n1042), .B(KEYINPUT124), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n368), .A2(new_n924), .ZN(new_n1044));
  OAI21_X1  g858(.A(new_n784), .B1(new_n794), .B2(new_n1044), .ZN(new_n1045));
  OR4_X1    g859(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .A4(new_n1045), .ZN(new_n1046));
  AND2_X1   g860(.A1(new_n1046), .A2(new_n219), .ZN(new_n1047));
  NOR2_X1   g861(.A1(new_n219), .A2(G900), .ZN(new_n1048));
  XNOR2_X1  g862(.A(new_n1048), .B(KEYINPUT126), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1039), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  NOR3_X1   g864(.A1(new_n1043), .A2(new_n729), .A3(KEYINPUT62), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n646), .A2(new_n875), .ZN(new_n1052));
  NOR3_X1   g866(.A1(new_n897), .A2(new_n707), .A3(new_n770), .ZN(new_n1053));
  AOI211_X1 g867(.A(new_n1041), .B(new_n1051), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g868(.A(KEYINPUT62), .B1(new_n1043), .B2(new_n729), .ZN(new_n1055));
  XNOR2_X1  g869(.A(new_n1055), .B(KEYINPUT125), .ZN(new_n1056));
  AND2_X1   g870(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g871(.A1(new_n1057), .A2(G953), .ZN(new_n1058));
  OAI21_X1  g872(.A(new_n1050), .B1(new_n1058), .B2(new_n1039), .ZN(new_n1059));
  AOI21_X1  g873(.A(new_n219), .B1(G227), .B2(G900), .ZN(new_n1060));
  XNOR2_X1  g874(.A(new_n1059), .B(new_n1060), .ZN(G72));
  NAND2_X1  g875(.A1(new_n1057), .A2(new_n1032), .ZN(new_n1062));
  XNOR2_X1  g876(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1063));
  NOR2_X1   g877(.A1(new_n678), .A2(new_n443), .ZN(new_n1064));
  XNOR2_X1  g878(.A(new_n1063), .B(new_n1064), .ZN(new_n1065));
  AOI21_X1  g879(.A(new_n719), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g880(.A(new_n1065), .B1(new_n1046), .B2(new_n1031), .ZN(new_n1067));
  NAND4_X1  g881(.A1(new_n1067), .A2(new_n341), .A3(new_n313), .A4(new_n305), .ZN(new_n1068));
  OAI221_X1 g882(.A(new_n1065), .B1(new_n343), .B2(new_n357), .C1(new_n944), .C2(new_n945), .ZN(new_n1069));
  NAND3_X1  g883(.A1(new_n1068), .A2(new_n967), .A3(new_n1069), .ZN(new_n1070));
  NOR2_X1   g884(.A1(new_n1066), .A2(new_n1070), .ZN(G57));
endmodule


