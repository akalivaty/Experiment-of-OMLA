//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 0 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968;
  INV_X1    g000(.A(G127gat), .ZN(new_n202));
  INV_X1    g001(.A(G134gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G127gat), .A2(G134gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT72), .ZN(new_n207));
  AOI21_X1  g006(.A(KEYINPUT1), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT71), .ZN(new_n209));
  INV_X1    g008(.A(G113gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n209), .B1(new_n210), .B2(G120gat), .ZN(new_n211));
  INV_X1    g010(.A(G120gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n212), .A2(KEYINPUT71), .A3(G113gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n211), .B(new_n213), .C1(G113gat), .C2(new_n212), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n204), .A2(KEYINPUT72), .A3(new_n205), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n208), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G113gat), .B(G120gat), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n204), .B(new_n205), .C1(new_n217), .C2(KEYINPUT1), .ZN(new_n218));
  AND2_X1   g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT2), .ZN(new_n220));
  AOI22_X1  g019(.A1(new_n220), .A2(KEYINPUT82), .B1(G155gat), .B2(G162gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(G141gat), .B(G148gat), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n220), .B1(G155gat), .B2(G162gat), .ZN(new_n223));
  OAI221_X1 g022(.A(new_n221), .B1(G155gat), .B2(G162gat), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n222), .A2(new_n223), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n221), .B1(G155gat), .B2(G162gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n219), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n230), .B(KEYINPUT4), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n216), .A2(new_n218), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n224), .A2(new_n227), .A3(new_n233), .ZN(new_n234));
  NOR3_X1   g033(.A1(new_n229), .A2(KEYINPUT83), .A3(new_n233), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT83), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n236), .B1(new_n228), .B2(KEYINPUT3), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n232), .B(new_n234), .C1(new_n235), .C2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n231), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G225gat), .A2(G233gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT5), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n232), .A2(new_n228), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n240), .B1(new_n230), .B2(new_n243), .ZN(new_n244));
  OAI22_X1  g043(.A1(new_n239), .A2(new_n241), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n231), .A2(new_n238), .A3(KEYINPUT5), .A4(new_n240), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G1gat), .B(G29gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT0), .ZN(new_n249));
  XNOR2_X1  g048(.A(G57gat), .B(G85gat), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n249), .B(new_n250), .Z(new_n251));
  NAND2_X1  g050(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT6), .ZN(new_n253));
  INV_X1    g052(.A(new_n251), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n245), .A2(new_n254), .A3(new_n246), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n252), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  OR2_X1    g055(.A1(new_n255), .A2(new_n253), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G8gat), .B(G36gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(G64gat), .B(G92gat), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n259), .B(new_n260), .Z(new_n261));
  NAND2_X1  g060(.A1(G226gat), .A2(G233gat), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G183gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(KEYINPUT24), .ZN(new_n265));
  NAND2_X1  g064(.A1(G183gat), .A2(G190gat), .ZN(new_n266));
  AOI22_X1  g065(.A1(new_n265), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n268));
  INV_X1    g067(.A(G190gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(new_n264), .A3(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT23), .ZN(new_n275));
  INV_X1    g074(.A(G169gat), .ZN(new_n276));
  INV_X1    g075(.A(G176gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(G169gat), .A2(G176gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT23), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n279), .A2(KEYINPUT25), .A3(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT67), .B1(new_n273), .B2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n281), .A2(KEYINPUT65), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT65), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n280), .A2(new_n286), .A3(KEYINPUT23), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n285), .A2(new_n287), .A3(new_n279), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n266), .A2(KEYINPUT24), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT24), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(G183gat), .A3(G190gat), .ZN(new_n291));
  AOI22_X1  g090(.A1(new_n289), .A2(new_n291), .B1(new_n264), .B2(new_n269), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n284), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n289), .A2(new_n291), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n294), .A2(new_n271), .A3(new_n270), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT67), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n281), .A2(KEYINPUT25), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n295), .A2(new_n296), .A3(new_n279), .A4(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n283), .A2(new_n293), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n274), .ZN(new_n303));
  OAI22_X1  g102(.A1(new_n303), .A2(KEYINPUT70), .B1(new_n278), .B2(KEYINPUT26), .ZN(new_n304));
  OR2_X1    g103(.A1(new_n278), .A2(KEYINPUT26), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n302), .B(new_n304), .C1(KEYINPUT70), .C2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n307));
  XOR2_X1   g106(.A(KEYINPUT27), .B(G183gat), .Z(new_n308));
  OAI21_X1  g107(.A(new_n307), .B1(new_n308), .B2(G190gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT68), .ZN(new_n310));
  OR2_X1    g109(.A1(new_n310), .A2(KEYINPUT28), .ZN(new_n311));
  OR3_X1    g110(.A1(new_n308), .A2(G190gat), .A3(new_n311), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n306), .A2(new_n309), .A3(new_n312), .A4(new_n266), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n299), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n263), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n316), .B1(new_n263), .B2(new_n314), .ZN(new_n317));
  XOR2_X1   g116(.A(G211gat), .B(G218gat), .Z(new_n318));
  AND2_X1   g117(.A1(new_n318), .A2(KEYINPUT79), .ZN(new_n319));
  XOR2_X1   g118(.A(KEYINPUT78), .B(G218gat), .Z(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT77), .B(G211gat), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT22), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  XOR2_X1   g121(.A(G197gat), .B(G204gat), .Z(new_n323));
  OAI21_X1  g122(.A(new_n319), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n318), .A2(KEYINPUT79), .ZN(new_n325));
  INV_X1    g124(.A(new_n323), .ZN(new_n326));
  XOR2_X1   g125(.A(KEYINPUT77), .B(G211gat), .Z(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT78), .B(G218gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n325), .B(new_n326), .C1(new_n329), .C2(KEYINPUT22), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n324), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n317), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n314), .A2(new_n263), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT80), .B(KEYINPUT29), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n334), .B1(new_n299), .B2(new_n313), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n333), .B1(new_n263), .B2(new_n335), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n324), .A2(new_n330), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n261), .B1(new_n332), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n332), .A2(new_n338), .A3(new_n261), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n339), .B1(new_n341), .B2(KEYINPUT30), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT30), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n340), .A2(KEYINPUT81), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT81), .B1(new_n340), .B2(new_n343), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n258), .B(new_n342), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G228gat), .A2(G233gat), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT29), .B1(new_n324), .B2(new_n330), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n228), .B1(new_n350), .B2(KEYINPUT3), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT85), .ZN(new_n352));
  INV_X1    g151(.A(new_n334), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n234), .A2(new_n353), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n337), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n352), .B1(new_n337), .B2(new_n354), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n349), .B(new_n351), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n348), .B(KEYINPUT84), .Z(new_n358));
  INV_X1    g157(.A(new_n318), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n359), .B1(new_n322), .B2(new_n323), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n318), .B(new_n326), .C1(new_n329), .C2(KEYINPUT22), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(new_n361), .A3(new_n353), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n229), .B1(new_n362), .B2(new_n233), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n331), .B1(new_n234), .B2(new_n353), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n358), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n357), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT86), .B1(new_n366), .B2(G22gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(G78gat), .B(G106gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT31), .B(G50gat), .ZN(new_n369));
  XOR2_X1   g168(.A(new_n368), .B(new_n369), .Z(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G22gat), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n372), .B1(new_n357), .B2(new_n365), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n357), .A2(new_n372), .A3(new_n365), .ZN(new_n374));
  OAI22_X1  g173(.A1(new_n367), .A2(new_n371), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n373), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n357), .A2(new_n372), .A3(new_n365), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n376), .A2(KEYINPUT86), .A3(new_n377), .A4(new_n370), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(KEYINPUT75), .B(KEYINPUT34), .Z(new_n381));
  NAND3_X1  g180(.A1(new_n299), .A2(new_n313), .A3(new_n219), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT73), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n299), .A2(new_n313), .A3(KEYINPUT73), .A4(new_n219), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT74), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n387), .B1(new_n314), .B2(new_n232), .ZN(new_n388));
  AOI211_X1 g187(.A(KEYINPUT74), .B(new_n219), .C1(new_n299), .C2(new_n313), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n386), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(G227gat), .A2(G233gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n381), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n314), .A2(new_n232), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT74), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n314), .A2(new_n387), .A3(new_n232), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n395), .A2(new_n396), .B1(new_n384), .B2(new_n385), .ZN(new_n397));
  INV_X1    g196(.A(new_n381), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(new_n391), .A3(new_n398), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n393), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(KEYINPUT32), .B1(new_n397), .B2(new_n391), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT33), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n402), .B1(new_n397), .B2(new_n391), .ZN(new_n403));
  XOR2_X1   g202(.A(G15gat), .B(G43gat), .Z(new_n404));
  XNOR2_X1  g203(.A(G71gat), .B(G99gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n404), .B(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n401), .A2(new_n403), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n406), .ZN(new_n408));
  OAI221_X1 g207(.A(KEYINPUT32), .B1(new_n402), .B2(new_n408), .C1(new_n397), .C2(new_n391), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n400), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n407), .A2(new_n409), .B1(new_n393), .B2(new_n399), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n380), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT91), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n407), .A2(new_n409), .ZN(new_n415));
  INV_X1    g214(.A(new_n400), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n400), .A2(new_n407), .A3(new_n409), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n419), .A2(KEYINPUT91), .A3(new_n380), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n347), .B1(new_n414), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT92), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT35), .ZN(new_n423));
  NOR3_X1   g222(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n258), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n342), .B1(new_n345), .B2(new_n346), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT91), .B1(new_n419), .B2(new_n380), .ZN(new_n428));
  AOI211_X1 g227(.A(new_n413), .B(new_n379), .C1(new_n417), .C2(new_n418), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT92), .B1(new_n430), .B2(KEYINPUT35), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n256), .A2(KEYINPUT88), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT88), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n252), .A2(new_n433), .A3(new_n253), .A4(new_n255), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n255), .A2(new_n253), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(KEYINPUT90), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n426), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(new_n423), .A3(new_n439), .ZN(new_n440));
  OAI22_X1  g239(.A1(new_n424), .A2(new_n431), .B1(new_n412), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n317), .A2(new_n337), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT37), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n443), .B1(new_n336), .B2(new_n331), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT38), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n261), .A2(new_n443), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n445), .B1(new_n339), .B2(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(KEYINPUT89), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n332), .A2(new_n338), .ZN(new_n449));
  OAI22_X1  g248(.A1(new_n449), .A2(new_n443), .B1(new_n339), .B2(new_n446), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n341), .B1(new_n450), .B2(KEYINPUT38), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n435), .A2(new_n437), .A3(new_n448), .A4(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT40), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n239), .A2(new_n241), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n230), .A2(new_n240), .A3(new_n243), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n454), .A2(KEYINPUT39), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n251), .B1(new_n454), .B2(KEYINPUT39), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n453), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n255), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n456), .A2(new_n457), .A3(new_n453), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT87), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n461), .A2(new_n426), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n462), .B1(new_n461), .B2(new_n426), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n452), .B(new_n380), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n347), .A2(new_n379), .ZN(new_n466));
  INV_X1    g265(.A(new_n419), .ZN(new_n467));
  XOR2_X1   g266(.A(KEYINPUT76), .B(KEYINPUT36), .Z(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT76), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n419), .B1(new_n470), .B2(KEYINPUT36), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n465), .A2(new_n466), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n441), .A2(KEYINPUT93), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT93), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n440), .A2(new_n412), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n422), .B1(new_n421), .B2(new_n423), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n430), .A2(KEYINPUT92), .A3(KEYINPUT35), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n473), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n475), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT98), .ZN(new_n482));
  XNOR2_X1  g281(.A(G43gat), .B(G50gat), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NOR3_X1   g284(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n486));
  OAI22_X1  g285(.A1(new_n483), .A2(KEYINPUT15), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(G50gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(G43gat), .ZN(new_n489));
  INV_X1    g288(.A(G43gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(G50gat), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n489), .A2(new_n491), .A3(KEYINPUT15), .ZN(new_n492));
  NAND2_X1  g291(.A1(G29gat), .A2(G36gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n487), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT94), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n484), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(KEYINPUT94), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n499));
  INV_X1    g298(.A(G36gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n497), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n492), .B1(new_n502), .B2(new_n493), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT17), .B1(new_n495), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n491), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT15), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n501), .A2(new_n484), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n507), .A2(new_n492), .A3(new_n493), .A4(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT17), .ZN(new_n510));
  AOI22_X1  g309(.A1(new_n484), .A2(new_n496), .B1(new_n499), .B2(new_n500), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n511), .A2(new_n498), .B1(G29gat), .B2(G36gat), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n509), .B(new_n510), .C1(new_n512), .C2(new_n492), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n504), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT96), .ZN(new_n515));
  XOR2_X1   g314(.A(KEYINPUT95), .B(G8gat), .Z(new_n516));
  INV_X1    g315(.A(G15gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(G22gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n372), .A2(G15gat), .ZN(new_n519));
  INV_X1    g318(.A(G1gat), .ZN(new_n520));
  AND4_X1   g319(.A1(KEYINPUT16), .A2(new_n518), .A3(new_n519), .A4(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n520), .B1(new_n518), .B2(new_n519), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n515), .B(new_n516), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n518), .A2(new_n519), .A3(KEYINPUT16), .A4(new_n520), .ZN(new_n524));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n524), .B(G8gat), .C1(new_n520), .C2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n524), .B1(new_n520), .B2(new_n525), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n515), .B1(new_n528), .B2(new_n516), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n530), .ZN(new_n531));
  OAI22_X1  g330(.A1(new_n527), .A2(new_n529), .B1(new_n503), .B2(new_n495), .ZN(new_n532));
  NAND2_X1  g331(.A1(G229gat), .A2(G233gat), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT18), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n534), .A2(KEYINPUT97), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT97), .B1(new_n534), .B2(new_n535), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n531), .A2(KEYINPUT18), .A3(new_n532), .A4(new_n533), .ZN(new_n538));
  INV_X1    g337(.A(new_n529), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n495), .A2(new_n503), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n539), .A2(new_n540), .A3(new_n526), .A4(new_n523), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(new_n532), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n533), .B(KEYINPUT13), .Z(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  NOR3_X1   g344(.A1(new_n536), .A2(new_n537), .A3(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G113gat), .B(G141gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(G197gat), .ZN(new_n548));
  XOR2_X1   g347(.A(KEYINPUT11), .B(G169gat), .Z(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT12), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n482), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n551), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n534), .A2(new_n535), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT97), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n545), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g357(.A(KEYINPUT98), .B(new_n553), .C1(new_n558), .C2(new_n536), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n552), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n557), .A2(new_n551), .A3(new_n554), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n474), .A2(new_n481), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G71gat), .B(G78gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(G57gat), .B(G64gat), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n564), .B1(new_n566), .B2(KEYINPUT9), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n565), .A2(KEYINPUT99), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(KEYINPUT99), .ZN(new_n569));
  AND3_X1   g368(.A1(new_n568), .A2(new_n564), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n571), .B(KEYINPUT100), .Z(new_n572));
  AOI21_X1  g371(.A(new_n567), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n573), .A2(KEYINPUT21), .ZN(new_n574));
  XNOR2_X1  g373(.A(G127gat), .B(G155gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  AOI211_X1 g375(.A(new_n529), .B(new_n527), .C1(new_n573), .C2(KEYINPUT21), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT101), .ZN(new_n580));
  XOR2_X1   g379(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G183gat), .B(G211gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n578), .B(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G85gat), .A2(G92gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n587), .B(new_n588), .Z(new_n589));
  INV_X1    g388(.A(KEYINPUT103), .ZN(new_n590));
  INV_X1    g389(.A(G92gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(G85gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(KEYINPUT103), .A2(G92gat), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT104), .ZN(new_n596));
  INV_X1    g395(.A(G99gat), .ZN(new_n597));
  INV_X1    g396(.A(G106gat), .ZN(new_n598));
  OAI21_X1  g397(.A(KEYINPUT8), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n595), .A2(new_n596), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n596), .B1(new_n595), .B2(new_n599), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n589), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G99gat), .B(G106gat), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n603), .B(new_n589), .C1(new_n600), .C2(new_n601), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n605), .A2(KEYINPUT105), .A3(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT105), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n602), .A2(new_n608), .A3(new_n604), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n607), .A2(new_n514), .A3(new_n609), .ZN(new_n610));
  AND2_X1   g409(.A1(G232gat), .A2(G233gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT41), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n540), .B1(new_n607), .B2(new_n609), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(G190gat), .B(G218gat), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n615), .B(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(G134gat), .B(G162gat), .Z(new_n619));
  NOR2_X1   g418(.A1(new_n611), .A2(KEYINPUT41), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n618), .A2(new_n621), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G120gat), .B(G148gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(G176gat), .B(G204gat), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n626), .B(new_n627), .Z(new_n628));
  NAND3_X1  g427(.A1(new_n573), .A2(new_n605), .A3(new_n606), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n570), .A2(new_n572), .ZN(new_n631));
  INV_X1    g430(.A(new_n567), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n607), .A2(new_n633), .A3(new_n609), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT106), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT106), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n607), .A2(new_n636), .A3(new_n633), .A4(new_n609), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n630), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G230gat), .A2(G233gat), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n628), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n635), .A2(new_n637), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT10), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n641), .A2(new_n642), .A3(new_n629), .ZN(new_n643));
  AOI211_X1 g442(.A(new_n642), .B(new_n633), .C1(new_n607), .C2(new_n609), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n640), .B1(new_n646), .B2(new_n639), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n638), .A2(new_n639), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n644), .B1(new_n638), .B2(new_n642), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n639), .B(KEYINPUT107), .Z(new_n650));
  OAI21_X1  g449(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n628), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n647), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n586), .A2(new_n625), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT108), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n563), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n656), .A2(new_n258), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(new_n520), .ZN(G1324gat));
  NAND3_X1  g457(.A1(new_n563), .A2(new_n426), .A3(new_n655), .ZN(new_n659));
  AND2_X1   g458(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n660));
  NOR2_X1   g459(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n659), .A2(G8gat), .ZN(new_n663));
  OAI21_X1  g462(.A(KEYINPUT42), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n664), .B1(KEYINPUT42), .B2(new_n662), .ZN(G1325gat));
  OAI21_X1  g464(.A(G15gat), .B1(new_n656), .B2(new_n472), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n419), .A2(new_n517), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n666), .B1(new_n656), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT109), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n666), .B(KEYINPUT109), .C1(new_n656), .C2(new_n667), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(G1326gat));
  OAI21_X1  g471(.A(KEYINPUT110), .B1(new_n656), .B2(new_n380), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT110), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n563), .A2(new_n674), .A3(new_n379), .A4(new_n655), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT43), .B(G22gat), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n673), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n676), .B1(new_n673), .B2(new_n675), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(G1327gat));
  NAND2_X1  g478(.A1(new_n653), .A2(new_n585), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(new_n625), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n563), .A2(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n258), .A2(G29gat), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT45), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n625), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n474), .A2(new_n481), .A3(new_n688), .ZN(new_n689));
  AOI211_X1 g488(.A(KEYINPUT111), .B(new_n380), .C1(new_n439), .C2(new_n258), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT111), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n691), .B1(new_n347), .B2(new_n379), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n693), .A2(new_n465), .A3(new_n472), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n479), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n687), .B1(new_n695), .B2(new_n625), .ZN(new_n696));
  INV_X1    g495(.A(new_n562), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n680), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n689), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT112), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT112), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n689), .A2(new_n696), .A3(new_n701), .A4(new_n698), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n700), .A2(new_n425), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(G29gat), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n686), .A2(new_n704), .ZN(G1328gat));
  NOR3_X1   g504(.A1(new_n682), .A2(G36gat), .A3(new_n439), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT113), .B(KEYINPUT46), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n700), .A2(new_n426), .A3(new_n702), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(G36gat), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n706), .A2(new_n708), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n709), .A2(new_n711), .A3(new_n712), .ZN(G1329gat));
  OAI21_X1  g512(.A(G43gat), .B1(new_n699), .B2(new_n472), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n419), .A2(new_n490), .ZN(new_n715));
  OAI211_X1 g514(.A(new_n714), .B(KEYINPUT47), .C1(new_n682), .C2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n682), .A2(new_n715), .ZN(new_n717));
  INV_X1    g516(.A(new_n472), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n700), .A2(new_n718), .A3(new_n702), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n717), .B1(new_n719), .B2(G43gat), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n716), .B1(new_n720), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g520(.A(G50gat), .B1(new_n699), .B2(new_n380), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n379), .A2(new_n488), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n722), .B(KEYINPUT48), .C1(new_n682), .C2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n682), .A2(new_n723), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n700), .A2(new_n379), .A3(new_n702), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n725), .B1(new_n726), .B2(G50gat), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n724), .B1(new_n727), .B2(KEYINPUT48), .ZN(G1331gat));
  OR2_X1    g527(.A1(new_n479), .A2(new_n694), .ZN(new_n729));
  NOR4_X1   g528(.A1(new_n562), .A2(new_n624), .A3(new_n653), .A4(new_n585), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n425), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(G57gat), .ZN(G1332gat));
  INV_X1    g532(.A(KEYINPUT49), .ZN(new_n734));
  INV_X1    g533(.A(G64gat), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n731), .B(new_n426), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n735), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1333gat));
  XNOR2_X1  g537(.A(new_n419), .B(KEYINPUT115), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n731), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n729), .A2(G71gat), .A3(new_n718), .A4(new_n730), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n742), .A2(KEYINPUT114), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(KEYINPUT114), .ZN(new_n744));
  OAI22_X1  g543(.A1(new_n741), .A2(G71gat), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n379), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g547(.A1(new_n586), .A2(new_n562), .A3(new_n653), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n689), .A2(new_n696), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G85gat), .B1(new_n750), .B2(new_n258), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n586), .A2(new_n562), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n624), .B(new_n752), .C1(new_n479), .C2(new_n694), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n653), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n425), .A2(new_n593), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n751), .B1(new_n757), .B2(new_n758), .ZN(G1336gat));
  NAND2_X1  g558(.A1(new_n592), .A2(new_n594), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n750), .B2(new_n439), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n426), .A2(new_n591), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n761), .B(new_n762), .C1(new_n757), .C2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT116), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n753), .A2(new_n765), .A3(new_n754), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n763), .A2(new_n653), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n766), .B(new_n767), .C1(new_n755), .C2(new_n765), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n768), .A2(new_n761), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n764), .B1(new_n769), .B2(new_n762), .ZN(G1337gat));
  NOR3_X1   g569(.A1(new_n750), .A2(new_n597), .A3(new_n472), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n755), .A2(new_n419), .A3(new_n756), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n771), .B1(new_n597), .B2(new_n772), .ZN(G1338gat));
  NOR3_X1   g572(.A1(new_n653), .A2(new_n380), .A3(G106gat), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n766), .B(new_n774), .C1(new_n755), .C2(new_n765), .ZN(new_n775));
  OAI21_X1  g574(.A(G106gat), .B1(new_n750), .B2(new_n380), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT53), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT53), .B1(new_n755), .B2(new_n774), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n776), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(G1339gat));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n782), .B1(new_n646), .B2(new_n639), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT117), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n649), .A2(new_n784), .A3(new_n650), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n643), .A2(new_n650), .A3(new_n645), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT117), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n783), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n650), .ZN(new_n789));
  AOI211_X1 g588(.A(KEYINPUT10), .B(new_n630), .C1(new_n635), .C2(new_n637), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n782), .B(new_n789), .C1(new_n790), .C2(new_n644), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n791), .A2(KEYINPUT55), .A3(new_n652), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n647), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n531), .A2(new_n532), .ZN(new_n795));
  OAI22_X1  g594(.A1(new_n795), .A2(new_n533), .B1(new_n542), .B2(new_n543), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n550), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n561), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n793), .A2(new_n624), .A3(new_n794), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n791), .A2(new_n652), .ZN(new_n800));
  INV_X1    g599(.A(new_n639), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT54), .B1(new_n649), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n784), .B1(new_n649), .B2(new_n650), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n800), .B1(new_n804), .B2(new_n785), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT118), .B1(new_n805), .B2(KEYINPUT55), .ZN(new_n806));
  INV_X1    g605(.A(new_n800), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT55), .B1(new_n788), .B2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n799), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n647), .B1(new_n560), .B2(new_n561), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n793), .A2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n805), .A2(KEYINPUT118), .A3(KEYINPUT55), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n808), .A2(new_n809), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n756), .A2(new_n798), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n811), .B1(new_n819), .B2(new_n625), .ZN(new_n820));
  OAI22_X1  g619(.A1(new_n820), .A2(new_n586), .B1(new_n562), .B2(new_n654), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n821), .A2(new_n380), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n426), .A2(new_n258), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(new_n419), .A3(new_n823), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n824), .A2(new_n210), .A3(new_n697), .ZN(new_n825));
  INV_X1    g624(.A(new_n821), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n428), .A2(new_n429), .ZN(new_n827));
  NOR4_X1   g626(.A1(new_n826), .A2(new_n258), .A3(new_n426), .A4(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(G113gat), .B1(new_n828), .B2(new_n562), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n825), .A2(new_n829), .ZN(G1340gat));
  NOR3_X1   g629(.A1(new_n824), .A2(new_n212), .A3(new_n653), .ZN(new_n831));
  AOI21_X1  g630(.A(G120gat), .B1(new_n828), .B2(new_n756), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n831), .A2(new_n832), .ZN(G1341gat));
  OAI21_X1  g632(.A(G127gat), .B1(new_n824), .B2(new_n585), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n828), .A2(new_n202), .A3(new_n586), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(G1342gat));
  NAND3_X1  g635(.A1(new_n828), .A2(new_n203), .A3(new_n624), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n837), .A2(KEYINPUT56), .ZN(new_n838));
  OAI21_X1  g637(.A(G134gat), .B1(new_n824), .B2(new_n625), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(KEYINPUT56), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(G1343gat));
  NOR2_X1   g640(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(KEYINPUT122), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(G141gat), .ZN(new_n845));
  INV_X1    g644(.A(new_n823), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n718), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n654), .A2(new_n562), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n818), .B1(new_n813), .B2(new_n808), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n625), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n811), .B1(new_n851), .B2(KEYINPUT119), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n793), .B(new_n812), .C1(new_n805), .C2(KEYINPUT55), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n624), .B1(new_n853), .B2(new_n818), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n586), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n849), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n815), .A2(new_n816), .ZN(new_n860));
  OAI22_X1  g659(.A1(new_n854), .A2(new_n855), .B1(new_n860), .B2(new_n799), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n851), .A2(KEYINPUT119), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n585), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(KEYINPUT120), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n380), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT57), .B1(new_n821), .B2(new_n379), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n848), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n845), .B1(new_n871), .B2(new_n562), .ZN(new_n872));
  NAND2_X1  g671(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n826), .A2(new_n258), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n718), .A2(new_n426), .A3(new_n380), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n697), .A2(G141gat), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n873), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n844), .B1(new_n872), .B2(new_n879), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n874), .A2(new_n875), .ZN(new_n881));
  AOI22_X1  g680(.A1(new_n881), .A2(new_n877), .B1(KEYINPUT121), .B2(KEYINPUT58), .ZN(new_n882));
  AOI211_X1 g681(.A(new_n697), .B(new_n848), .C1(new_n868), .C2(new_n870), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n882), .B(new_n843), .C1(new_n883), .C2(new_n845), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n880), .A2(new_n884), .ZN(G1344gat));
  AND2_X1   g684(.A1(new_n821), .A2(new_n867), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n655), .A2(new_n697), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n585), .B1(new_n854), .B2(new_n811), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT57), .B1(new_n889), .B2(new_n379), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n847), .A2(new_n756), .ZN(new_n892));
  OAI21_X1  g691(.A(G148gat), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT59), .ZN(new_n894));
  INV_X1    g693(.A(new_n867), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n895), .B1(new_n859), .B2(new_n864), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n756), .B(new_n847), .C1(new_n896), .C2(new_n869), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT123), .ZN(new_n898));
  INV_X1    g697(.A(G148gat), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(KEYINPUT59), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n897), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n898), .B1(new_n897), .B2(new_n900), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n894), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n881), .A2(new_n899), .A3(new_n756), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1345gat));
  NOR3_X1   g704(.A1(new_n876), .A2(KEYINPUT124), .A3(new_n585), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n906), .A2(G155gat), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT124), .B1(new_n876), .B2(new_n585), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n586), .A2(G155gat), .ZN(new_n909));
  AOI22_X1  g708(.A1(new_n907), .A2(new_n908), .B1(new_n871), .B2(new_n909), .ZN(G1346gat));
  INV_X1    g709(.A(G162gat), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n624), .B(new_n847), .C1(new_n896), .C2(new_n869), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n911), .B1(new_n912), .B2(KEYINPUT125), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n913), .B1(KEYINPUT125), .B2(new_n912), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n881), .A2(new_n911), .A3(new_n624), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1347gat));
  AND2_X1   g715(.A1(new_n821), .A2(new_n258), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n827), .A2(new_n439), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(new_n276), .A3(new_n562), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT126), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n439), .A2(new_n425), .ZN(new_n923));
  AND4_X1   g722(.A1(new_n380), .A2(new_n821), .A3(new_n739), .A4(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n562), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n922), .B1(new_n925), .B2(G169gat), .ZN(new_n926));
  AOI211_X1 g725(.A(KEYINPUT126), .B(new_n276), .C1(new_n924), .C2(new_n562), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n921), .B1(new_n926), .B2(new_n927), .ZN(G1348gat));
  NAND3_X1  g727(.A1(new_n920), .A2(new_n277), .A3(new_n756), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n924), .A2(new_n756), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n929), .B1(new_n277), .B2(new_n930), .ZN(G1349gat));
  NOR3_X1   g730(.A1(new_n919), .A2(new_n308), .A3(new_n585), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n264), .B1(new_n924), .B2(new_n586), .ZN(new_n933));
  OR3_X1    g732(.A1(new_n932), .A2(KEYINPUT60), .A3(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(KEYINPUT60), .B1(new_n932), .B2(new_n933), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1350gat));
  NAND3_X1  g735(.A1(new_n920), .A2(new_n269), .A3(new_n624), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT61), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n924), .A2(new_n624), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n939), .B2(G190gat), .ZN(new_n940));
  AOI211_X1 g739(.A(KEYINPUT61), .B(new_n269), .C1(new_n924), .C2(new_n624), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(G1351gat));
  OR2_X1    g741(.A1(new_n886), .A2(new_n890), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n472), .A2(new_n923), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(G197gat), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n945), .A2(new_n946), .A3(new_n697), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n718), .A2(new_n439), .A3(new_n380), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n917), .A2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(G197gat), .B1(new_n950), .B2(new_n562), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n947), .A2(new_n951), .ZN(G1352gat));
  NOR3_X1   g751(.A1(new_n949), .A2(G204gat), .A3(new_n653), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT62), .ZN(new_n954));
  OAI21_X1  g753(.A(G204gat), .B1(new_n945), .B2(new_n653), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1353gat));
  NAND3_X1  g755(.A1(new_n950), .A2(new_n327), .A3(new_n586), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n943), .A2(new_n586), .A3(new_n944), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n958), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT63), .B1(new_n958), .B2(G211gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(G1354gat));
  INV_X1    g760(.A(G218gat), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n962), .B1(new_n949), .B2(new_n625), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n624), .A2(new_n320), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n963), .B1(new_n945), .B2(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT127), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI211_X1 g766(.A(KEYINPUT127), .B(new_n963), .C1(new_n945), .C2(new_n964), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(G1355gat));
endmodule


