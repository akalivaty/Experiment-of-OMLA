//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G469), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(new_n193), .A3(G128), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT67), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  AND2_X1   g010(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n197));
  NOR2_X1   g011(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(G143), .B(G146), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT67), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n199), .A2(new_n200), .A3(new_n201), .A4(G128), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n196), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n200), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  INV_X1    g019(.A(new_n193), .ZN(new_n206));
  AOI22_X1  g020(.A1(new_n204), .A2(new_n205), .B1(KEYINPUT1), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G101), .ZN(new_n209));
  INV_X1    g023(.A(G104), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G107), .ZN(new_n211));
  INV_X1    g025(.A(G107), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G104), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n209), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT3), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT78), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(KEYINPUT78), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n217), .B1(new_n218), .B2(new_n213), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n216), .A2(new_n212), .A3(KEYINPUT78), .A4(G104), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n219), .A2(new_n209), .A3(new_n211), .A4(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n208), .A2(new_n215), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT10), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G134), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT11), .B1(new_n225), .B2(G137), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT11), .ZN(new_n227));
  INV_X1    g041(.A(G137), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n228), .A3(G134), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n226), .A2(new_n229), .B1(new_n225), .B2(G137), .ZN(new_n230));
  XOR2_X1   g044(.A(KEYINPUT64), .B(G131), .Z(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G131), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n232), .B1(new_n233), .B2(new_n230), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT79), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT78), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(KEYINPUT3), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n210), .A2(G107), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(KEYINPUT3), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n220), .A2(new_n211), .ZN(new_n242));
  NOR3_X1   g056(.A1(new_n241), .A2(new_n242), .A3(G101), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n236), .B1(new_n243), .B2(new_n214), .ZN(new_n244));
  INV_X1    g058(.A(new_n191), .ZN(new_n245));
  OAI21_X1  g059(.A(G128), .B1(new_n199), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n204), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n203), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n221), .A2(KEYINPUT79), .A3(new_n215), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n244), .A2(KEYINPUT10), .A3(new_n248), .A4(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(G101), .B1(new_n241), .B2(new_n242), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(KEYINPUT4), .A3(new_n221), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT0), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n200), .B1(new_n253), .B2(new_n205), .ZN(new_n254));
  XOR2_X1   g068(.A(KEYINPUT0), .B(G128), .Z(new_n255));
  OAI21_X1  g069(.A(new_n254), .B1(new_n200), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n257), .B(G101), .C1(new_n241), .C2(new_n242), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n252), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n224), .A2(new_n235), .A3(new_n250), .A4(new_n259), .ZN(new_n260));
  XOR2_X1   g074(.A(G110), .B(G140), .Z(new_n261));
  XNOR2_X1  g075(.A(new_n261), .B(KEYINPUT77), .ZN(new_n262));
  INV_X1    g076(.A(G953), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G227), .ZN(new_n264));
  XOR2_X1   g078(.A(new_n262), .B(new_n264), .Z(new_n265));
  NAND2_X1  g079(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT80), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n196), .A2(new_n202), .B1(new_n246), .B2(new_n204), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n221), .A2(KEYINPUT79), .A3(new_n215), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT79), .B1(new_n221), .B2(new_n215), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n267), .B(new_n268), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n222), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n244), .A2(new_n249), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n267), .B1(new_n273), .B2(new_n268), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n234), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT12), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI211_X1 g091(.A(KEYINPUT12), .B(new_n234), .C1(new_n272), .C2(new_n274), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n266), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n224), .A2(new_n250), .A3(new_n259), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n234), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n265), .B1(new_n281), .B2(new_n260), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n188), .B(new_n189), .C1(new_n279), .C2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n281), .A2(new_n265), .A3(new_n260), .ZN(new_n284));
  INV_X1    g098(.A(new_n260), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n285), .B1(new_n277), .B2(new_n278), .ZN(new_n286));
  OAI211_X1 g100(.A(G469), .B(new_n284), .C1(new_n286), .C2(new_n265), .ZN(new_n287));
  NAND2_X1  g101(.A1(G469), .A2(G902), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n283), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT9), .B(G234), .ZN(new_n290));
  OAI21_X1  g104(.A(G221), .B1(new_n290), .B2(G902), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n291), .B(KEYINPUT76), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(G210), .B1(G237), .B2(G902), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  AND2_X1   g110(.A1(KEYINPUT69), .A2(G116), .ZN(new_n297));
  NOR2_X1   g111(.A1(KEYINPUT69), .A2(G116), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G119), .ZN(new_n300));
  INV_X1    g114(.A(G116), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n301), .A2(G119), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n300), .A2(KEYINPUT5), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G113), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT5), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n305), .B1(new_n302), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G119), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n297), .A2(new_n298), .A3(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n309), .A2(new_n302), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT2), .B(G113), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n304), .A2(new_n307), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n244), .A2(new_n313), .A3(new_n249), .ZN(new_n314));
  XNOR2_X1  g128(.A(G110), .B(G122), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n300), .A2(new_n303), .A3(new_n312), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n311), .B1(new_n309), .B2(new_n302), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n252), .A2(new_n318), .A3(new_n258), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n314), .A2(new_n315), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G125), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n268), .A2(new_n322), .ZN(new_n323));
  OR2_X1    g137(.A1(new_n256), .A2(new_n322), .ZN(new_n324));
  INV_X1    g138(.A(G224), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n325), .A2(G953), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT7), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n323), .A2(new_n324), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n323), .A2(new_n324), .ZN(new_n330));
  INV_X1    g144(.A(new_n328), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n304), .A2(new_n307), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n316), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n221), .A2(new_n215), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n314), .A2(new_n336), .ZN(new_n337));
  XOR2_X1   g151(.A(new_n315), .B(KEYINPUT8), .Z(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n329), .A2(new_n332), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n321), .B1(new_n340), .B2(KEYINPUT84), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n332), .A2(new_n329), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n337), .A2(new_n339), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT84), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(G902), .B1(new_n341), .B2(new_n346), .ZN(new_n347));
  XOR2_X1   g161(.A(KEYINPUT82), .B(KEYINPUT6), .Z(new_n348));
  AOI211_X1 g162(.A(new_n315), .B(new_n348), .C1(new_n314), .C2(new_n319), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n330), .B(new_n327), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n320), .A2(KEYINPUT6), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n315), .B1(new_n314), .B2(new_n319), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n314), .A2(new_n319), .ZN(new_n355));
  INV_X1    g169(.A(new_n315), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n357), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(new_n320), .ZN(new_n358));
  AOI211_X1 g172(.A(new_n349), .B(new_n350), .C1(new_n354), .C2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT83), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n347), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n354), .A2(new_n358), .ZN(new_n362));
  INV_X1    g176(.A(new_n349), .ZN(new_n363));
  INV_X1    g177(.A(new_n350), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n362), .A2(new_n360), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n296), .B1(new_n361), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT83), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n369), .A2(new_n295), .A3(new_n365), .A4(new_n347), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT92), .ZN(new_n372));
  XNOR2_X1  g186(.A(KEYINPUT88), .B(G122), .ZN(new_n373));
  OR2_X1    g187(.A1(new_n373), .A2(new_n301), .ZN(new_n374));
  INV_X1    g188(.A(G122), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n297), .A2(new_n298), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n374), .A2(new_n212), .A3(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n373), .A2(new_n301), .ZN(new_n379));
  OAI21_X1  g193(.A(G107), .B1(new_n379), .B2(new_n376), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT89), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n382), .B1(new_n205), .B2(G143), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n192), .A2(KEYINPUT89), .A3(G128), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n385), .B1(G128), .B2(new_n192), .ZN(new_n386));
  OR2_X1    g200(.A1(new_n386), .A2(G134), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n381), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(KEYINPUT13), .B1(new_n383), .B2(new_n384), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT90), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n192), .A2(G128), .ZN(new_n392));
  OR3_X1    g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n391), .B1(new_n390), .B2(new_n392), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT91), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT13), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n395), .B1(new_n385), .B2(new_n396), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n383), .A2(new_n384), .A3(KEYINPUT91), .A4(KEYINPUT13), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n393), .A2(new_n394), .A3(new_n397), .A4(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G134), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n374), .B1(new_n377), .B2(KEYINPUT14), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n377), .A2(KEYINPUT14), .ZN(new_n402));
  OAI21_X1  g216(.A(G107), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n379), .A2(G107), .A3(new_n376), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n386), .A2(G134), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n404), .B1(new_n387), .B2(new_n405), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n389), .A2(new_n400), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G217), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n290), .A2(new_n408), .A3(G953), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n372), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n409), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n388), .B1(G134), .B2(new_n399), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n406), .A2(new_n403), .ZN(new_n413));
  OAI211_X1 g227(.A(KEYINPUT92), .B(new_n411), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n389), .A2(new_n400), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n406), .A2(new_n403), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n416), .A3(new_n409), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n410), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n189), .ZN(new_n419));
  INV_X1    g233(.A(G478), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n420), .A2(KEYINPUT15), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n419), .B(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(G113), .B(G122), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(G104), .ZN(new_n424));
  INV_X1    g238(.A(G237), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(new_n263), .A3(G214), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n192), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n425), .A2(new_n263), .A3(G143), .A4(G214), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(KEYINPUT18), .A3(G131), .ZN(new_n430));
  XNOR2_X1  g244(.A(G125), .B(G140), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(new_n190), .ZN(new_n432));
  NAND2_X1  g246(.A1(KEYINPUT18), .A2(G131), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n427), .A2(new_n428), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n430), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n231), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n429), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT85), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT17), .ZN(new_n441));
  AOI21_X1  g255(.A(KEYINPUT85), .B1(new_n429), .B2(new_n437), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n440), .B(new_n441), .C1(new_n438), .C2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n429), .A2(new_n437), .A3(KEYINPUT17), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n431), .A2(KEYINPUT16), .ZN(new_n446));
  OR3_X1    g260(.A1(new_n322), .A2(KEYINPUT16), .A3(G140), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(G146), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(G146), .B1(new_n446), .B2(new_n447), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n445), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  AOI211_X1 g265(.A(new_n424), .B(new_n436), .C1(new_n443), .C2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n424), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n443), .A2(new_n451), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n453), .B1(new_n454), .B2(new_n435), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n189), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(G475), .ZN(new_n457));
  NOR2_X1   g271(.A1(G475), .A2(G902), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n431), .A2(KEYINPUT86), .A3(KEYINPUT19), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n460), .B1(new_n431), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n190), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n442), .A2(new_n438), .ZN(new_n464));
  NOR3_X1   g278(.A1(new_n429), .A2(new_n437), .A3(KEYINPUT85), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n448), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n435), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n424), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n454), .A2(new_n453), .A3(new_n435), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n459), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT20), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(KEYINPUT87), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n453), .B1(new_n466), .B2(new_n435), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n458), .B1(new_n452), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT20), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT87), .B1(new_n470), .B2(new_n471), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n457), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(G234), .A2(G237), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n479), .A2(G952), .A3(new_n263), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n479), .A2(G902), .A3(G953), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT21), .B(G898), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR3_X1   g297(.A1(new_n422), .A2(new_n478), .A3(new_n483), .ZN(new_n484));
  AND4_X1   g298(.A1(new_n187), .A2(new_n294), .A3(new_n371), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n226), .A2(new_n229), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n225), .A2(G137), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n231), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT65), .B1(new_n228), .B2(G134), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT65), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(new_n225), .A3(G137), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n228), .A2(G134), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n233), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT71), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n488), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n490), .B1(new_n225), .B2(G137), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n228), .A2(KEYINPUT65), .A3(G134), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n493), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(G131), .ZN(new_n500));
  AOI21_X1  g314(.A(KEYINPUT71), .B1(new_n500), .B2(new_n232), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n248), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n318), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n230), .A2(new_n233), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n256), .B1(new_n488), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT70), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g321(.A(KEYINPUT70), .B(new_n256), .C1(new_n488), .C2(new_n504), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n502), .A2(new_n503), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT72), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n508), .ZN(new_n512));
  AOI21_X1  g326(.A(KEYINPUT70), .B1(new_n234), .B2(new_n256), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n514), .A2(KEYINPUT72), .A3(new_n503), .A4(new_n502), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n425), .A2(new_n263), .A3(G210), .ZN(new_n517));
  XOR2_X1   g331(.A(new_n517), .B(KEYINPUT27), .Z(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT26), .B(G101), .ZN(new_n519));
  XOR2_X1   g333(.A(new_n518), .B(new_n519), .Z(new_n520));
  NAND4_X1  g334(.A1(new_n248), .A2(KEYINPUT68), .A3(new_n232), .A4(new_n500), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT68), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n500), .A2(new_n232), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n522), .B1(new_n268), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n521), .A2(new_n524), .A3(new_n505), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT30), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n502), .A2(KEYINPUT30), .A3(new_n507), .A4(new_n508), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(new_n318), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n516), .A2(new_n520), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT31), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n516), .A2(new_n529), .A3(KEYINPUT31), .A4(new_n520), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT28), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI22_X1  g351(.A1(new_n511), .A2(new_n515), .B1(new_n318), .B2(new_n525), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n537), .B1(new_n538), .B2(new_n536), .ZN(new_n539));
  INV_X1    g353(.A(new_n520), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI211_X1 g355(.A(G472), .B(G902), .C1(new_n534), .C2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT73), .B1(new_n542), .B2(KEYINPUT32), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n534), .A2(new_n541), .ZN(new_n544));
  INV_X1    g358(.A(G472), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n545), .A3(new_n189), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT73), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT32), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n542), .A2(KEYINPUT32), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n520), .B(new_n537), .C1(new_n538), .C2(new_n536), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n520), .B1(new_n516), .B2(new_n529), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT29), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n503), .B1(new_n514), .B2(new_n502), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n555), .B1(new_n511), .B2(new_n515), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n537), .B1(new_n556), .B2(new_n536), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n520), .A2(KEYINPUT29), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n189), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(G472), .B1(new_n554), .B2(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n543), .A2(new_n549), .A3(new_n550), .A4(new_n560), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n205), .B(G119), .C1(KEYINPUT74), .C2(KEYINPUT23), .ZN(new_n562));
  AOI21_X1  g376(.A(KEYINPUT23), .B1(new_n205), .B2(G119), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n205), .A2(G119), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n562), .B1(new_n565), .B2(KEYINPUT74), .ZN(new_n566));
  XNOR2_X1  g380(.A(G119), .B(G128), .ZN(new_n567));
  XOR2_X1   g381(.A(KEYINPUT24), .B(G110), .Z(new_n568));
  OAI22_X1  g382(.A1(new_n566), .A2(G110), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n431), .A2(new_n190), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(new_n448), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n566), .A2(G110), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n568), .A2(new_n567), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n572), .B(new_n573), .C1(new_n449), .C2(new_n450), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT75), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT22), .B(G137), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n263), .A2(G221), .A3(G234), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT75), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n571), .A2(new_n574), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n576), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n571), .A2(new_n574), .A3(new_n579), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(KEYINPUT25), .B1(new_n586), .B2(G902), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT25), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n585), .A2(new_n588), .A3(new_n189), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n408), .B1(G234), .B2(new_n189), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n590), .A2(G902), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n585), .A2(new_n592), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n485), .A2(new_n561), .A3(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT93), .B(G101), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(G3));
  NAND2_X1  g411(.A1(new_n294), .A2(new_n594), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n544), .A2(new_n189), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(G472), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n546), .ZN(new_n601));
  OR3_X1    g415(.A1(new_n598), .A2(new_n601), .A3(KEYINPUT94), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT97), .ZN(new_n603));
  INV_X1    g417(.A(new_n478), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT96), .B(G478), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n605), .B1(new_n418), .B2(new_n189), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n607), .A2(KEYINPUT33), .A3(new_n417), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT33), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n608), .B1(new_n418), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n420), .A2(G902), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n606), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n603), .B1(new_n604), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n610), .A2(new_n611), .ZN(new_n614));
  INV_X1    g428(.A(new_n606), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n616), .A2(KEYINPUT97), .A3(new_n478), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n483), .B1(new_n613), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT95), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n370), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n320), .B1(new_n344), .B2(new_n345), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n340), .A2(KEYINPUT84), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n189), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(KEYINPUT83), .B2(new_n368), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n624), .A2(KEYINPUT95), .A3(new_n295), .A4(new_n365), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n620), .A2(new_n625), .A3(new_n367), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n618), .A2(new_n187), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(KEYINPUT94), .B1(new_n598), .B2(new_n601), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n602), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT34), .B(G104), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  NAND2_X1  g445(.A1(new_n626), .A2(new_n187), .ZN(new_n632));
  INV_X1    g446(.A(new_n483), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n470), .A2(new_n471), .ZN(new_n634));
  AOI22_X1  g448(.A1(new_n634), .A2(new_n475), .B1(G475), .B2(new_n456), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n422), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n602), .A2(new_n628), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT35), .B(G107), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  INV_X1    g454(.A(KEYINPUT99), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n576), .A2(new_n582), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT98), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT98), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n576), .A2(new_n644), .A3(new_n582), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n580), .A2(KEYINPUT36), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n643), .B(new_n645), .C1(KEYINPUT36), .C2(new_n580), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n641), .B1(new_n650), .B2(new_n592), .ZN(new_n651));
  INV_X1    g465(.A(new_n592), .ZN(new_n652));
  AOI211_X1 g466(.A(KEYINPUT99), .B(new_n652), .C1(new_n648), .C2(new_n649), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n591), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n485), .A2(new_n546), .A3(new_n600), .A4(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT37), .B(G110), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  INV_X1    g471(.A(new_n632), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n294), .A2(new_n654), .ZN(new_n659));
  INV_X1    g473(.A(G900), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n480), .B1(new_n481), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  AOI211_X1 g476(.A(KEYINPUT15), .B(new_n420), .C1(new_n418), .C2(new_n189), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n419), .A2(new_n421), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n635), .B(new_n662), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(KEYINPUT100), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT100), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n422), .A2(new_n667), .A3(new_n635), .A4(new_n662), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n659), .A2(new_n669), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n658), .A2(new_n670), .A3(new_n561), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(new_n205), .ZN(G30));
  XOR2_X1   g486(.A(KEYINPUT101), .B(KEYINPUT39), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n661), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n294), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n675), .B(KEYINPUT40), .Z(new_n676));
  INV_X1    g490(.A(new_n530), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n556), .A2(new_n520), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n189), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(G472), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n543), .A2(new_n549), .A3(new_n550), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n371), .B(KEYINPUT38), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n422), .A2(new_n478), .ZN(new_n683));
  INV_X1    g497(.A(new_n187), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n654), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n676), .A2(new_n681), .A3(new_n682), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G143), .ZN(G45));
  INV_X1    g501(.A(new_n611), .ZN(new_n688));
  AOI211_X1 g502(.A(new_n688), .B(new_n608), .C1(new_n609), .C2(new_n418), .ZN(new_n689));
  OAI211_X1 g503(.A(new_n478), .B(new_n662), .C1(new_n689), .C2(new_n606), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n659), .A2(new_n690), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n658), .A2(new_n691), .A3(new_n561), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT102), .B(G146), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G48));
  NOR2_X1   g508(.A1(new_n279), .A2(new_n282), .ZN(new_n695));
  OAI21_X1  g509(.A(G469), .B1(new_n695), .B2(G902), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n696), .A2(new_n293), .A3(new_n283), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n627), .A2(new_n561), .A3(new_n594), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT41), .B(G113), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G15));
  NAND4_X1  g514(.A1(new_n637), .A2(new_n561), .A3(new_n594), .A4(new_n697), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G116), .ZN(G18));
  AND3_X1   g516(.A1(new_n626), .A2(new_n187), .A3(new_n697), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n703), .A2(new_n561), .A3(new_n484), .A4(new_n654), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G119), .ZN(G21));
  NAND4_X1  g519(.A1(new_n626), .A2(new_n187), .A3(new_n478), .A4(new_n422), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n557), .A2(new_n540), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n534), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(G472), .A2(G902), .ZN(new_n709));
  AOI22_X1  g523(.A1(new_n599), .A2(G472), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  AND4_X1   g524(.A1(new_n293), .A2(new_n696), .A3(new_n283), .A4(new_n633), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(new_n711), .A3(new_n594), .ZN(new_n712));
  OR3_X1    g526(.A1(new_n706), .A2(KEYINPUT103), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g527(.A(KEYINPUT103), .B1(new_n706), .B2(new_n712), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G122), .ZN(G24));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n690), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n616), .A2(KEYINPUT104), .A3(new_n478), .A4(new_n662), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n710), .A2(new_n718), .A3(new_n654), .A4(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n703), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n626), .A2(new_n187), .A3(new_n697), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT105), .B1(new_n720), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G125), .ZN(G27));
  OR3_X1    g541(.A1(new_n542), .A2(KEYINPUT109), .A3(KEYINPUT32), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT109), .B1(new_n542), .B2(KEYINPUT32), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n728), .A2(new_n550), .A3(new_n560), .A4(new_n729), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n730), .A2(new_n594), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n718), .A2(new_n719), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n367), .A2(new_n187), .A3(new_n370), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT107), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT107), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n367), .A2(new_n736), .A3(new_n187), .A4(new_n370), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n289), .B(KEYINPUT106), .ZN(new_n738));
  AND4_X1   g552(.A1(new_n293), .A2(new_n735), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n731), .A2(KEYINPUT42), .A3(new_n733), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n561), .A2(new_n594), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n735), .A2(new_n738), .A3(new_n293), .A4(new_n737), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n741), .A2(new_n742), .A3(new_n732), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n744), .A3(KEYINPUT42), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n739), .A2(new_n561), .A3(new_n594), .A4(new_n733), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT42), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT108), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n740), .B1(new_n745), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G131), .ZN(G33));
  NOR3_X1   g564(.A1(new_n741), .A2(new_n742), .A3(new_n669), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n225), .ZN(G36));
  XNOR2_X1  g566(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n753));
  OR2_X1    g567(.A1(KEYINPUT111), .A2(KEYINPUT43), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n612), .A2(new_n478), .ZN(new_n755));
  MUX2_X1   g569(.A(new_n753), .B(new_n754), .S(new_n755), .Z(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(new_n601), .A3(new_n654), .ZN(new_n757));
  XOR2_X1   g571(.A(new_n757), .B(KEYINPUT44), .Z(new_n758));
  NAND2_X1  g572(.A1(new_n735), .A2(new_n737), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n284), .B1(new_n286), .B2(new_n265), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT45), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(G469), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n288), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT110), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n763), .A2(new_n767), .A3(new_n764), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n762), .A2(KEYINPUT46), .A3(new_n288), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n766), .A2(new_n283), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n293), .A3(new_n674), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n758), .A2(new_n759), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(new_n228), .ZN(G39));
  NOR4_X1   g587(.A1(new_n561), .A2(new_n759), .A3(new_n594), .A4(new_n690), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT47), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n770), .A2(new_n293), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n776), .A2(KEYINPUT112), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(KEYINPUT112), .ZN(new_n778));
  AOI211_X1 g592(.A(KEYINPUT113), .B(new_n775), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n775), .A2(KEYINPUT113), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT47), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n777), .A2(new_n780), .A3(new_n778), .A4(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n774), .B1(new_n779), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G140), .ZN(G42));
  AND2_X1   g600(.A1(new_n696), .A2(new_n283), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT114), .ZN(new_n788));
  XOR2_X1   g602(.A(new_n788), .B(KEYINPUT49), .Z(new_n789));
  INV_X1    g603(.A(new_n681), .ZN(new_n790));
  INV_X1    g604(.A(new_n682), .ZN(new_n791));
  AND4_X1   g605(.A1(new_n594), .A2(new_n755), .A3(new_n187), .A4(new_n293), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n789), .A2(new_n790), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n777), .A2(new_n780), .A3(new_n778), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n781), .A3(KEYINPUT47), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n795), .B(new_n783), .C1(new_n293), .C2(new_n788), .ZN(new_n796));
  INV_X1    g610(.A(new_n759), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n756), .A2(new_n594), .A3(new_n480), .A4(new_n710), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n796), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(KEYINPUT119), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n797), .A2(new_n293), .A3(new_n787), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(new_n594), .A3(new_n480), .A4(new_n790), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n803), .A2(new_n478), .A3(new_n616), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n791), .A2(new_n684), .A3(new_n697), .ZN(new_n805));
  OAI21_X1  g619(.A(KEYINPUT118), .B1(new_n805), .B2(new_n798), .ZN(new_n806));
  XOR2_X1   g620(.A(new_n806), .B(KEYINPUT50), .Z(new_n807));
  NAND2_X1  g621(.A1(new_n710), .A2(new_n654), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n802), .A2(new_n480), .A3(new_n756), .ZN(new_n810));
  AOI211_X1 g624(.A(new_n804), .B(new_n807), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n800), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n801), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n800), .B(new_n811), .C1(KEYINPUT119), .C2(KEYINPUT51), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n810), .A2(new_n731), .ZN(new_n816));
  XOR2_X1   g630(.A(new_n816), .B(KEYINPUT48), .Z(new_n817));
  AOI21_X1  g631(.A(new_n803), .B1(new_n613), .B2(new_n617), .ZN(new_n818));
  OAI211_X1 g632(.A(G952), .B(new_n263), .C1(new_n798), .C2(new_n724), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n814), .A2(new_n815), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n561), .B(new_n658), .C1(new_n670), .C2(new_n691), .ZN(new_n823));
  INV_X1    g637(.A(new_n706), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n293), .A2(new_n662), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n654), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n738), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n824), .A2(new_n681), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n722), .B1(new_n721), .B2(new_n703), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n720), .A2(new_n724), .A3(KEYINPUT105), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n823), .B(new_n828), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n726), .A2(KEYINPUT52), .A3(new_n828), .A4(new_n823), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n635), .A2(new_n662), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n659), .A2(new_n422), .A3(new_n836), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n797), .A2(new_n837), .A3(new_n561), .ZN(new_n838));
  AOI211_X1 g652(.A(new_n838), .B(new_n751), .C1(new_n721), .C2(new_n739), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n749), .A2(new_n835), .A3(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n715), .A2(new_n698), .A3(new_n701), .A4(new_n704), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(KEYINPUT115), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n698), .A2(new_n704), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n843), .A2(new_n844), .A3(new_n701), .A4(new_n715), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n604), .A2(new_n612), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n846), .B1(new_n604), .B2(new_n422), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n371), .A2(new_n187), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n847), .A2(new_n848), .A3(new_n483), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n602), .A2(new_n849), .A3(new_n628), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n850), .A2(new_n595), .A3(new_n655), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n842), .A2(new_n845), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n822), .B1(new_n840), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT116), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT54), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n850), .A2(KEYINPUT53), .A3(new_n595), .A4(new_n655), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n841), .A2(new_n856), .ZN(new_n857));
  AND4_X1   g671(.A1(new_n749), .A2(new_n857), .A3(new_n835), .A4(new_n839), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n860), .B(new_n822), .C1(new_n840), .C2(new_n852), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n854), .A2(new_n855), .A3(new_n859), .A4(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n749), .A2(new_n839), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n842), .A2(new_n845), .A3(new_n851), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT53), .A4(new_n835), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n853), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT54), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT117), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT117), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n862), .A2(new_n867), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n821), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(G952), .A2(G953), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n793), .B1(new_n873), .B2(new_n874), .ZN(G75));
  NOR2_X1   g689(.A1(new_n263), .A2(G952), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n858), .B1(new_n853), .B2(KEYINPUT116), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n189), .B1(new_n878), .B2(new_n861), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT56), .B1(new_n879), .B2(G210), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n362), .A2(new_n363), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(new_n364), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT55), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n877), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT56), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n879), .A2(G210), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n886), .B1(new_n887), .B2(KEYINPUT120), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n887), .A2(KEYINPUT120), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n884), .B1(new_n888), .B2(new_n889), .ZN(G51));
  INV_X1    g704(.A(new_n695), .ZN(new_n891));
  AOI211_X1 g705(.A(KEYINPUT121), .B(new_n855), .C1(new_n878), .C2(new_n861), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n878), .A2(new_n861), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT54), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n862), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n892), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n288), .B(KEYINPUT57), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n891), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n879), .A2(G469), .A3(new_n761), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n876), .B1(new_n899), .B2(new_n900), .ZN(G54));
  NAND2_X1  g715(.A1(new_n468), .A2(new_n469), .ZN(new_n902));
  NAND2_X1  g716(.A1(KEYINPUT58), .A2(G475), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT122), .Z(new_n904));
  AND3_X1   g718(.A1(new_n879), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n902), .B1(new_n879), .B2(new_n904), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n905), .A2(new_n906), .A3(new_n876), .ZN(G60));
  NAND2_X1  g721(.A1(G478), .A2(G902), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT59), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n610), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n877), .B1(new_n897), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n610), .B1(new_n872), .B2(new_n909), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n911), .A2(new_n912), .ZN(G63));
  XNOR2_X1  g727(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n408), .A2(new_n189), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n914), .B(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n917), .B1(new_n878), .B2(new_n861), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n876), .B1(new_n919), .B2(new_n586), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT124), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n918), .A2(new_n921), .A3(new_n650), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n921), .B1(new_n918), .B2(new_n650), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n920), .B(KEYINPUT61), .C1(new_n922), .C2(new_n923), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(G66));
  NAND3_X1  g742(.A1(new_n852), .A2(KEYINPUT125), .A3(new_n263), .ZN(new_n929));
  OAI21_X1  g743(.A(G953), .B1(new_n482), .B2(new_n325), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT125), .B1(new_n852), .B2(new_n263), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n881), .B1(G898), .B2(new_n263), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n933), .B(new_n934), .Z(G69));
  NAND2_X1  g749(.A1(new_n527), .A2(new_n528), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(new_n462), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(G900), .B2(G953), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n726), .A2(new_n823), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n731), .A2(new_n824), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n771), .A2(new_n940), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n772), .A2(new_n941), .A3(new_n751), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n785), .A2(new_n749), .A3(new_n939), .A4(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n938), .B1(new_n943), .B2(G953), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n939), .A2(new_n686), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT62), .Z(new_n946));
  XNOR2_X1  g760(.A(new_n847), .B(KEYINPUT126), .ZN(new_n947));
  NOR4_X1   g761(.A1(new_n947), .A2(new_n741), .A3(new_n675), .A4(new_n759), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n772), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n785), .A2(new_n946), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n263), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n951), .A2(new_n952), .A3(new_n937), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n952), .B1(new_n951), .B2(new_n937), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n944), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n263), .B1(G227), .B2(G900), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n956), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n958), .B(new_n944), .C1(new_n953), .C2(new_n954), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n959), .ZN(G72));
  NAND2_X1  g774(.A1(new_n516), .A2(new_n529), .ZN(new_n961));
  OR2_X1    g775(.A1(new_n943), .A2(new_n852), .ZN(new_n962));
  NAND2_X1  g776(.A1(G472), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT63), .Z(new_n964));
  AOI211_X1 g778(.A(new_n520), .B(new_n961), .C1(new_n962), .C2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n961), .A2(new_n520), .ZN(new_n966));
  OR2_X1    g780(.A1(new_n950), .A2(new_n852), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n966), .B1(new_n967), .B2(new_n964), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n964), .B1(new_n677), .B2(new_n553), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n865), .B2(new_n853), .ZN(new_n970));
  NOR4_X1   g784(.A1(new_n965), .A2(new_n968), .A3(new_n876), .A4(new_n970), .ZN(G57));
endmodule


