

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X1 U325 ( .A(n378), .B(n377), .ZN(n381) );
  XNOR2_X1 U326 ( .A(n376), .B(KEYINPUT11), .ZN(n377) );
  NOR2_X1 U327 ( .A1(n545), .A2(n457), .ZN(n531) );
  XNOR2_X1 U328 ( .A(n447), .B(n446), .ZN(n449) );
  OR2_X1 U329 ( .A1(n459), .A2(n458), .ZN(n293) );
  XOR2_X1 U330 ( .A(n372), .B(n371), .Z(n294) );
  NOR2_X1 U331 ( .A1(n364), .A2(n581), .ZN(n365) );
  XNOR2_X1 U332 ( .A(n387), .B(n386), .ZN(n388) );
  INV_X1 U333 ( .A(KEYINPUT23), .ZN(n434) );
  XNOR2_X1 U334 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n407) );
  XNOR2_X1 U335 ( .A(n435), .B(n434), .ZN(n436) );
  INV_X1 U336 ( .A(KEYINPUT32), .ZN(n340) );
  XNOR2_X1 U337 ( .A(n437), .B(n436), .ZN(n441) );
  XNOR2_X1 U338 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U339 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U340 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U341 ( .A(n470), .B(KEYINPUT97), .ZN(n485) );
  XNOR2_X1 U342 ( .A(KEYINPUT38), .B(n490), .ZN(n499) );
  XNOR2_X1 U343 ( .A(n453), .B(G190GAT), .ZN(n454) );
  XNOR2_X1 U344 ( .A(n455), .B(n454), .ZN(G1351GAT) );
  XOR2_X1 U345 ( .A(G176GAT), .B(G183GAT), .Z(n296) );
  XNOR2_X1 U346 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U348 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n298) );
  XNOR2_X1 U349 ( .A(G190GAT), .B(KEYINPUT84), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U351 ( .A(n300), .B(n299), .Z(n401) );
  XOR2_X1 U352 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n302) );
  NAND2_X1 U353 ( .A1(G227GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U354 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U355 ( .A(n303), .B(KEYINPUT65), .Z(n308) );
  XOR2_X1 U356 ( .A(G127GAT), .B(KEYINPUT81), .Z(n305) );
  XNOR2_X1 U357 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n305), .B(n304), .ZN(n427) );
  XNOR2_X1 U359 ( .A(G99GAT), .B(G120GAT), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n306), .B(G71GAT), .ZN(n337) );
  XNOR2_X1 U361 ( .A(n427), .B(n337), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U363 ( .A(n309), .B(KEYINPUT20), .Z(n311) );
  XOR2_X1 U364 ( .A(G43GAT), .B(G134GAT), .Z(n368) );
  XNOR2_X1 U365 ( .A(G15GAT), .B(n368), .ZN(n310) );
  XNOR2_X1 U366 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X2 U367 ( .A(n401), .B(n312), .Z(n529) );
  XOR2_X1 U368 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n318) );
  XOR2_X1 U369 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n314) );
  XNOR2_X1 U370 ( .A(G197GAT), .B(G22GAT), .ZN(n313) );
  XNOR2_X1 U371 ( .A(n314), .B(n313), .ZN(n316) );
  XNOR2_X1 U372 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n315) );
  XNOR2_X1 U373 ( .A(n315), .B(KEYINPUT8), .ZN(n371) );
  XNOR2_X1 U374 ( .A(n316), .B(n371), .ZN(n317) );
  XNOR2_X1 U375 ( .A(n318), .B(n317), .ZN(n324) );
  XOR2_X1 U376 ( .A(G15GAT), .B(KEYINPUT69), .Z(n320) );
  XNOR2_X1 U377 ( .A(G1GAT), .B(G8GAT), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n320), .B(n319), .ZN(n359) );
  XOR2_X1 U379 ( .A(G50GAT), .B(n359), .Z(n322) );
  NAND2_X1 U380 ( .A1(G229GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U381 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U382 ( .A(n324), .B(n323), .Z(n329) );
  XOR2_X1 U383 ( .A(G113GAT), .B(G141GAT), .Z(n326) );
  XNOR2_X1 U384 ( .A(G169GAT), .B(G43GAT), .ZN(n325) );
  XNOR2_X1 U385 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U386 ( .A(n327), .B(G36GAT), .ZN(n328) );
  XOR2_X1 U387 ( .A(n329), .B(n328), .Z(n572) );
  INV_X1 U388 ( .A(n572), .ZN(n559) );
  XNOR2_X1 U389 ( .A(G92GAT), .B(G64GAT), .ZN(n330) );
  XNOR2_X1 U390 ( .A(n330), .B(G204GAT), .ZN(n402) );
  XNOR2_X1 U391 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n331) );
  XOR2_X1 U392 ( .A(n331), .B(KEYINPUT13), .Z(n358) );
  XNOR2_X1 U393 ( .A(n402), .B(n358), .ZN(n345) );
  NAND2_X1 U394 ( .A1(G230GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U395 ( .A(KEYINPUT73), .B(KEYINPUT33), .ZN(n332) );
  XOR2_X1 U396 ( .A(n333), .B(n332), .Z(n334) );
  XOR2_X1 U397 ( .A(n334), .B(KEYINPUT31), .Z(n339) );
  XOR2_X1 U398 ( .A(KEYINPUT71), .B(G78GAT), .Z(n336) );
  XNOR2_X1 U399 ( .A(G148GAT), .B(G106GAT), .ZN(n335) );
  XNOR2_X1 U400 ( .A(n336), .B(n335), .ZN(n443) );
  XNOR2_X1 U401 ( .A(n337), .B(n443), .ZN(n338) );
  XNOR2_X1 U402 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U403 ( .A(G85GAT), .B(KEYINPUT72), .Z(n372) );
  XNOR2_X1 U404 ( .A(G176GAT), .B(n372), .ZN(n341) );
  XNOR2_X1 U405 ( .A(n345), .B(n344), .ZN(n577) );
  XNOR2_X1 U406 ( .A(KEYINPUT41), .B(n577), .ZN(n563) );
  NOR2_X1 U407 ( .A1(n559), .A2(n563), .ZN(n346) );
  XNOR2_X1 U408 ( .A(n346), .B(KEYINPUT46), .ZN(n364) );
  XOR2_X1 U409 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n348) );
  XNOR2_X1 U410 ( .A(G71GAT), .B(G78GAT), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n348), .B(n347), .ZN(n363) );
  XNOR2_X1 U412 ( .A(G22GAT), .B(G155GAT), .ZN(n448) );
  XOR2_X1 U413 ( .A(G211GAT), .B(G64GAT), .Z(n350) );
  XNOR2_X1 U414 ( .A(G183GAT), .B(G127GAT), .ZN(n349) );
  XNOR2_X1 U415 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U416 ( .A(n448), .B(n351), .ZN(n353) );
  NAND2_X1 U417 ( .A1(G231GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U418 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U419 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n355) );
  XNOR2_X1 U420 ( .A(KEYINPUT78), .B(KEYINPUT15), .ZN(n354) );
  XNOR2_X1 U421 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U422 ( .A(n357), .B(n356), .Z(n361) );
  XOR2_X1 U423 ( .A(n359), .B(n358), .Z(n360) );
  XNOR2_X1 U424 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U425 ( .A(n363), .B(n362), .Z(n567) );
  INV_X1 U426 ( .A(n567), .ZN(n581) );
  XNOR2_X1 U427 ( .A(n365), .B(KEYINPUT112), .ZN(n384) );
  XOR2_X1 U428 ( .A(KEYINPUT10), .B(KEYINPUT75), .Z(n367) );
  XNOR2_X1 U429 ( .A(G190GAT), .B(KEYINPUT74), .ZN(n366) );
  XNOR2_X1 U430 ( .A(n367), .B(n366), .ZN(n383) );
  XOR2_X1 U431 ( .A(G50GAT), .B(G162GAT), .Z(n444) );
  XOR2_X1 U432 ( .A(n444), .B(G106GAT), .Z(n370) );
  XNOR2_X1 U433 ( .A(n368), .B(KEYINPUT76), .ZN(n369) );
  XNOR2_X1 U434 ( .A(n370), .B(n369), .ZN(n375) );
  NAND2_X1 U435 ( .A1(G232GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U436 ( .A(n294), .B(n373), .ZN(n374) );
  XNOR2_X1 U437 ( .A(n375), .B(n374), .ZN(n378) );
  XOR2_X1 U438 ( .A(G99GAT), .B(G92GAT), .Z(n376) );
  XNOR2_X1 U439 ( .A(G36GAT), .B(G218GAT), .ZN(n379) );
  XNOR2_X1 U440 ( .A(n379), .B(KEYINPUT77), .ZN(n396) );
  XOR2_X1 U441 ( .A(n396), .B(KEYINPUT9), .Z(n380) );
  XNOR2_X1 U442 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U443 ( .A(n383), .B(n382), .ZN(n540) );
  INV_X1 U444 ( .A(n540), .ZN(n556) );
  NAND2_X1 U445 ( .A1(n384), .A2(n556), .ZN(n385) );
  XNOR2_X1 U446 ( .A(n385), .B(KEYINPUT47), .ZN(n391) );
  XNOR2_X1 U447 ( .A(KEYINPUT36), .B(n540), .ZN(n584) );
  NAND2_X1 U448 ( .A1(n584), .A2(n581), .ZN(n387) );
  XOR2_X1 U449 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n386) );
  NAND2_X1 U450 ( .A1(n388), .A2(n559), .ZN(n389) );
  NOR2_X1 U451 ( .A1(n577), .A2(n389), .ZN(n390) );
  NOR2_X1 U452 ( .A1(n391), .A2(n390), .ZN(n392) );
  XNOR2_X1 U453 ( .A(KEYINPUT48), .B(n392), .ZN(n528) );
  XOR2_X1 U454 ( .A(KEYINPUT91), .B(KEYINPUT93), .Z(n394) );
  NAND2_X1 U455 ( .A1(G226GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U456 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U457 ( .A(KEYINPUT92), .B(n395), .Z(n398) );
  XNOR2_X1 U458 ( .A(G8GAT), .B(n396), .ZN(n397) );
  XNOR2_X1 U459 ( .A(n398), .B(n397), .ZN(n400) );
  XNOR2_X1 U460 ( .A(G197GAT), .B(G211GAT), .ZN(n399) );
  XNOR2_X1 U461 ( .A(n399), .B(KEYINPUT21), .ZN(n442) );
  XOR2_X1 U462 ( .A(n400), .B(n442), .Z(n405) );
  INV_X1 U463 ( .A(n401), .ZN(n403) );
  XOR2_X1 U464 ( .A(n403), .B(n402), .Z(n404) );
  XOR2_X1 U465 ( .A(n405), .B(n404), .Z(n477) );
  XNOR2_X1 U466 ( .A(KEYINPUT119), .B(n477), .ZN(n406) );
  NOR2_X1 U467 ( .A1(n528), .A2(n406), .ZN(n408) );
  XNOR2_X1 U468 ( .A(n408), .B(n407), .ZN(n432) );
  XOR2_X1 U469 ( .A(KEYINPUT5), .B(G57GAT), .Z(n410) );
  XNOR2_X1 U470 ( .A(KEYINPUT1), .B(KEYINPUT86), .ZN(n409) );
  XNOR2_X1 U471 ( .A(n410), .B(n409), .ZN(n414) );
  XOR2_X1 U472 ( .A(G155GAT), .B(KEYINPUT90), .Z(n412) );
  XNOR2_X1 U473 ( .A(G120GAT), .B(KEYINPUT4), .ZN(n411) );
  XNOR2_X1 U474 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U475 ( .A(n414), .B(n413), .Z(n419) );
  XOR2_X1 U476 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n416) );
  NAND2_X1 U477 ( .A1(G225GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U478 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U479 ( .A(G148GAT), .B(n417), .ZN(n418) );
  XNOR2_X1 U480 ( .A(n419), .B(n418), .ZN(n431) );
  XOR2_X1 U481 ( .A(G162GAT), .B(G85GAT), .Z(n421) );
  XNOR2_X1 U482 ( .A(G134GAT), .B(KEYINPUT76), .ZN(n420) );
  XNOR2_X1 U483 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U484 ( .A(KEYINPUT6), .B(KEYINPUT89), .Z(n423) );
  XNOR2_X1 U485 ( .A(G29GAT), .B(G1GAT), .ZN(n422) );
  XNOR2_X1 U486 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U487 ( .A(n425), .B(n424), .Z(n429) );
  XNOR2_X1 U488 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n426) );
  XNOR2_X1 U489 ( .A(n426), .B(KEYINPUT2), .ZN(n437) );
  XNOR2_X1 U490 ( .A(n427), .B(n437), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U492 ( .A(n431), .B(n430), .Z(n474) );
  INV_X1 U493 ( .A(n474), .ZN(n545) );
  NAND2_X1 U494 ( .A1(n432), .A2(n545), .ZN(n433) );
  XNOR2_X1 U495 ( .A(n433), .B(KEYINPUT64), .ZN(n570) );
  NAND2_X1 U496 ( .A1(G228GAT), .A2(G233GAT), .ZN(n435) );
  XOR2_X1 U497 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n439) );
  XNOR2_X1 U498 ( .A(G204GAT), .B(G218GAT), .ZN(n438) );
  XNOR2_X1 U499 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U500 ( .A(n441), .B(n440), .Z(n447) );
  XNOR2_X1 U501 ( .A(n443), .B(n442), .ZN(n445) );
  XNOR2_X1 U502 ( .A(n449), .B(n448), .ZN(n463) );
  NOR2_X1 U503 ( .A1(n570), .A2(n463), .ZN(n450) );
  XNOR2_X1 U504 ( .A(n450), .B(KEYINPUT55), .ZN(n451) );
  NOR2_X1 U505 ( .A1(n529), .A2(n451), .ZN(n452) );
  XNOR2_X1 U506 ( .A(n452), .B(KEYINPUT121), .ZN(n566) );
  NOR2_X1 U507 ( .A1(n566), .A2(n556), .ZN(n455) );
  XNOR2_X1 U508 ( .A(KEYINPUT123), .B(KEYINPUT58), .ZN(n453) );
  NOR2_X1 U509 ( .A1(n559), .A2(n577), .ZN(n489) );
  INV_X1 U510 ( .A(n529), .ZN(n480) );
  XOR2_X1 U511 ( .A(n480), .B(KEYINPUT85), .Z(n459) );
  XNOR2_X1 U512 ( .A(n477), .B(KEYINPUT94), .ZN(n456) );
  XOR2_X1 U513 ( .A(KEYINPUT27), .B(n456), .Z(n461) );
  XNOR2_X1 U514 ( .A(KEYINPUT28), .B(n463), .ZN(n498) );
  OR2_X1 U515 ( .A1(n461), .A2(n498), .ZN(n457) );
  XNOR2_X1 U516 ( .A(KEYINPUT95), .B(n531), .ZN(n458) );
  NAND2_X1 U517 ( .A1(n463), .A2(n529), .ZN(n460) );
  XNOR2_X1 U518 ( .A(n460), .B(KEYINPUT26), .ZN(n569) );
  NOR2_X1 U519 ( .A1(n569), .A2(n461), .ZN(n547) );
  INV_X1 U520 ( .A(n477), .ZN(n517) );
  NOR2_X1 U521 ( .A1(n529), .A2(n517), .ZN(n462) );
  NOR2_X1 U522 ( .A1(n463), .A2(n462), .ZN(n464) );
  XOR2_X1 U523 ( .A(KEYINPUT25), .B(n464), .Z(n465) );
  NOR2_X1 U524 ( .A1(n547), .A2(n465), .ZN(n466) );
  NOR2_X1 U525 ( .A1(n474), .A2(n466), .ZN(n467) );
  XNOR2_X1 U526 ( .A(KEYINPUT96), .B(n467), .ZN(n468) );
  INV_X1 U527 ( .A(n468), .ZN(n469) );
  NAND2_X1 U528 ( .A1(n293), .A2(n469), .ZN(n470) );
  NOR2_X1 U529 ( .A1(n567), .A2(n540), .ZN(n471) );
  XOR2_X1 U530 ( .A(KEYINPUT16), .B(n471), .Z(n472) );
  NOR2_X1 U531 ( .A1(n485), .A2(n472), .ZN(n502) );
  NAND2_X1 U532 ( .A1(n489), .A2(n502), .ZN(n473) );
  XOR2_X1 U533 ( .A(KEYINPUT98), .B(n473), .Z(n483) );
  NAND2_X1 U534 ( .A1(n483), .A2(n474), .ZN(n475) );
  XNOR2_X1 U535 ( .A(n475), .B(KEYINPUT34), .ZN(n476) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(n476), .ZN(G1324GAT) );
  XOR2_X1 U537 ( .A(G8GAT), .B(KEYINPUT99), .Z(n479) );
  NAND2_X1 U538 ( .A1(n483), .A2(n477), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n479), .B(n478), .ZN(G1325GAT) );
  XOR2_X1 U540 ( .A(G15GAT), .B(KEYINPUT35), .Z(n482) );
  NAND2_X1 U541 ( .A1(n483), .A2(n480), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n482), .B(n481), .ZN(G1326GAT) );
  NAND2_X1 U543 ( .A1(n483), .A2(n498), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n484), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U545 ( .A1(n485), .A2(n581), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n486), .B(KEYINPUT100), .ZN(n487) );
  NAND2_X1 U547 ( .A1(n487), .A2(n584), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n488), .B(KEYINPUT37), .ZN(n514) );
  NAND2_X1 U549 ( .A1(n514), .A2(n489), .ZN(n490) );
  NOR2_X1 U550 ( .A1(n499), .A2(n545), .ZN(n492) );
  XNOR2_X1 U551 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(G1328GAT) );
  XNOR2_X1 U553 ( .A(G36GAT), .B(KEYINPUT101), .ZN(n494) );
  NOR2_X1 U554 ( .A1(n517), .A2(n499), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(G1329GAT) );
  XNOR2_X1 U556 ( .A(KEYINPUT40), .B(KEYINPUT102), .ZN(n496) );
  NOR2_X1 U557 ( .A1(n529), .A2(n499), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U559 ( .A(G43GAT), .B(n497), .Z(G1330GAT) );
  INV_X1 U560 ( .A(n498), .ZN(n525) );
  NOR2_X1 U561 ( .A1(n499), .A2(n525), .ZN(n501) );
  XNOR2_X1 U562 ( .A(G50GAT), .B(KEYINPUT103), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(G1331GAT) );
  NOR2_X1 U564 ( .A1(n563), .A2(n572), .ZN(n513) );
  NAND2_X1 U565 ( .A1(n513), .A2(n502), .ZN(n510) );
  NOR2_X1 U566 ( .A1(n545), .A2(n510), .ZN(n504) );
  XNOR2_X1 U567 ( .A(KEYINPUT42), .B(KEYINPUT104), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U569 ( .A(G57GAT), .B(n505), .Z(G1332GAT) );
  NOR2_X1 U570 ( .A1(n517), .A2(n510), .ZN(n507) );
  XNOR2_X1 U571 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U573 ( .A(G64GAT), .B(n508), .ZN(G1333GAT) );
  NOR2_X1 U574 ( .A1(n529), .A2(n510), .ZN(n509) );
  XOR2_X1 U575 ( .A(G71GAT), .B(n509), .Z(G1334GAT) );
  NOR2_X1 U576 ( .A1(n525), .A2(n510), .ZN(n512) );
  XNOR2_X1 U577 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  NAND2_X1 U579 ( .A1(n514), .A2(n513), .ZN(n524) );
  NOR2_X1 U580 ( .A1(n545), .A2(n524), .ZN(n516) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(KEYINPUT107), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(G1336GAT) );
  NOR2_X1 U583 ( .A1(n517), .A2(n524), .ZN(n518) );
  XOR2_X1 U584 ( .A(KEYINPUT108), .B(n518), .Z(n519) );
  XNOR2_X1 U585 ( .A(G92GAT), .B(n519), .ZN(G1337GAT) );
  NOR2_X1 U586 ( .A1(n529), .A2(n524), .ZN(n521) );
  XNOR2_X1 U587 ( .A(G99GAT), .B(KEYINPUT109), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(G1338GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT110), .B(KEYINPUT44), .Z(n523) );
  XNOR2_X1 U590 ( .A(G106GAT), .B(KEYINPUT111), .ZN(n522) );
  XNOR2_X1 U591 ( .A(n523), .B(n522), .ZN(n527) );
  NOR2_X1 U592 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U593 ( .A(n527), .B(n526), .Z(G1339GAT) );
  NOR2_X1 U594 ( .A1(n528), .A2(n529), .ZN(n530) );
  NAND2_X1 U595 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U596 ( .A(KEYINPUT113), .B(n532), .ZN(n541) );
  NAND2_X1 U597 ( .A1(n572), .A2(n541), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n533), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT49), .Z(n536) );
  INV_X1 U600 ( .A(n563), .ZN(n534) );
  NAND2_X1 U601 ( .A1(n541), .A2(n534), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(G1341GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n538) );
  NAND2_X1 U604 ( .A1(n541), .A2(n581), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U606 ( .A(G127GAT), .B(n539), .Z(G1342GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U608 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U610 ( .A(G134GAT), .B(n544), .Z(G1343GAT) );
  NOR2_X1 U611 ( .A1(n545), .A2(n528), .ZN(n546) );
  NAND2_X1 U612 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U613 ( .A(KEYINPUT116), .B(n548), .ZN(n555) );
  NOR2_X1 U614 ( .A1(n559), .A2(n555), .ZN(n549) );
  XOR2_X1 U615 ( .A(G141GAT), .B(n549), .Z(G1344GAT) );
  NOR2_X1 U616 ( .A1(n555), .A2(n563), .ZN(n553) );
  XOR2_X1 U617 ( .A(KEYINPUT117), .B(KEYINPUT52), .Z(n551) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  NOR2_X1 U621 ( .A1(n567), .A2(n555), .ZN(n554) );
  XOR2_X1 U622 ( .A(G155GAT), .B(n554), .Z(G1346GAT) );
  NOR2_X1 U623 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U624 ( .A(KEYINPUT118), .B(n557), .Z(n558) );
  XNOR2_X1 U625 ( .A(G162GAT), .B(n558), .ZN(G1347GAT) );
  NOR2_X1 U626 ( .A1(n559), .A2(n566), .ZN(n560) );
  XOR2_X1 U627 ( .A(G169GAT), .B(n560), .Z(G1348GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT122), .B(KEYINPUT56), .Z(n562) );
  XNOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(n565) );
  NOR2_X1 U631 ( .A1(n563), .A2(n566), .ZN(n564) );
  XOR2_X1 U632 ( .A(n565), .B(n564), .Z(G1349GAT) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U634 ( .A(G183GAT), .B(n568), .Z(G1350GAT) );
  NOR2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(KEYINPUT124), .B(n571), .ZN(n583) );
  AND2_X1 U637 ( .A1(n583), .A2(n572), .ZN(n576) );
  XOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n574) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n579) );
  NAND2_X1 U643 ( .A1(n583), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(n580), .ZN(G1353GAT) );
  NAND2_X1 U646 ( .A1(n583), .A2(n581), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n586) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

