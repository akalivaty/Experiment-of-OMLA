//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  XOR2_X1   g0011(.A(KEYINPUT65), .B(G238), .Z(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G107), .A2(G264), .ZN(new_n218));
  NAND4_X1  g0018(.A1(new_n215), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n211), .B1(new_n214), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT66), .Z(new_n222));
  NOR2_X1   g0022(.A1(new_n211), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT0), .ZN(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT64), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n228), .A2(new_n209), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n225), .B(new_n230), .C1(KEYINPUT1), .C2(new_n220), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n222), .A2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT67), .Z(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n236), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XOR2_X1   g0045(.A(new_n245), .B(KEYINPUT68), .Z(new_n246));
  NAND2_X1  g0046(.A1(new_n202), .A2(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n213), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n246), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(G13), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G1), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT71), .ZN(new_n256));
  NOR3_X1   g0056(.A1(new_n253), .A2(new_n209), .A3(G1), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT71), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n228), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n208), .A2(G20), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(G68), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n256), .A2(new_n259), .ZN(new_n266));
  OAI21_X1  g0066(.A(KEYINPUT12), .B1(new_n266), .B2(G68), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n213), .A2(G20), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT12), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n254), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n267), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G20), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G50), .ZN(new_n273));
  INV_X1    g0073(.A(G77), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n209), .A2(G33), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n273), .B(new_n268), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n262), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n277), .B(KEYINPUT11), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n265), .A2(new_n271), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G238), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT69), .ZN(new_n285));
  INV_X1    g0085(.A(G33), .ZN(new_n286));
  INV_X1    g0086(.A(G41), .ZN(new_n287));
  OAI211_X1 g0087(.A(G1), .B(G13), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(KEYINPUT69), .B1(new_n288), .B2(new_n282), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n280), .B1(new_n285), .B2(new_n290), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n288), .A2(G274), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n283), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G226), .A2(G1698), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n294), .B1(new_n238), .B2(G1698), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT3), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n286), .ZN(new_n297));
  NAND2_X1  g0097(.A1(KEYINPUT3), .A2(G33), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n295), .A2(new_n299), .B1(G33), .B2(G97), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n293), .B1(new_n300), .B2(new_n288), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT13), .B1(new_n291), .B2(new_n301), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n300), .A2(new_n288), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT69), .ZN(new_n304));
  NOR3_X1   g0104(.A1(new_n281), .A2(new_n283), .A3(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(G238), .B1(new_n305), .B2(new_n289), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT13), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n303), .A2(new_n306), .A3(new_n307), .A4(new_n293), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n279), .B1(new_n309), .B2(G200), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n302), .A2(KEYINPUT72), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT72), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n312), .B(KEYINPUT13), .C1(new_n291), .C2(new_n301), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n311), .A2(G190), .A3(new_n313), .A4(new_n308), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n309), .A2(G169), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT73), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT14), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n311), .A2(G179), .A3(new_n313), .A4(new_n308), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(KEYINPUT14), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n309), .A2(G169), .A3(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n316), .B1(new_n323), .B2(new_n279), .ZN(new_n324));
  AND2_X1   g0124(.A1(KEYINPUT3), .A2(G33), .ZN(new_n325));
  NOR2_X1   g0125(.A1(KEYINPUT3), .A2(G33), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G107), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n299), .A2(G1698), .ZN(new_n329));
  INV_X1    g0129(.A(G1698), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n299), .A2(new_n330), .ZN(new_n331));
  OAI221_X1 g0131(.A(new_n328), .B1(new_n329), .B2(new_n212), .C1(new_n238), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n281), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n285), .A2(new_n290), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G244), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(new_n293), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G169), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n263), .A2(G77), .A3(new_n264), .ZN(new_n339));
  XOR2_X1   g0139(.A(KEYINPUT8), .B(G58), .Z(new_n340));
  AOI22_X1  g0140(.A1(new_n340), .A2(new_n272), .B1(G20), .B2(G77), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT15), .B(G87), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n341), .B1(new_n275), .B2(new_n342), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n343), .A2(new_n262), .B1(new_n274), .B2(new_n260), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n338), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n336), .ZN(new_n347));
  INV_X1    g0147(.A(G179), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G200), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G190), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n339), .B(new_n344), .C1(new_n336), .C2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n324), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT16), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n297), .A2(new_n209), .A3(new_n298), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT7), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n297), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n298), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n213), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G58), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n365), .A2(new_n213), .ZN(new_n366));
  OAI21_X1  g0166(.A(G20), .B1(new_n366), .B2(new_n201), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n272), .A2(G159), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n359), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n262), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n367), .A2(KEYINPUT16), .A3(new_n368), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT74), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n363), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n327), .A2(KEYINPUT74), .A3(KEYINPUT7), .A4(new_n209), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n374), .A2(new_n375), .A3(new_n362), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n372), .B1(new_n376), .B2(G68), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT75), .B1(new_n371), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n377), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT75), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n379), .A2(new_n380), .A3(new_n262), .A4(new_n370), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n257), .A2(new_n262), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n340), .A2(new_n264), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n384), .A2(new_n385), .B1(new_n255), .B2(new_n340), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  OAI211_X1 g0187(.A(G226), .B(G1698), .C1(new_n325), .C2(new_n326), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT76), .ZN(new_n389));
  XNOR2_X1  g0189(.A(new_n388), .B(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n327), .A2(G1698), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n391), .A2(G223), .B1(G33), .B2(G87), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n288), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n283), .A2(new_n292), .B1(new_n284), .B2(G232), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n352), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G223), .ZN(new_n397));
  INV_X1    g0197(.A(G87), .ZN(new_n398));
  OAI22_X1  g0198(.A1(new_n331), .A2(new_n397), .B1(new_n286), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n388), .A2(new_n389), .ZN(new_n400));
  OR2_X1    g0200(.A1(new_n388), .A2(new_n389), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n394), .B1(new_n402), .B2(new_n288), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n354), .A2(KEYINPUT77), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n354), .A2(KEYINPUT77), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n396), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n382), .A2(new_n387), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT17), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n262), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT7), .B1(new_n327), .B2(new_n209), .ZN(new_n413));
  INV_X1    g0213(.A(new_n363), .ZN(new_n414));
  OAI21_X1  g0214(.A(G68), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n369), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n412), .B1(new_n417), .B2(new_n359), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n380), .B1(new_n418), .B2(new_n379), .ZN(new_n419));
  NOR3_X1   g0219(.A1(new_n371), .A2(KEYINPUT75), .A3(new_n377), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n387), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT18), .ZN(new_n422));
  OAI21_X1  g0222(.A(G169), .B1(new_n393), .B2(new_n395), .ZN(new_n423));
  OAI211_X1 g0223(.A(G179), .B(new_n394), .C1(new_n402), .C2(new_n288), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n421), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n386), .B1(new_n378), .B2(new_n381), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n423), .A2(new_n424), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT18), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n427), .A2(KEYINPUT17), .A3(new_n408), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n411), .A2(new_n426), .A3(new_n429), .A4(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n327), .A2(G77), .ZN(new_n433));
  INV_X1    g0233(.A(G222), .ZN(new_n434));
  OAI221_X1 g0234(.A(new_n433), .B1(new_n329), .B2(new_n397), .C1(new_n434), .C2(new_n331), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n281), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n334), .A2(G226), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n293), .A3(new_n437), .ZN(new_n438));
  OR2_X1    g0238(.A1(new_n438), .A2(G179), .ZN(new_n439));
  INV_X1    g0239(.A(new_n275), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n340), .A2(new_n440), .B1(G150), .B2(new_n272), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n203), .A2(G20), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n412), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(KEYINPUT70), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(KEYINPUT70), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n202), .B1(new_n208), .B2(G20), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n383), .A2(new_n447), .B1(new_n202), .B2(new_n257), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n445), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n438), .A2(new_n337), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n439), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n446), .A2(new_n448), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT9), .B1(new_n453), .B2(new_n444), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT9), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n445), .A2(new_n455), .A3(new_n446), .A4(new_n448), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n438), .A2(G200), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n436), .A2(G190), .A3(new_n293), .A4(new_n437), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT10), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n454), .A2(new_n456), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT10), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n462), .A2(new_n463), .A3(new_n458), .A4(new_n459), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n452), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n358), .A2(KEYINPUT78), .A3(new_n432), .A4(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT78), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n324), .A2(new_n357), .A3(new_n465), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n467), .B1(new_n468), .B2(new_n431), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n327), .A2(new_n330), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n471), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n299), .A2(G244), .A3(new_n330), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT4), .ZN(new_n474));
  OAI21_X1  g0274(.A(KEYINPUT79), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT79), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n391), .A2(new_n476), .A3(KEYINPUT4), .A4(G244), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n473), .A2(new_n474), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n472), .A2(new_n475), .A3(new_n477), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n281), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT5), .B(G41), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n208), .A2(G45), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n288), .ZN(new_n485));
  INV_X1    g0285(.A(G257), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n292), .A2(new_n483), .A3(new_n481), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n480), .A2(new_n348), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(G107), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(KEYINPUT6), .A3(G97), .ZN(new_n492));
  INV_X1    g0292(.A(G97), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n493), .A2(new_n491), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(new_n205), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n492), .B1(new_n495), .B2(KEYINPUT6), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n496), .A2(G20), .B1(G77), .B2(new_n272), .ZN(new_n497));
  OAI21_X1  g0297(.A(G107), .B1(new_n413), .B2(new_n414), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n412), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n257), .A2(new_n493), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n208), .A2(G33), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n383), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n500), .B1(new_n502), .B2(new_n493), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n288), .A2(G274), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n484), .A2(new_n506), .ZN(new_n507));
  AOI211_X1 g0307(.A(new_n487), .B(new_n507), .C1(new_n479), .C2(new_n281), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n490), .B(new_n505), .C1(new_n508), .C2(G169), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n299), .A2(new_n209), .A3(G68), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT19), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n275), .B2(new_n493), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n209), .A2(new_n514), .B1(new_n205), .B2(new_n398), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n262), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n260), .A2(new_n342), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n383), .A2(G87), .A3(new_n501), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n288), .A2(G250), .A3(new_n482), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n506), .B2(new_n482), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n299), .A2(G238), .A3(new_n330), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G33), .A2(G116), .ZN(new_n523));
  INV_X1    g0323(.A(G244), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n522), .B(new_n523), .C1(new_n329), .C2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n521), .B1(new_n525), .B2(new_n281), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G190), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n519), .B(new_n527), .C1(new_n352), .C2(new_n526), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n516), .B(new_n517), .C1(new_n342), .C2(new_n502), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n526), .A2(new_n348), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n529), .B(new_n530), .C1(G169), .C2(new_n526), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n480), .A2(G190), .A3(new_n488), .A4(new_n489), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n533), .B(new_n504), .C1(new_n508), .C2(new_n352), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n509), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n299), .A2(new_n209), .A3(G87), .ZN(new_n536));
  XOR2_X1   g0336(.A(KEYINPUT81), .B(KEYINPUT22), .Z(new_n537));
  OR2_X1    g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT22), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n536), .A2(KEYINPUT81), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n523), .A2(G20), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT23), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(new_n209), .B2(G107), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n491), .A2(KEYINPUT23), .A3(G20), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n538), .A2(new_n540), .A3(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT24), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n538), .A2(KEYINPUT24), .A3(new_n540), .A4(new_n545), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n548), .A2(new_n262), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n383), .A2(G107), .A3(new_n501), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT82), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n552), .B(KEYINPUT25), .C1(new_n255), .C2(G107), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT25), .ZN(new_n554));
  AOI21_X1  g0354(.A(G107), .B1(new_n554), .B2(KEYINPUT82), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n257), .B(new_n555), .C1(KEYINPUT82), .C2(new_n554), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n551), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT83), .ZN(new_n558));
  XNOR2_X1  g0358(.A(new_n557), .B(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n550), .A2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(G264), .ZN(new_n561));
  OAI22_X1  g0361(.A1(new_n485), .A2(new_n561), .B1(new_n506), .B2(new_n484), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n299), .A2(G257), .A3(G1698), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n299), .A2(G250), .A3(new_n330), .ZN(new_n564));
  NAND2_X1  g0364(.A1(G33), .A2(G294), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT84), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n288), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT84), .A4(new_n565), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n562), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n348), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n568), .A2(new_n569), .ZN(new_n572));
  INV_X1    g0372(.A(new_n562), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n337), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n560), .A2(new_n571), .A3(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT21), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n266), .A2(G116), .A3(new_n412), .A4(new_n501), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(G116), .B2(new_n266), .ZN(new_n580));
  AOI21_X1  g0380(.A(G20), .B1(G33), .B2(G283), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(G33), .B2(new_n493), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n582), .B(new_n262), .C1(new_n209), .C2(G116), .ZN(new_n583));
  XNOR2_X1  g0383(.A(new_n583), .B(KEYINPUT20), .ZN(new_n584));
  OAI21_X1  g0384(.A(G169), .B1(new_n580), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(G270), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n489), .B1(new_n586), .B2(new_n485), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n327), .A2(new_n486), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n588), .A2(new_n330), .B1(G303), .B2(new_n327), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT80), .B1(new_n471), .B2(G264), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT80), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n329), .A2(new_n591), .A3(new_n561), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n589), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n587), .B1(new_n593), .B2(new_n281), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n578), .B1(new_n585), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT20), .ZN(new_n596));
  XNOR2_X1  g0396(.A(new_n583), .B(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n597), .B(new_n579), .C1(G116), .C2(new_n266), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n598), .A2(G179), .A3(new_n594), .ZN(new_n599));
  INV_X1    g0399(.A(new_n485), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n507), .B1(new_n600), .B2(G270), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n299), .A2(G257), .ZN(new_n602));
  INV_X1    g0402(.A(G303), .ZN(new_n603));
  OAI22_X1  g0403(.A1(new_n602), .A2(G1698), .B1(new_n603), .B2(new_n299), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n591), .B1(new_n329), .B2(new_n561), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n471), .A2(KEYINPUT80), .A3(G264), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n601), .B1(new_n607), .B2(new_n288), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n598), .A2(new_n608), .A3(KEYINPUT21), .A4(G169), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n595), .A2(new_n599), .A3(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n577), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n574), .A2(G200), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n570), .A2(G190), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n612), .A2(new_n559), .A3(new_n550), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n608), .A2(G200), .ZN(new_n615));
  INV_X1    g0415(.A(new_n598), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n615), .B(new_n616), .C1(new_n406), .C2(new_n608), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  AND4_X1   g0419(.A1(new_n470), .A2(new_n535), .A3(new_n611), .A4(new_n619), .ZN(G372));
  NAND4_X1  g0420(.A1(new_n509), .A2(new_n532), .A3(new_n534), .A4(new_n614), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n610), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT85), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(new_n624), .A3(new_n576), .ZN(new_n625));
  OAI21_X1  g0425(.A(KEYINPUT85), .B1(new_n577), .B2(new_n610), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n622), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n531), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n528), .A2(new_n531), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n629), .B1(new_n509), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n480), .A2(new_n488), .A3(new_n489), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n504), .B1(new_n632), .B2(new_n337), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n532), .A2(KEYINPUT26), .A3(new_n490), .A4(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n628), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n627), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n470), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n422), .B1(new_n421), .B2(new_n425), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n427), .A2(KEYINPUT18), .A3(new_n428), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n351), .A2(new_n315), .B1(new_n323), .B2(new_n279), .ZN(new_n641));
  AND4_X1   g0441(.A1(KEYINPUT17), .A2(new_n382), .A3(new_n387), .A4(new_n408), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT17), .B1(new_n427), .B2(new_n408), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n640), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n461), .A2(new_n464), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n452), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n637), .A2(new_n648), .ZN(G369));
  NAND2_X1  g0449(.A1(new_n254), .A2(new_n209), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(G213), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(G343), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n616), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n610), .B(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n658), .A2(new_n617), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n560), .A2(new_n655), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n577), .B1(new_n614), .B2(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n576), .A2(new_n655), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n659), .A2(G330), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n610), .A2(new_n656), .ZN(new_n666));
  OAI22_X1  g0466(.A1(new_n661), .A2(new_n666), .B1(new_n576), .B2(new_n655), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g0468(.A(new_n668), .B(KEYINPUT86), .Z(G399));
  INV_X1    g0469(.A(new_n223), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(G41), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G1), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n227), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n674), .B1(new_n675), .B2(new_n672), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT28), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n655), .B1(new_n627), .B2(new_n635), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT29), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n611), .A2(new_n621), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n655), .B1(new_n680), .B2(new_n635), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(KEYINPUT29), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT87), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n480), .A2(new_n488), .A3(new_n526), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n608), .A2(new_n348), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n685), .A2(new_n686), .A3(KEYINPUT30), .A4(new_n570), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT30), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n594), .A2(G179), .A3(new_n570), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n480), .A2(new_n488), .A3(new_n526), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n526), .A2(G179), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n632), .A2(new_n692), .A3(new_n608), .A4(new_n574), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n687), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n694), .A2(KEYINPUT31), .A3(new_n655), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(KEYINPUT31), .B1(new_n694), .B2(new_n655), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n684), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n694), .A2(new_n655), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT31), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(KEYINPUT87), .A3(new_n695), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n535), .A2(new_n611), .A3(new_n619), .A4(new_n656), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G330), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n683), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(KEYINPUT88), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT88), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n683), .A2(new_n709), .A3(new_n706), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n677), .B1(new_n711), .B2(G1), .ZN(G364));
  NOR2_X1   g0512(.A1(new_n253), .A2(G20), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n208), .B1(new_n713), .B2(G45), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n671), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n670), .A2(new_n327), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT89), .ZN(new_n719));
  XNOR2_X1  g0519(.A(G355), .B(KEYINPUT90), .ZN(new_n720));
  INV_X1    g0520(.A(G116), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n719), .A2(new_n720), .B1(new_n721), .B2(new_n670), .ZN(new_n722));
  INV_X1    g0522(.A(G45), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n251), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n670), .A2(new_n299), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(new_n675), .B2(G45), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n722), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(G13), .A2(G33), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G20), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n228), .B1(G20), .B2(new_n337), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n717), .B1(new_n727), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n730), .ZN(new_n734));
  OAI21_X1  g0534(.A(KEYINPUT92), .B1(new_n209), .B2(G190), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n209), .A2(KEYINPUT92), .A3(G190), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G179), .A2(G200), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g0541(.A(KEYINPUT93), .B(G159), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT94), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n744), .A2(KEYINPUT32), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n209), .A2(new_n348), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G200), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G190), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n209), .B1(new_n740), .B2(G190), .ZN(new_n750));
  OAI22_X1  g0550(.A1(new_n749), .A2(new_n213), .B1(new_n493), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n352), .A2(G179), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n753), .A2(new_n209), .A3(new_n354), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n406), .A2(new_n747), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n299), .B1(new_n755), .B2(new_n398), .C1(new_n757), .C2(new_n202), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n738), .A2(new_n753), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n751), .B(new_n758), .C1(G107), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n744), .A2(KEYINPUT32), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n746), .A2(KEYINPUT91), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n746), .A2(KEYINPUT91), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n763), .A2(new_n407), .A3(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n763), .A2(new_n354), .A3(new_n764), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(G58), .A2(new_n766), .B1(new_n768), .B2(G77), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n745), .A2(new_n760), .A3(new_n761), .A4(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT95), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n741), .A2(KEYINPUT97), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n741), .A2(KEYINPUT97), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G329), .ZN(new_n778));
  XNOR2_X1  g0578(.A(KEYINPUT33), .B(G317), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n756), .A2(G326), .B1(new_n748), .B2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G294), .ZN(new_n781));
  INV_X1    g0581(.A(G311), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n780), .B1(new_n781), .B2(new_n750), .C1(new_n782), .C2(new_n767), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(G322), .B2(new_n766), .ZN(new_n784));
  INV_X1    g0584(.A(new_n759), .ZN(new_n785));
  INV_X1    g0585(.A(G283), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n299), .B1(new_n754), .B2(G303), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n785), .A2(new_n786), .B1(new_n787), .B2(KEYINPUT96), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(KEYINPUT96), .B2(new_n787), .ZN(new_n789));
  AND3_X1   g0589(.A1(new_n778), .A2(new_n784), .A3(new_n789), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n772), .A2(new_n773), .A3(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n731), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n733), .B1(new_n659), .B2(new_n734), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n659), .A2(G330), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n717), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n659), .A2(G330), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n793), .B1(new_n795), .B2(new_n796), .ZN(G396));
  NAND2_X1  g0597(.A1(new_n345), .A2(new_n655), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(new_n353), .B2(new_n355), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n350), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n346), .A2(new_n349), .A3(new_n656), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n678), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n678), .A2(new_n803), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n717), .B1(new_n806), .B2(new_n706), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n807), .A2(KEYINPUT101), .B1(new_n706), .B2(new_n806), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(KEYINPUT101), .B2(new_n807), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n731), .A2(new_n728), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n717), .B1(new_n274), .B2(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n756), .A2(G137), .B1(new_n748), .B2(G150), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n742), .B2(new_n767), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(G143), .B2(new_n766), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT99), .Z(new_n815));
  INV_X1    g0615(.A(KEYINPUT34), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n299), .B1(new_n750), .B2(new_n365), .C1(new_n755), .C2(new_n202), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n785), .A2(new_n213), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(G132), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n820), .B1(new_n776), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(new_n815), .B2(new_n816), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n776), .A2(new_n782), .B1(new_n398), .B2(new_n785), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT98), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n767), .A2(new_n721), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n327), .B1(new_n750), .B2(new_n493), .C1(new_n755), .C2(new_n491), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n757), .A2(new_n603), .B1(new_n749), .B2(new_n786), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n765), .A2(new_n781), .ZN(new_n829));
  NOR4_X1   g0629(.A1(new_n826), .A2(new_n827), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n817), .A2(new_n823), .B1(new_n825), .B2(new_n830), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n811), .B1(new_n803), .B2(new_n729), .C1(new_n831), .C2(new_n792), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT100), .Z(new_n833));
  NAND2_X1  g0633(.A1(new_n809), .A2(new_n833), .ZN(G384));
  OR2_X1    g0634(.A1(new_n496), .A2(KEYINPUT35), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n496), .A2(KEYINPUT35), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n835), .A2(G116), .A3(new_n229), .A4(new_n836), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT36), .Z(new_n838));
  OAI211_X1 g0638(.A(new_n227), .B(G77), .C1(new_n365), .C2(new_n213), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n208), .B(G13), .C1(new_n839), .C2(new_n247), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n805), .A2(new_n801), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n279), .A2(new_n655), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n324), .A2(new_n843), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n279), .B(new_n655), .C1(new_n323), .C2(new_n316), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n653), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n379), .A2(new_n262), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n376), .A2(G68), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT16), .B1(new_n850), .B2(new_n416), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n387), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n431), .A2(new_n848), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n409), .B1(new_n427), .B2(new_n428), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT37), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n653), .B(KEYINPUT102), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n855), .B1(new_n427), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n423), .A2(new_n424), .A3(new_n653), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n427), .A2(new_n408), .B1(new_n852), .B2(new_n859), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n854), .A2(new_n858), .B1(new_n860), .B2(new_n855), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n853), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT38), .ZN(new_n863));
  OR2_X1    g0663(.A1(new_n860), .A2(new_n855), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n421), .A2(new_n425), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n421), .A2(new_n856), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n865), .A2(new_n866), .A3(new_n855), .A4(new_n409), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n863), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n862), .A2(new_n863), .B1(new_n853), .B2(new_n868), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n847), .A2(new_n869), .B1(new_n640), .B2(new_n856), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n861), .A2(KEYINPUT38), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n852), .A2(new_n848), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n640), .B2(new_n644), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT104), .ZN(new_n874));
  NOR3_X1   g0674(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT104), .B1(new_n868), .B2(new_n853), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n427), .A2(new_n857), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n431), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT103), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT103), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n431), .A2(new_n881), .A3(new_n878), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT37), .B1(new_n854), .B2(new_n878), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n867), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n880), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n863), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT105), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT39), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n877), .A2(new_n886), .A3(new_n887), .A4(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n874), .B1(new_n871), .B2(new_n873), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n868), .A2(KEYINPUT104), .A3(new_n853), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n890), .A2(new_n891), .A3(new_n888), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n879), .A2(KEYINPUT103), .B1(new_n867), .B2(new_n883), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT38), .B1(new_n893), .B2(new_n882), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT105), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n869), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT39), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n889), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n323), .A2(new_n279), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n899), .A2(new_n655), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n870), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n679), .A2(new_n470), .A3(new_n682), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n648), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n901), .B(new_n903), .Z(new_n904));
  NAND3_X1  g0704(.A1(new_n704), .A2(new_n701), .A3(new_n695), .ZN(new_n905));
  AND4_X1   g0705(.A1(KEYINPUT40), .A2(new_n905), .A3(new_n846), .A4(new_n803), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n890), .A2(new_n891), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n906), .B1(new_n894), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT40), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n905), .A2(new_n846), .A3(new_n803), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n909), .B1(new_n869), .B2(new_n910), .ZN(new_n911));
  AND4_X1   g0711(.A1(new_n470), .A2(new_n908), .A3(new_n905), .A4(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n908), .A2(G330), .A3(new_n911), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n470), .A2(G330), .A3(new_n905), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n912), .B1(KEYINPUT106), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(KEYINPUT106), .B2(new_n915), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n904), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n208), .B2(new_n713), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n904), .A2(new_n917), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n841), .B1(new_n919), .B2(new_n920), .ZN(G367));
  OAI21_X1  g0721(.A(new_n327), .B1(new_n749), .B2(new_n781), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n785), .A2(new_n493), .ZN(new_n923));
  INV_X1    g0723(.A(new_n741), .ZN(new_n924));
  AOI211_X1 g0724(.A(new_n922), .B(new_n923), .C1(G317), .C2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n768), .A2(G283), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n766), .A2(G303), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n754), .A2(G116), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n928), .B(KEYINPUT46), .Z(new_n929));
  OAI22_X1  g0729(.A1(new_n757), .A2(new_n782), .B1(new_n491), .B2(new_n750), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n925), .A2(new_n926), .A3(new_n927), .A4(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n299), .B1(new_n755), .B2(new_n365), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(G143), .B2(new_n756), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n924), .A2(G137), .B1(new_n759), .B2(G77), .ZN(new_n935));
  INV_X1    g0735(.A(new_n742), .ZN(new_n936));
  INV_X1    g0736(.A(new_n750), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n748), .A2(new_n936), .B1(G68), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n934), .A2(new_n935), .A3(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(G150), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n202), .A2(new_n767), .B1(new_n765), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n932), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n943));
  XNOR2_X1  g0743(.A(new_n942), .B(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n731), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n519), .A2(new_n656), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n630), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n628), .A2(new_n946), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n947), .A2(new_n730), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n725), .A2(new_n235), .ZN(new_n950));
  INV_X1    g0750(.A(new_n732), .ZN(new_n951));
  INV_X1    g0751(.A(new_n342), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n951), .B1(new_n670), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n717), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n945), .A2(new_n949), .A3(new_n954), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n509), .B(new_n534), .C1(new_n504), .C2(new_n656), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n633), .A2(new_n490), .A3(new_n655), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n667), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT45), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n667), .A2(new_n959), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT44), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(new_n665), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n794), .B(KEYINPUT108), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n663), .B(new_n666), .Z(new_n968));
  AND2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n968), .B1(KEYINPUT108), .B2(new_n794), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n711), .B1(new_n966), .B2(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n671), .B(KEYINPUT41), .Z(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n715), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  OR3_X1    g0775(.A1(new_n664), .A2(KEYINPUT107), .A3(new_n959), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT107), .B1(new_n664), .B2(new_n959), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n947), .A2(new_n948), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n979), .A2(KEYINPUT43), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n978), .A2(new_n980), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n663), .A2(new_n610), .A3(new_n656), .A4(new_n958), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n984), .A2(KEYINPUT42), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n956), .A2(new_n576), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n655), .B1(new_n986), .B2(new_n509), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(new_n984), .B2(KEYINPUT42), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n985), .A2(new_n988), .B1(KEYINPUT43), .B2(new_n979), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n983), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n981), .A2(new_n989), .A3(new_n982), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n955), .B1(new_n975), .B2(new_n993), .ZN(G387));
  NAND3_X1  g0794(.A1(new_n971), .A2(new_n710), .A3(new_n708), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n969), .A2(new_n970), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n672), .B1(new_n711), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n725), .B1(new_n241), .B2(new_n723), .ZN(new_n999));
  INV_X1    g0799(.A(new_n719), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n999), .B1(new_n1000), .B2(new_n673), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n340), .ZN(new_n1002));
  OR3_X1    g0802(.A1(new_n1002), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1003));
  OAI21_X1  g0803(.A(KEYINPUT50), .B1(new_n1002), .B2(G50), .ZN(new_n1004));
  AOI21_X1  g0804(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1003), .A2(new_n673), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n1001), .A2(new_n1006), .B1(new_n491), .B2(new_n670), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n716), .B1(new_n1007), .B2(new_n951), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n755), .A2(new_n274), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(new_n924), .B2(G150), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT110), .ZN(new_n1011));
  INV_X1    g0811(.A(G159), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n299), .B1(new_n757), .B2(new_n1012), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n749), .A2(new_n1002), .B1(new_n342), .B2(new_n750), .ZN(new_n1014));
  NOR3_X1   g0814(.A1(new_n923), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G50), .A2(new_n766), .B1(new_n768), .B2(G68), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1011), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n299), .B1(new_n924), .B2(G326), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n755), .A2(new_n781), .B1(new_n750), .B2(new_n786), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n756), .A2(G322), .B1(new_n748), .B2(G311), .ZN(new_n1020));
  INV_X1    g0820(.A(G317), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1020), .B1(new_n765), .B2(new_n1021), .C1(new_n603), .C2(new_n767), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT48), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1019), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n1023), .B2(new_n1022), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT49), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1018), .B1(new_n721), .B2(new_n785), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1017), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1008), .B1(new_n1029), .B2(new_n731), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n663), .B2(new_n734), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n998), .B(new_n1031), .C1(new_n714), .C2(new_n971), .ZN(G393));
  XNOR2_X1  g0832(.A(new_n965), .B(new_n664), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n959), .A2(new_n730), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n725), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n732), .B1(new_n493), .B2(new_n223), .C1(new_n1035), .C2(new_n245), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n716), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n327), .B1(new_n749), .B2(new_n603), .C1(new_n786), .C2(new_n755), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(G116), .B2(new_n937), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n924), .A2(G322), .B1(new_n759), .B2(G107), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(new_n781), .C2(new_n767), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n765), .A2(new_n782), .B1(new_n757), .B2(new_n1021), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT52), .Z(new_n1043));
  NOR2_X1   g0843(.A1(new_n750), .A2(new_n274), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n299), .B1(new_n755), .B2(new_n213), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1044), .B(new_n1045), .C1(G50), .C2(new_n748), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n924), .A2(G143), .B1(new_n759), .B2(G87), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1046), .B(new_n1047), .C1(new_n1002), .C2(new_n767), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n765), .A2(new_n1012), .B1(new_n757), .B2(new_n940), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT51), .Z(new_n1050));
  OAI22_X1  g0850(.A1(new_n1041), .A2(new_n1043), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1037), .B1(new_n1051), .B2(new_n731), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n1033), .A2(new_n715), .B1(new_n1034), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n711), .A2(new_n996), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n671), .B1(new_n1054), .B2(new_n966), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1033), .B1(new_n711), .B2(new_n996), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1053), .B1(new_n1055), .B2(new_n1056), .ZN(G390));
  INV_X1    g0857(.A(new_n900), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n801), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n678), .B2(new_n803), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n846), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1058), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n889), .A2(new_n895), .A3(new_n897), .A4(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(G330), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n802), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n705), .A2(new_n846), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1059), .B1(new_n681), .B2(new_n800), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1058), .B1(new_n1067), .B2(new_n1061), .C1(new_n894), .C2(new_n907), .ZN(new_n1068));
  AND3_X1   g0868(.A1(new_n1063), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n910), .A2(new_n1064), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n1063), .B2(new_n1068), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n902), .A2(new_n914), .A3(new_n648), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1065), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n703), .B2(new_n704), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1070), .B1(new_n846), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n681), .A2(new_n800), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n801), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n1074), .B2(new_n846), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n905), .A2(new_n1065), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n1061), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT111), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1079), .A2(KEYINPUT111), .A3(new_n1061), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n1075), .A2(new_n842), .B1(new_n1078), .B2(new_n1084), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n1069), .A2(new_n1071), .B1(new_n1072), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1063), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1074), .A2(new_n846), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n910), .A2(new_n1064), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n842), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1083), .ZN(new_n1091));
  AOI21_X1  g0891(.A(KEYINPUT111), .B1(new_n1079), .B2(new_n1061), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1066), .B(new_n1067), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1072), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n1063), .A2(new_n1068), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1087), .B(new_n1094), .C1(new_n1095), .C2(new_n1070), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1086), .A2(new_n1096), .A3(new_n671), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n810), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n716), .B1(new_n340), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n777), .A2(G294), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n819), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n757), .A2(new_n786), .B1(new_n749), .B2(new_n491), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n327), .B1(new_n755), .B2(new_n398), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n1103), .A2(new_n1104), .A3(new_n1044), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G97), .A2(new_n768), .B1(new_n766), .B2(G116), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1101), .A2(new_n1102), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n777), .A2(G125), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n766), .A2(G132), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n299), .B1(new_n750), .B2(new_n1012), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n756), .B2(G128), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT53), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n755), .B2(new_n940), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n754), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1113), .A2(new_n1114), .B1(G50), .B2(new_n759), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1108), .A2(new_n1109), .A3(new_n1111), .A4(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT54), .B(G143), .ZN(new_n1117));
  INV_X1    g0917(.A(G137), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n767), .A2(new_n1117), .B1(new_n749), .B2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT112), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1107), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1100), .B1(new_n1121), .B2(new_n731), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n898), .B2(new_n729), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(KEYINPUT113), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT113), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1125), .B(new_n1122), .C1(new_n898), .C2(new_n729), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1098), .A2(new_n715), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1097), .A2(new_n1127), .ZN(G378));
  INV_X1    g0928(.A(new_n1072), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1096), .A2(new_n1129), .ZN(new_n1130));
  XOR2_X1   g0930(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n647), .A2(new_n451), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n449), .A2(new_n848), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT115), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n465), .A2(new_n1134), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1137), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1132), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1141), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1143), .A2(new_n1131), .A3(new_n1139), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1145), .A2(G330), .A3(new_n911), .A4(new_n908), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n913), .A2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n892), .A2(new_n894), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1149), .A2(new_n887), .B1(KEYINPUT39), .B2(new_n896), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1058), .B1(new_n1150), .B2(new_n895), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1146), .B(new_n1148), .C1(new_n1151), .C2(new_n870), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1148), .A2(new_n1146), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n901), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1152), .A2(KEYINPUT116), .A3(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1153), .A2(new_n901), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT116), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1130), .A2(new_n1155), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT57), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1160), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n672), .B1(new_n1162), .B2(new_n1130), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1155), .A2(new_n715), .A3(new_n1158), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n717), .B1(new_n202), .B2(new_n810), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n749), .A2(new_n821), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n755), .A2(new_n1117), .B1(new_n750), .B2(new_n940), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1167), .B(new_n1168), .C1(G125), .C2(new_n756), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n766), .A2(G128), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1169), .B(new_n1170), .C1(new_n1118), .C2(new_n767), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n1171), .A2(KEYINPUT59), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(KEYINPUT59), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n759), .A2(new_n936), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT114), .B(G124), .ZN(new_n1175));
  AOI211_X1 g0975(.A(G33), .B(G41), .C1(new_n924), .C2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .A4(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n299), .A2(G41), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1179), .B(new_n1009), .C1(G68), .C2(new_n937), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n759), .A2(G58), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n756), .A2(G116), .B1(new_n748), .B2(G97), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(G107), .A2(new_n766), .B1(new_n768), .B2(new_n952), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(new_n786), .C2(new_n776), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT58), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1179), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1189));
  AND4_X1   g0989(.A1(new_n1177), .A2(new_n1187), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1166), .B1(new_n792), .B2(new_n1190), .C1(new_n1147), .C2(new_n729), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1165), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1164), .A2(new_n1193), .ZN(G375));
  AOI21_X1  g0994(.A(new_n714), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1061), .A2(new_n728), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n716), .B1(G68), .B2(new_n1099), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT117), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n756), .A2(G294), .B1(new_n748), .B2(G116), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n754), .A2(G97), .B1(new_n952), .B2(new_n937), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(new_n786), .C2(new_n765), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(G107), .B2(new_n768), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n299), .B1(new_n759), .B2(G77), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT118), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1202), .B(new_n1204), .C1(new_n603), .C2(new_n776), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT119), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n777), .A2(G128), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n299), .B1(new_n755), .B2(new_n1012), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n757), .A2(new_n821), .B1(new_n749), .B2(new_n1117), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1209), .B(new_n1210), .C1(G50), .C2(new_n937), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(G137), .A2(new_n766), .B1(new_n768), .B2(G150), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1208), .A2(new_n1181), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1207), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1198), .B1(new_n1215), .B2(new_n731), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1196), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(KEYINPUT120), .B1(new_n1195), .B2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT120), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1220), .B(new_n1217), .C1(new_n1085), .C2(new_n714), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1094), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1090), .A2(new_n1093), .A3(new_n1072), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1223), .A2(new_n974), .A3(new_n1224), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1222), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(G381));
  INV_X1    g1027(.A(G387), .ZN(new_n1228));
  INV_X1    g1028(.A(G384), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1229), .B(new_n1053), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(G393), .A2(G396), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1228), .A2(new_n1231), .A3(new_n1232), .A4(new_n1226), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT121), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1192), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1235));
  INV_X1    g1035(.A(G378), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1234), .A2(new_n1238), .ZN(G407));
  INV_X1    g1039(.A(G213), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(new_n1234), .B2(new_n1238), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1240), .A2(G343), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1235), .A2(new_n1236), .A3(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT122), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1243), .B(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1241), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT123), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1241), .A2(new_n1245), .A3(KEYINPUT123), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(G409));
  INV_X1    g1050(.A(G390), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(G387), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(KEYINPUT125), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(G393), .B(G396), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1228), .A2(G390), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1252), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1253), .A2(new_n1254), .A3(new_n1256), .A4(new_n1252), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G375), .A2(G378), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1153), .A2(new_n901), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n715), .B1(new_n1263), .B2(new_n1156), .ZN(new_n1264));
  AND4_X1   g1064(.A1(new_n1097), .A2(new_n1127), .A3(new_n1264), .A4(new_n1191), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1130), .A2(new_n1155), .A3(new_n974), .A4(new_n1158), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1242), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1090), .A2(new_n1072), .A3(new_n1093), .A4(KEYINPUT60), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1268), .A2(new_n671), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT60), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1224), .B1(new_n1094), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n1272), .A2(new_n1222), .A3(G384), .ZN(new_n1273));
  AOI21_X1  g1073(.A(G384), .B1(new_n1272), .B2(new_n1222), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  AND2_X1   g1075(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1262), .A2(new_n1267), .A3(new_n1275), .A4(new_n1278), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1267), .B(new_n1275), .C1(new_n1235), .C2(new_n1236), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1276), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1267), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1282));
  OAI21_X1  g1082(.A(KEYINPUT124), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1272), .A2(new_n1222), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1229), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT124), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1272), .A2(new_n1222), .A3(G384), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1285), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1242), .A2(G2897), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1283), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1275), .A2(new_n1286), .A3(G2897), .A4(new_n1242), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(KEYINPUT61), .B1(new_n1282), .B2(new_n1292), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1279), .B(new_n1281), .C1(new_n1293), .C2(KEYINPUT126), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT126), .ZN(new_n1295));
  AOI211_X1 g1095(.A(new_n1295), .B(KEYINPUT61), .C1(new_n1282), .C2(new_n1292), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1261), .B1(new_n1294), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT63), .ZN(new_n1298));
  OR2_X1    g1098(.A1(new_n1280), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1280), .A2(new_n1298), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1299), .A2(new_n1260), .A3(new_n1293), .A4(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1297), .A2(new_n1301), .ZN(G405));
  NAND2_X1  g1102(.A1(new_n1262), .A2(new_n1237), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1261), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1303), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1305), .A2(new_n1260), .ZN(new_n1306));
  OAI22_X1  g1106(.A1(new_n1304), .A2(new_n1306), .B1(new_n1274), .B2(new_n1273), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1261), .A2(new_n1303), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1305), .A2(new_n1260), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1308), .A2(new_n1275), .A3(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1307), .A2(new_n1310), .ZN(G402));
endmodule


