//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 0 1 1 0 0 1 1 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n806, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n993, new_n994, new_n995,
    new_n996;
  INV_X1    g000(.A(KEYINPUT88), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT35), .ZN(new_n203));
  INV_X1    g002(.A(G134gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G127gat), .ZN(new_n205));
  INV_X1    g004(.A(G127gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G134gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT70), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n210));
  OAI22_X1  g009(.A1(new_n210), .A2(KEYINPUT71), .B1(G113gat), .B2(G120gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT71), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n212), .A2(KEYINPUT1), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  AND2_X1   g013(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n216));
  OAI21_X1  g015(.A(G113gat), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT70), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n205), .A2(new_n207), .A3(new_n218), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n209), .A2(new_n214), .A3(new_n217), .A4(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(KEYINPUT67), .A2(G127gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT68), .ZN(new_n222));
  NAND2_X1  g021(.A1(KEYINPUT67), .A2(G127gat), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n221), .A2(new_n222), .A3(G134gat), .A4(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT1), .B1(G113gat), .B2(G120gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G113gat), .B2(G120gat), .ZN(new_n226));
  AND2_X1   g025(.A1(KEYINPUT67), .A2(G127gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(KEYINPUT67), .A2(G127gat), .ZN(new_n228));
  NOR3_X1   g027(.A1(new_n227), .A2(new_n228), .A3(new_n204), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n205), .A2(KEYINPUT68), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n224), .B(new_n226), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n220), .A2(new_n231), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n232), .A2(KEYINPUT72), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT27), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n234), .A2(G183gat), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(G190gat), .B1(new_n234), .B2(G183gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(KEYINPUT28), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G190gat), .ZN(new_n239));
  INV_X1    g038(.A(G183gat), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n240), .B2(KEYINPUT27), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT65), .B(G183gat), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n241), .B1(new_n242), .B2(KEYINPUT27), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n238), .B1(new_n243), .B2(KEYINPUT28), .ZN(new_n244));
  NAND2_X1  g043(.A1(G183gat), .A2(G190gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(G169gat), .A2(G176gat), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT26), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G169gat), .ZN(new_n249));
  INV_X1    g048(.A(G176gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n248), .A2(KEYINPUT66), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(G169gat), .A2(G176gat), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n247), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n252), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n244), .A2(new_n245), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT25), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n249), .A2(KEYINPUT64), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT64), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G169gat), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n261), .A2(new_n263), .A3(KEYINPUT23), .A4(new_n250), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n246), .A2(KEYINPUT23), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(new_n251), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(G183gat), .A2(G190gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n245), .A2(KEYINPUT24), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT24), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(G183gat), .A3(G190gat), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n268), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n260), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n242), .A2(new_n239), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n269), .A2(new_n271), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n255), .B1(KEYINPUT23), .B2(new_n246), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n249), .A2(new_n250), .A3(KEYINPUT23), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT25), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n273), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n259), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n232), .A2(KEYINPUT72), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n233), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n259), .A2(new_n282), .A3(KEYINPUT72), .A4(new_n232), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT34), .ZN(new_n288));
  NAND2_X1  g087(.A1(G227gat), .A2(G233gat), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n288), .B1(new_n287), .B2(new_n289), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n285), .A2(G227gat), .A3(G233gat), .A4(new_n286), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT32), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT33), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(G15gat), .B(G43gat), .Z(new_n297));
  XNOR2_X1  g096(.A(G71gat), .B(G99gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n294), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n299), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n293), .B(KEYINPUT32), .C1(new_n295), .C2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n292), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n292), .A2(new_n300), .A3(new_n302), .ZN(new_n305));
  XNOR2_X1  g104(.A(G197gat), .B(G204gat), .ZN(new_n306));
  INV_X1    g105(.A(G211gat), .ZN(new_n307));
  INV_X1    g106(.A(G218gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n306), .B1(KEYINPUT22), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G211gat), .B(G218gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT3), .ZN(new_n313));
  NAND2_X1  g112(.A1(G155gat), .A2(G162gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G141gat), .B(G148gat), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n317), .B1(new_n318), .B2(KEYINPUT2), .ZN(new_n319));
  INV_X1    g118(.A(G148gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G141gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  AND2_X1   g121(.A1(KEYINPUT76), .A2(G141gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(KEYINPUT76), .A2(G141gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n322), .B1(new_n325), .B2(G148gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT2), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n316), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(new_n314), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n313), .B(new_n319), .C1(new_n326), .C2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n312), .B1(new_n332), .B2(KEYINPUT29), .ZN(new_n333));
  INV_X1    g132(.A(new_n312), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT29), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT3), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT76), .ZN(new_n337));
  INV_X1    g136(.A(G141gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(KEYINPUT76), .A2(G141gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(G148gat), .A3(new_n340), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n341), .A2(new_n321), .B1(new_n314), .B2(new_n328), .ZN(new_n342));
  XNOR2_X1  g141(.A(G155gat), .B(G162gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n338), .A2(G148gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n321), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n343), .B1(new_n327), .B2(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n333), .B1(new_n336), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G78gat), .B(G106gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G228gat), .A2(G233gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(G22gat), .ZN(new_n352));
  XOR2_X1   g151(.A(KEYINPUT31), .B(G50gat), .Z(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n350), .B(new_n354), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n304), .A2(new_n305), .A3(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n347), .A2(new_n231), .A3(new_n220), .A4(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT3), .B1(new_n342), .B2(new_n346), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n232), .A2(new_n359), .A3(new_n331), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n341), .A2(new_n321), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n329), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(new_n319), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT4), .B1(new_n232), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n358), .B1(new_n360), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G225gat), .A2(G233gat), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n367), .A2(KEYINPUT5), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n357), .B1(new_n232), .B2(new_n363), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n232), .A2(new_n359), .A3(new_n331), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n347), .A2(KEYINPUT4), .A3(new_n231), .A4(new_n220), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n370), .A2(new_n371), .A3(new_n366), .A4(new_n372), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n232), .A2(new_n363), .ZN(new_n374));
  AOI22_X1  g173(.A1(new_n231), .A2(new_n220), .B1(new_n362), .B2(new_n319), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n367), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n373), .A2(KEYINPUT5), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n369), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G1gat), .B(G29gat), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT0), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G57gat), .B(G85gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n381), .B(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n378), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT6), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n369), .A2(new_n377), .A3(new_n383), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n373), .A2(KEYINPUT5), .A3(new_n376), .ZN(new_n389));
  INV_X1    g188(.A(new_n368), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n347), .A2(new_n231), .A3(new_n220), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n371), .A2(KEYINPUT4), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n390), .B1(new_n392), .B2(new_n358), .ZN(new_n393));
  OAI211_X1 g192(.A(KEYINPUT6), .B(new_n384), .C1(new_n389), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT78), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT78), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n378), .A2(new_n396), .A3(KEYINPUT6), .A4(new_n384), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n388), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G8gat), .B(G36gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(G64gat), .B(G92gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n400), .B(new_n401), .Z(new_n402));
  INV_X1    g201(.A(KEYINPUT28), .ZN(new_n403));
  NOR3_X1   g202(.A1(new_n241), .A2(new_n235), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n240), .A2(KEYINPUT65), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT65), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(G183gat), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n407), .A3(KEYINPUT27), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n237), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n404), .B1(new_n409), .B2(new_n403), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n258), .A2(new_n245), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n240), .A2(KEYINPUT24), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n413), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n245), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n266), .B(new_n264), .C1(new_n414), .C2(new_n268), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n415), .A2(new_n260), .B1(new_n276), .B2(new_n280), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT74), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT74), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n259), .A2(new_n282), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(G226gat), .ZN(new_n420));
  INV_X1    g219(.A(G233gat), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n422), .A2(KEYINPUT29), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n417), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n259), .A2(new_n282), .A3(new_n422), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(new_n312), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n423), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n427), .B1(new_n259), .B2(new_n282), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n417), .A2(new_n419), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n428), .B1(new_n429), .B2(new_n422), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n402), .B(new_n426), .C1(new_n430), .C2(new_n312), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT30), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n422), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n434), .B1(new_n417), .B2(new_n419), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n334), .B1(new_n435), .B2(new_n428), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n436), .A2(KEYINPUT30), .A3(new_n402), .A4(new_n426), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n426), .ZN(new_n438));
  XOR2_X1   g237(.A(new_n402), .B(KEYINPUT75), .Z(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n433), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n399), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n203), .B1(new_n356), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT73), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n305), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n292), .A2(new_n300), .A3(KEYINPUT73), .A4(new_n302), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n447), .A2(new_n203), .A3(new_n304), .A4(new_n355), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT80), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n441), .A2(new_n450), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n431), .A2(new_n432), .B1(new_n438), .B2(new_n439), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n452), .A2(KEYINPUT80), .A3(new_n437), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT5), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n232), .A2(new_n363), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n391), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n455), .B1(new_n457), .B2(new_n367), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n373), .A2(new_n458), .B1(new_n365), .B2(new_n368), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT81), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n383), .B(new_n460), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n387), .B(new_n386), .C1(new_n459), .C2(new_n461), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n395), .A2(new_n397), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT86), .B1(new_n454), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT86), .ZN(new_n466));
  AOI211_X1 g265(.A(new_n466), .B(new_n463), .C1(new_n451), .C2(new_n453), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n449), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT87), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT80), .B1(new_n452), .B2(new_n437), .ZN(new_n470));
  AND4_X1   g269(.A1(KEYINPUT80), .A2(new_n433), .A3(new_n437), .A4(new_n440), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n466), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n454), .A2(KEYINPUT86), .A3(new_n464), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT87), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(new_n476), .A3(new_n449), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n443), .B1(new_n469), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n304), .A2(KEYINPUT36), .A3(new_n305), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n303), .B1(new_n445), .B2(new_n446), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n479), .B1(new_n480), .B2(KEYINPUT36), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT79), .ZN(new_n482));
  INV_X1    g281(.A(new_n355), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n483), .B1(new_n399), .B2(new_n441), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n459), .A2(new_n461), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT39), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n392), .A2(new_n488), .A3(new_n367), .A4(new_n358), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n461), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT82), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT39), .B1(new_n457), .B2(new_n367), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT83), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n494), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n495), .B(new_n496), .C1(new_n366), .C2(new_n365), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n487), .B1(new_n498), .B2(KEYINPUT40), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n492), .A2(new_n497), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT40), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n499), .A2(new_n451), .A3(new_n453), .A4(new_n502), .ZN(new_n503));
  XOR2_X1   g302(.A(KEYINPUT84), .B(KEYINPUT38), .Z(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(KEYINPUT85), .B(KEYINPUT37), .ZN(new_n506));
  OR2_X1    g305(.A1(new_n438), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n402), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n438), .A2(KEYINPUT37), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n505), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n424), .A2(new_n334), .A3(new_n425), .ZN(new_n512));
  OAI211_X1 g311(.A(KEYINPUT37), .B(new_n512), .C1(new_n430), .C2(new_n334), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n507), .A2(new_n439), .A3(new_n504), .A4(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n511), .A2(new_n463), .A3(new_n431), .A4(new_n514), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n503), .A2(new_n355), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n482), .B1(new_n481), .B2(new_n484), .ZN(new_n517));
  NOR3_X1   g316(.A1(new_n486), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n202), .B1(new_n478), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n443), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n476), .B1(new_n475), .B2(new_n449), .ZN(new_n521));
  AOI211_X1 g320(.A(KEYINPUT87), .B(new_n448), .C1(new_n473), .C2(new_n474), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n516), .A2(new_n517), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n485), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(KEYINPUT88), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT15), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT89), .B(G36gat), .ZN(new_n528));
  INV_X1    g327(.A(G29gat), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(G29gat), .A2(G36gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT14), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n527), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT14), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n531), .B(new_n534), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n535), .B(KEYINPUT15), .C1(new_n529), .C2(new_n528), .ZN(new_n536));
  XNOR2_X1  g335(.A(G43gat), .B(G50gat), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n533), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n530), .A2(new_n532), .ZN(new_n539));
  INV_X1    g338(.A(new_n537), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(KEYINPUT15), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(G8gat), .ZN(new_n543));
  XOR2_X1   g342(.A(G15gat), .B(G22gat), .Z(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(G1gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(G15gat), .B(G22gat), .ZN(new_n546));
  INV_X1    g345(.A(G1gat), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(KEYINPUT16), .A3(new_n547), .ZN(new_n548));
  AOI211_X1 g347(.A(KEYINPUT90), .B(new_n543), .C1(new_n545), .C2(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n543), .A2(KEYINPUT90), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n543), .A2(KEYINPUT90), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n545), .A2(new_n548), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n542), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT92), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n555), .A3(KEYINPUT92), .ZN(new_n559));
  NOR4_X1   g358(.A1(new_n530), .A2(new_n532), .A3(new_n527), .A4(new_n537), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n540), .B1(new_n539), .B2(KEYINPUT15), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n560), .B1(new_n561), .B2(new_n533), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n545), .A2(new_n548), .A3(new_n552), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n550), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n553), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT93), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  AND4_X1   g365(.A1(KEYINPUT93), .A2(new_n565), .A3(new_n538), .A4(new_n541), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n558), .B(new_n559), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n569), .B(KEYINPUT13), .Z(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT94), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n568), .A2(KEYINPUT94), .A3(new_n570), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT17), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n538), .A2(new_n576), .A3(new_n541), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n576), .B1(new_n538), .B2(new_n541), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n565), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n579), .A2(new_n569), .A3(new_n556), .ZN(new_n580));
  NOR2_X1   g379(.A1(KEYINPUT91), .A2(KEYINPUT18), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n579), .A2(new_n569), .A3(new_n556), .A4(new_n581), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n575), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G113gat), .B(G141gat), .ZN(new_n587));
  INV_X1    g386(.A(G197gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(KEYINPUT11), .B(G169gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT12), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n568), .A2(KEYINPUT94), .A3(new_n570), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT94), .B1(new_n568), .B2(new_n570), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n585), .B(new_n592), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n597), .A2(KEYINPUT95), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n597), .A2(KEYINPUT95), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n594), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AND3_X1   g399(.A1(new_n519), .A2(new_n526), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT96), .ZN(new_n603));
  XOR2_X1   g402(.A(G57gat), .B(G64gat), .Z(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G71gat), .B(G78gat), .Z(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(G64gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(G57gat), .ZN(new_n609));
  XOR2_X1   g408(.A(KEYINPUT97), .B(G57gat), .Z(new_n610));
  OAI21_X1  g409(.A(new_n609), .B1(new_n610), .B2(new_n608), .ZN(new_n611));
  INV_X1    g410(.A(new_n606), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(new_n612), .A3(new_n603), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT98), .B(KEYINPUT21), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT99), .ZN(new_n617));
  XOR2_X1   g416(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n603), .A2(new_n612), .ZN(new_n620));
  AOI22_X1  g419(.A1(new_n620), .A2(new_n611), .B1(new_n605), .B2(new_n606), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n555), .B1(KEYINPUT21), .B2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n619), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G127gat), .B(G155gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(G231gat), .A2(G233gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G183gat), .B(G211gat), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n628), .B(new_n629), .Z(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n625), .B(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT104), .ZN(new_n633));
  XNOR2_X1  g432(.A(G99gat), .B(G106gat), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT103), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G85gat), .A2(G92gat), .ZN(new_n637));
  NAND2_X1  g436(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n637), .B(new_n638), .Z(new_n639));
  NAND2_X1  g438(.A1(new_n634), .A2(new_n635), .ZN(new_n640));
  NAND2_X1  g439(.A1(G99gat), .A2(G106gat), .ZN(new_n641));
  INV_X1    g440(.A(G85gat), .ZN(new_n642));
  INV_X1    g441(.A(G92gat), .ZN(new_n643));
  AOI22_X1  g442(.A1(KEYINPUT8), .A2(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n636), .A2(new_n639), .A3(new_n640), .A4(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  AOI22_X1  g445(.A1(new_n640), .A2(new_n636), .B1(new_n639), .B2(new_n644), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n633), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n636), .A2(new_n640), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n639), .A2(new_n644), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n651), .A2(KEYINPUT104), .A3(new_n645), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(G232gat), .A2(G233gat), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  AOI22_X1  g454(.A1(new_n653), .A2(new_n542), .B1(KEYINPUT41), .B2(new_n655), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n648), .B(new_n652), .C1(new_n577), .C2(new_n578), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(G190gat), .B(G218gat), .Z(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n655), .A2(KEYINPUT41), .ZN(new_n661));
  XNOR2_X1  g460(.A(G134gat), .B(G162gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n659), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n656), .A2(new_n664), .A3(new_n657), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n660), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n663), .B1(new_n660), .B2(new_n665), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT106), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n607), .A2(KEYINPUT10), .A3(new_n613), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n671), .B1(new_n648), .B2(new_n652), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n650), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n674), .A2(new_n607), .A3(new_n613), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n675), .B1(new_n647), .B2(new_n646), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n621), .A2(new_n651), .A3(new_n645), .A4(new_n674), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT10), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n672), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(G230gat), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(new_n421), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n670), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n678), .A2(new_n681), .A3(new_n421), .ZN(new_n684));
  XNOR2_X1  g483(.A(G120gat), .B(G148gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(G176gat), .B(G204gat), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n685), .B(new_n686), .Z(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT10), .B1(new_n676), .B2(new_n677), .ZN(new_n690));
  OAI221_X1 g489(.A(KEYINPUT106), .B1(new_n681), .B2(new_n421), .C1(new_n690), .C2(new_n672), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n683), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n687), .B(KEYINPUT107), .Z(new_n693));
  NOR2_X1   g492(.A1(new_n680), .A2(new_n682), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n693), .B1(new_n694), .B2(new_n684), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n632), .A2(new_n669), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n601), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n398), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(new_n547), .ZN(G1324gat));
  INV_X1    g501(.A(new_n454), .ZN(new_n703));
  XOR2_X1   g502(.A(KEYINPUT16), .B(G8gat), .Z(new_n704));
  NAND4_X1  g503(.A1(new_n601), .A2(new_n703), .A3(new_n699), .A4(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT108), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(KEYINPUT42), .ZN(new_n707));
  OAI21_X1  g506(.A(G8gat), .B1(new_n700), .B2(new_n454), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n705), .A2(KEYINPUT108), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n707), .A2(new_n708), .A3(new_n710), .ZN(G1325gat));
  OAI21_X1  g510(.A(G15gat), .B1(new_n700), .B2(new_n481), .ZN(new_n712));
  INV_X1    g511(.A(new_n480), .ZN(new_n713));
  OR2_X1    g512(.A1(new_n713), .A2(G15gat), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n712), .B1(new_n700), .B2(new_n714), .ZN(G1326gat));
  NOR2_X1   g514(.A1(new_n700), .A2(new_n355), .ZN(new_n716));
  XOR2_X1   g515(.A(KEYINPUT43), .B(G22gat), .Z(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1327gat));
  NOR3_X1   g517(.A1(new_n632), .A2(new_n669), .A3(new_n696), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT109), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n519), .A2(new_n526), .A3(new_n600), .A4(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n722), .A2(new_n529), .A3(new_n399), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT45), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n669), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n519), .A2(new_n526), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n481), .A2(new_n484), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n516), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n668), .B1(new_n478), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n725), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n632), .A2(KEYINPUT110), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n625), .B(new_n630), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n597), .A2(KEYINPUT95), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT95), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n575), .A2(new_n739), .A3(new_n592), .A4(new_n585), .ZN(new_n740));
  AOI22_X1  g539(.A1(new_n738), .A2(new_n740), .B1(new_n593), .B2(new_n586), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n737), .A2(new_n741), .A3(new_n696), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT111), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n732), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(G29gat), .B1(new_n744), .B2(new_n398), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n724), .A2(new_n745), .ZN(G1328gat));
  INV_X1    g545(.A(new_n528), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n721), .A2(new_n454), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT46), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n744), .B2(new_n454), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(G1329gat));
  INV_X1    g550(.A(new_n481), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n727), .A2(new_n731), .A3(new_n752), .A4(new_n743), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G43gat), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n713), .A2(G43gat), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n722), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT47), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  AOI22_X1  g558(.A1(new_n753), .A2(G43gat), .B1(new_n722), .B2(new_n755), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT47), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n760), .A2(KEYINPUT112), .A3(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n759), .A2(new_n762), .ZN(G1330gat));
  INV_X1    g562(.A(KEYINPUT48), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n355), .A2(G50gat), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n764), .B1(new_n722), .B2(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n727), .A2(new_n731), .A3(new_n483), .A4(new_n743), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G50gat), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n766), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n769), .B1(new_n766), .B2(new_n768), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n772));
  INV_X1    g571(.A(new_n765), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n721), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n722), .A2(KEYINPUT113), .A3(new_n765), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n768), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  OAI22_X1  g575(.A1(new_n770), .A2(new_n771), .B1(new_n776), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g576(.A1(new_n478), .A2(new_n729), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT115), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n632), .A2(new_n741), .A3(new_n669), .A4(new_n696), .ZN(new_n780));
  OR3_X1    g579(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n778), .B2(new_n780), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n399), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(new_n610), .ZN(G1332gat));
  AOI21_X1  g585(.A(new_n454), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT116), .B1(new_n783), .B2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n781), .A2(new_n790), .A3(new_n782), .A4(new_n787), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT49), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n608), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n789), .A2(new_n793), .A3(new_n608), .A4(new_n791), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(G1333gat));
  OAI21_X1  g596(.A(G71gat), .B1(new_n783), .B2(new_n481), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n713), .A2(G71gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n781), .A2(new_n782), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n798), .A2(KEYINPUT50), .A3(new_n800), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(G1334gat));
  NAND2_X1  g604(.A1(new_n784), .A2(new_n483), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g606(.A1(new_n632), .A2(new_n600), .A3(new_n697), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n732), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(G85gat), .B1(new_n809), .B2(new_n398), .ZN(new_n810));
  INV_X1    g609(.A(new_n729), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n669), .B1(new_n523), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n632), .A2(new_n600), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(KEYINPUT51), .A3(new_n813), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n668), .B(new_n813), .C1(new_n478), .C2(new_n729), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT51), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n818), .A2(new_n642), .A3(new_n399), .A4(new_n696), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n810), .A2(new_n819), .ZN(G1336gat));
  NAND4_X1  g619(.A1(new_n727), .A2(new_n731), .A3(new_n703), .A4(new_n808), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(G92gat), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n454), .A2(G92gat), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n818), .A2(new_n696), .A3(new_n823), .ZN(new_n824));
  AOI211_X1 g623(.A(KEYINPUT117), .B(KEYINPUT52), .C1(new_n822), .C2(new_n824), .ZN(new_n825));
  OR2_X1    g624(.A1(KEYINPUT117), .A2(KEYINPUT52), .ZN(new_n826));
  NAND2_X1  g625(.A1(KEYINPUT117), .A2(KEYINPUT52), .ZN(new_n827));
  AND4_X1   g626(.A1(new_n826), .A2(new_n822), .A3(new_n824), .A4(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n825), .A2(new_n828), .ZN(G1337gat));
  OAI21_X1  g628(.A(G99gat), .B1(new_n809), .B2(new_n481), .ZN(new_n830));
  INV_X1    g629(.A(G99gat), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n713), .A2(new_n697), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n818), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n830), .A2(new_n833), .ZN(G1338gat));
  NAND4_X1  g633(.A1(new_n727), .A2(new_n731), .A3(new_n483), .A4(new_n808), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(G106gat), .ZN(new_n836));
  INV_X1    g635(.A(new_n818), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n697), .A2(G106gat), .A3(new_n355), .ZN(new_n838));
  XOR2_X1   g637(.A(new_n838), .B(KEYINPUT118), .Z(new_n839));
  OAI21_X1  g638(.A(new_n836), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT53), .ZN(new_n841));
  INV_X1    g640(.A(new_n838), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n842), .B1(new_n814), .B2(new_n817), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT53), .B1(new_n843), .B2(KEYINPUT119), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n844), .B(new_n836), .C1(KEYINPUT119), .C2(new_n843), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n841), .A2(new_n845), .ZN(G1339gat));
  NAND2_X1  g645(.A1(new_n699), .A2(new_n741), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n579), .A2(new_n556), .ZN(new_n848));
  OAI22_X1  g647(.A1(new_n848), .A2(new_n569), .B1(new_n568), .B2(new_n570), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n591), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n850), .B1(new_n598), .B2(new_n599), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n852), .B1(new_n680), .B2(new_n682), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n683), .A2(new_n853), .A3(new_n691), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n687), .B1(new_n694), .B2(new_n852), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT55), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n854), .A2(new_n855), .A3(KEYINPUT55), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n858), .A2(new_n668), .A3(new_n692), .A4(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n851), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n858), .A2(new_n692), .A3(new_n859), .ZN(new_n862));
  OAI22_X1  g661(.A1(new_n851), .A2(new_n697), .B1(new_n741), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n861), .B1(new_n863), .B2(new_n669), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n847), .B1(new_n864), .B2(new_n737), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n703), .A2(new_n398), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n356), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(G113gat), .B1(new_n869), .B2(new_n600), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n865), .A2(new_n355), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n480), .A3(new_n866), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n600), .A2(G113gat), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n870), .B1(new_n874), .B2(new_n875), .ZN(G1340gat));
  OAI21_X1  g675(.A(G120gat), .B1(new_n873), .B2(new_n697), .ZN(new_n877));
  OR3_X1    g676(.A1(new_n697), .A2(new_n216), .A3(new_n215), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n877), .B1(new_n868), .B2(new_n878), .ZN(G1341gat));
  INV_X1    g678(.A(new_n737), .ZN(new_n880));
  OAI22_X1  g679(.A1(new_n873), .A2(new_n880), .B1(new_n228), .B2(new_n227), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n632), .A2(new_n221), .A3(new_n223), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n868), .B2(new_n882), .ZN(G1342gat));
  NOR3_X1   g682(.A1(new_n868), .A2(G134gat), .A3(new_n669), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(KEYINPUT56), .ZN(new_n885));
  OAI21_X1  g684(.A(G134gat), .B1(new_n873), .B2(new_n669), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(G1343gat));
  AND2_X1   g686(.A1(new_n866), .A2(new_n481), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT57), .B1(new_n865), .B2(new_n483), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n355), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n858), .A2(new_n692), .A3(new_n859), .ZN(new_n893));
  AOI22_X1  g692(.A1(new_n738), .A2(new_n740), .B1(new_n591), .B2(new_n849), .ZN(new_n894));
  AOI22_X1  g693(.A1(new_n600), .A2(new_n893), .B1(new_n894), .B2(new_n696), .ZN(new_n895));
  OAI22_X1  g694(.A1(new_n895), .A2(new_n668), .B1(new_n851), .B2(new_n860), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n734), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n892), .B1(new_n897), .B2(new_n847), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n600), .B(new_n888), .C1(new_n889), .C2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n698), .A2(new_n600), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n902), .B1(new_n896), .B2(new_n880), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n890), .B1(new_n903), .B2(new_n355), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n864), .A2(new_n632), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n891), .B1(new_n905), .B2(new_n902), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n907), .A2(KEYINPUT120), .A3(new_n600), .A4(new_n888), .ZN(new_n908));
  INV_X1    g707(.A(new_n325), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n901), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n752), .A2(new_n355), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n867), .A2(new_n338), .A3(new_n600), .A4(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT58), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n909), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n912), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(KEYINPUT58), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n916), .A2(new_n919), .A3(KEYINPUT121), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n325), .B1(new_n899), .B2(new_n900), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n914), .B1(new_n922), .B2(new_n908), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n913), .B1(new_n917), .B2(new_n912), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n920), .A2(new_n925), .ZN(G1344gat));
  NAND2_X1  g725(.A1(new_n907), .A2(new_n888), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n927), .A2(new_n697), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n928), .A2(KEYINPUT59), .A3(new_n320), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT59), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n897), .A2(new_n847), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT57), .B1(new_n931), .B2(new_n483), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n903), .A2(new_n892), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n696), .B(new_n888), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n930), .B1(new_n934), .B2(G148gat), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n867), .A2(new_n911), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n696), .A2(new_n320), .ZN(new_n937));
  OAI22_X1  g736(.A1(new_n929), .A2(new_n935), .B1(new_n936), .B2(new_n937), .ZN(G1345gat));
  OAI21_X1  g737(.A(G155gat), .B1(new_n927), .B2(new_n880), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n734), .A2(G155gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n936), .B2(new_n940), .ZN(G1346gat));
  NOR3_X1   g740(.A1(new_n936), .A2(G162gat), .A3(new_n669), .ZN(new_n942));
  XOR2_X1   g741(.A(new_n942), .B(KEYINPUT122), .Z(new_n943));
  OAI21_X1  g742(.A(G162gat), .B1(new_n927), .B2(new_n669), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1347gat));
  NOR2_X1   g744(.A1(new_n454), .A2(new_n399), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n865), .A2(new_n356), .A3(new_n946), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n947), .A2(new_n261), .A3(new_n263), .A4(new_n600), .ZN(new_n948));
  XOR2_X1   g747(.A(new_n948), .B(KEYINPUT123), .Z(new_n949));
  NAND3_X1  g748(.A1(new_n872), .A2(new_n480), .A3(new_n946), .ZN(new_n950));
  OAI21_X1  g749(.A(G169gat), .B1(new_n950), .B2(new_n741), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(G1348gat));
  AOI21_X1  g751(.A(G176gat), .B1(new_n947), .B2(new_n696), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n832), .A2(G176gat), .A3(new_n946), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n872), .B2(new_n954), .ZN(G1349gat));
  NAND2_X1  g754(.A1(new_n234), .A2(G183gat), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n947), .A2(new_n956), .A3(new_n236), .A4(new_n632), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n950), .A2(new_n880), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n957), .B1(new_n958), .B2(new_n242), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g759(.A1(new_n947), .A2(new_n239), .A3(new_n668), .ZN(new_n961));
  OR2_X1    g760(.A1(new_n950), .A2(new_n669), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT124), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT61), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n962), .A2(new_n963), .A3(new_n964), .A4(G190gat), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n239), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n967));
  AOI22_X1  g766(.A1(new_n962), .A2(new_n967), .B1(new_n963), .B2(new_n964), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n961), .B1(new_n966), .B2(new_n968), .ZN(G1351gat));
  NAND2_X1  g768(.A1(new_n481), .A2(new_n946), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n865), .A2(new_n483), .A3(new_n971), .ZN(new_n972));
  XOR2_X1   g771(.A(new_n972), .B(KEYINPUT125), .Z(new_n973));
  AOI21_X1  g772(.A(G197gat), .B1(new_n973), .B2(new_n600), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n932), .A2(new_n933), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(KEYINPUT126), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n977), .B1(new_n932), .B2(new_n933), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n970), .A2(new_n588), .A3(new_n741), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n974), .B1(new_n979), .B2(new_n980), .ZN(G1352gat));
  NOR3_X1   g780(.A1(new_n972), .A2(G204gat), .A3(new_n697), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n982), .B(KEYINPUT62), .ZN(new_n983));
  AOI211_X1 g782(.A(new_n697), .B(new_n970), .C1(new_n976), .C2(new_n978), .ZN(new_n984));
  INV_X1    g783(.A(G204gat), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(G1353gat));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n632), .ZN(new_n987));
  OAI21_X1  g786(.A(G211gat), .B1(new_n975), .B2(new_n987), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT63), .ZN(new_n989));
  XNOR2_X1  g788(.A(new_n988), .B(new_n989), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n973), .A2(new_n307), .A3(new_n632), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(G1354gat));
  AOI21_X1  g791(.A(G218gat), .B1(new_n973), .B2(new_n668), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n668), .A2(G218gat), .ZN(new_n994));
  XOR2_X1   g793(.A(new_n994), .B(KEYINPUT127), .Z(new_n995));
  NOR2_X1   g794(.A1(new_n995), .A2(new_n970), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n993), .B1(new_n979), .B2(new_n996), .ZN(G1355gat));
endmodule


