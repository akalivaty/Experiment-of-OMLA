

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757;

  XNOR2_X1 U373 ( .A(n378), .B(G113), .ZN(n538) );
  XOR2_X1 U374 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n351) );
  NOR2_X2 U375 ( .A1(n427), .A2(n425), .ZN(n424) );
  AND2_X1 U376 ( .A1(n561), .A2(n560), .ZN(n547) );
  OR2_X2 U377 ( .A1(n742), .A2(KEYINPUT2), .ZN(n634) );
  OR2_X2 U378 ( .A1(n479), .A2(G902), .ZN(n437) );
  XNOR2_X2 U379 ( .A(n611), .B(KEYINPUT35), .ZN(n750) );
  XNOR2_X2 U380 ( .A(n521), .B(n520), .ZN(n376) );
  NOR2_X1 U381 ( .A1(n616), .A2(n637), .ZN(n609) );
  NOR2_X1 U382 ( .A1(n554), .A2(n568), .ZN(n555) );
  INV_X2 U383 ( .A(G953), .ZN(n490) );
  AND2_X1 U384 ( .A1(n634), .A2(n635), .ZN(n625) );
  XNOR2_X1 U385 ( .A(n352), .B(KEYINPUT82), .ZN(n742) );
  XNOR2_X1 U386 ( .A(n555), .B(n388), .ZN(n756) );
  XNOR2_X1 U387 ( .A(n560), .B(KEYINPUT102), .ZN(n544) );
  NOR2_X1 U388 ( .A1(n674), .A2(G953), .ZN(n677) );
  OR2_X1 U389 ( .A1(n734), .A2(KEYINPUT2), .ZN(n635) );
  AND2_X1 U390 ( .A1(n463), .A2(n467), .ZN(n390) );
  XNOR2_X1 U391 ( .A(n391), .B(n361), .ZN(n368) );
  NAND2_X1 U392 ( .A1(n451), .A2(n452), .ZN(n616) );
  NAND2_X1 U393 ( .A1(n453), .A2(n452), .ZN(n391) );
  AND2_X1 U394 ( .A1(n461), .A2(n454), .ZN(n453) );
  NAND2_X1 U395 ( .A1(n458), .A2(n456), .ZN(n452) );
  AND2_X1 U396 ( .A1(n558), .A2(n522), .ZN(n523) );
  XNOR2_X1 U397 ( .A(n643), .B(KEYINPUT80), .ZN(n619) );
  NAND2_X1 U398 ( .A1(n701), .A2(n626), .ZN(n521) );
  INV_X1 U399 ( .A(n544), .ZN(n545) );
  XNOR2_X1 U400 ( .A(n533), .B(G478), .ZN(n561) );
  XNOR2_X1 U401 ( .A(n505), .B(n355), .ZN(n653) );
  XNOR2_X1 U402 ( .A(n719), .B(n718), .ZN(n720) );
  XNOR2_X1 U403 ( .A(n529), .B(n396), .ZN(n719) );
  XNOR2_X1 U404 ( .A(n406), .B(n514), .ZN(n516) );
  XNOR2_X1 U405 ( .A(n537), .B(n534), .ZN(n431) );
  XNOR2_X1 U406 ( .A(n414), .B(G131), .ZN(n534) );
  XNOR2_X1 U407 ( .A(n386), .B(G146), .ZN(n515) );
  XNOR2_X1 U408 ( .A(G134), .B(G137), .ZN(n405) );
  NOR2_X1 U409 ( .A1(n587), .A2(n380), .ZN(n352) );
  XNOR2_X2 U410 ( .A(n740), .B(G146), .ZN(n379) );
  XNOR2_X2 U411 ( .A(n393), .B(n517), .ZN(n740) );
  AND2_X1 U412 ( .A1(n756), .A2(n557), .ZN(n419) );
  XNOR2_X1 U413 ( .A(n515), .B(n356), .ZN(n406) );
  XNOR2_X1 U414 ( .A(n434), .B(KEYINPUT71), .ZN(n571) );
  NAND2_X1 U415 ( .A1(n619), .A2(n435), .ZN(n434) );
  INV_X1 U416 ( .A(KEYINPUT47), .ZN(n435) );
  XNOR2_X1 U417 ( .A(G113), .B(G116), .ZN(n470) );
  XNOR2_X1 U418 ( .A(KEYINPUT67), .B(KEYINPUT48), .ZN(n581) );
  NOR2_X1 U419 ( .A1(n417), .A2(n415), .ZN(n582) );
  AND2_X1 U420 ( .A1(n467), .A2(n612), .ZN(n464) );
  NAND2_X1 U421 ( .A1(n390), .A2(n374), .ZN(n372) );
  AND2_X1 U422 ( .A1(n407), .A2(n621), .ZN(n374) );
  NOR2_X1 U423 ( .A1(n750), .A2(n612), .ZN(n407) );
  XNOR2_X1 U424 ( .A(G110), .B(KEYINPUT16), .ZN(n508) );
  INV_X1 U425 ( .A(KEYINPUT69), .ZN(n450) );
  XNOR2_X1 U426 ( .A(n377), .B(G119), .ZN(n509) );
  XNOR2_X1 U427 ( .A(G101), .B(KEYINPUT3), .ZN(n377) );
  XNOR2_X1 U428 ( .A(n413), .B(n534), .ZN(n393) );
  XNOR2_X1 U429 ( .A(n405), .B(n404), .ZN(n413) );
  INV_X1 U430 ( .A(KEYINPUT66), .ZN(n404) );
  NAND2_X1 U431 ( .A1(n653), .A2(n550), .ZN(n573) );
  INV_X1 U432 ( .A(n549), .ZN(n383) );
  INV_X1 U433 ( .A(KEYINPUT86), .ZN(n566) );
  XNOR2_X1 U434 ( .A(n448), .B(G107), .ZN(n527) );
  INV_X1 U435 ( .A(G116), .ZN(n448) );
  XNOR2_X1 U436 ( .A(n525), .B(n412), .ZN(n411) );
  INV_X1 U437 ( .A(KEYINPUT7), .ZN(n412) );
  XOR2_X1 U438 ( .A(KEYINPUT9), .B(KEYINPUT103), .Z(n525) );
  XNOR2_X1 U439 ( .A(G104), .B(G101), .ZN(n487) );
  XOR2_X1 U440 ( .A(G140), .B(G107), .Z(n488) );
  NAND2_X1 U441 ( .A1(n439), .A2(n387), .ZN(n701) );
  NAND2_X1 U442 ( .A1(n444), .A2(n443), .ZN(n387) );
  XNOR2_X1 U443 ( .A(n635), .B(n398), .ZN(n397) );
  INV_X1 U444 ( .A(KEYINPUT81), .ZN(n398) );
  INV_X1 U445 ( .A(G469), .ZN(n423) );
  NOR2_X1 U446 ( .A1(G902), .A2(n709), .ZN(n494) );
  INV_X1 U447 ( .A(n653), .ZN(n601) );
  XNOR2_X1 U448 ( .A(n572), .B(n426), .ZN(n425) );
  INV_X1 U449 ( .A(KEYINPUT70), .ZN(n426) );
  INV_X1 U450 ( .A(KEYINPUT4), .ZN(n392) );
  NAND2_X1 U451 ( .A1(G234), .A2(G237), .ZN(n481) );
  INV_X1 U452 ( .A(G125), .ZN(n386) );
  NOR2_X2 U453 ( .A1(G953), .A2(G237), .ZN(n535) );
  NAND2_X1 U454 ( .A1(n588), .A2(n375), .ZN(n381) );
  NOR2_X1 U455 ( .A1(G237), .A2(G902), .ZN(n477) );
  INV_X1 U456 ( .A(n573), .ZN(n389) );
  XNOR2_X1 U457 ( .A(n502), .B(n402), .ZN(n506) );
  XNOR2_X1 U458 ( .A(n503), .B(KEYINPUT96), .ZN(n402) );
  XOR2_X1 U459 ( .A(KEYINPUT97), .B(KEYINPUT20), .Z(n503) );
  NAND2_X1 U460 ( .A1(n460), .A2(KEYINPUT0), .ZN(n459) );
  INV_X1 U461 ( .A(n596), .ZN(n460) );
  AND2_X1 U462 ( .A1(n596), .A2(n457), .ZN(n456) );
  INV_X1 U463 ( .A(KEYINPUT0), .ZN(n457) );
  XNOR2_X1 U464 ( .A(n379), .B(n438), .ZN(n479) );
  NAND2_X1 U465 ( .A1(n375), .A2(n699), .ZN(n380) );
  INV_X1 U466 ( .A(KEYINPUT45), .ZN(n369) );
  NAND2_X1 U467 ( .A1(n372), .A2(n371), .ZN(n370) );
  NAND2_X1 U468 ( .A1(n466), .A2(n373), .ZN(n371) );
  XNOR2_X1 U469 ( .A(n510), .B(n511), .ZN(n728) );
  XNOR2_X1 U470 ( .A(n449), .B(n527), .ZN(n511) );
  XNOR2_X1 U471 ( .A(n508), .B(n450), .ZN(n449) );
  INV_X1 U472 ( .A(KEYINPUT65), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n429), .B(n515), .ZN(n739) );
  XNOR2_X1 U474 ( .A(n367), .B(n366), .ZN(n429) );
  INV_X1 U475 ( .A(G140), .ZN(n366) );
  XNOR2_X1 U476 ( .A(KEYINPUT64), .B(KEYINPUT10), .ZN(n367) );
  OR2_X2 U477 ( .A1(n694), .A2(n573), .ZN(n399) );
  XNOR2_X1 U478 ( .A(n385), .B(n384), .ZN(n558) );
  INV_X1 U479 ( .A(KEYINPUT76), .ZN(n384) );
  AND2_X1 U480 ( .A1(n601), .A2(n360), .ZN(n382) );
  XNOR2_X1 U481 ( .A(n480), .B(KEYINPUT30), .ZN(n559) );
  NOR2_X1 U482 ( .A1(n640), .A2(n615), .ZN(n480) );
  AND2_X1 U483 ( .A1(n601), .A2(n597), .ZN(n649) );
  XNOR2_X1 U484 ( .A(n479), .B(KEYINPUT62), .ZN(n629) );
  XNOR2_X1 U485 ( .A(n532), .B(n528), .ZN(n396) );
  XNOR2_X1 U486 ( .A(n526), .B(n411), .ZN(n529) );
  XNOR2_X1 U487 ( .A(n379), .B(n493), .ZN(n709) );
  XNOR2_X1 U488 ( .A(n701), .B(n363), .ZN(n702) );
  NOR2_X1 U489 ( .A1(G952), .A2(n490), .ZN(n727) );
  AND2_X1 U490 ( .A1(n638), .A2(n359), .ZN(n672) );
  INV_X1 U491 ( .A(KEYINPUT42), .ZN(n388) );
  NAND2_X1 U492 ( .A1(n546), .A2(n691), .ZN(n436) );
  INV_X1 U493 ( .A(n605), .ZN(n395) );
  XNOR2_X1 U494 ( .A(n408), .B(n548), .ZN(n663) );
  INV_X1 U495 ( .A(n467), .ZN(n465) );
  NAND2_X1 U496 ( .A1(n395), .A2(n358), .ZN(n467) );
  AND2_X1 U497 ( .A1(n690), .A2(n570), .ZN(n353) );
  AND2_X1 U498 ( .A1(n577), .A2(n649), .ZN(n354) );
  XOR2_X1 U499 ( .A(n504), .B(KEYINPUT25), .Z(n355) );
  INV_X1 U500 ( .A(n375), .ZN(n700) );
  AND2_X1 U501 ( .A1(G224), .A2(n490), .ZN(n356) );
  AND2_X1 U502 ( .A1(n648), .A2(n663), .ZN(n357) );
  AND2_X1 U503 ( .A1(n601), .A2(n607), .ZN(n358) );
  NOR2_X1 U504 ( .A1(n671), .A2(n357), .ZN(n359) );
  AND2_X1 U505 ( .A1(n597), .A2(n383), .ZN(n360) );
  XOR2_X1 U506 ( .A(KEYINPUT68), .B(KEYINPUT22), .Z(n361) );
  XOR2_X1 U507 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n362) );
  XNOR2_X1 U508 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n363) );
  XOR2_X1 U509 ( .A(n708), .B(n707), .Z(n364) );
  INV_X1 U510 ( .A(n739), .ZN(n428) );
  XNOR2_X2 U511 ( .A(n365), .B(n541), .ZN(n560) );
  NOR2_X2 U512 ( .A1(n714), .A2(G902), .ZN(n365) );
  NAND2_X1 U513 ( .A1(n368), .A2(n599), .ZN(n605) );
  NAND2_X1 U514 ( .A1(n368), .A2(n603), .ZN(n604) );
  XNOR2_X2 U515 ( .A(n370), .B(n369), .ZN(n734) );
  AND2_X1 U516 ( .A1(n464), .A2(n621), .ZN(n373) );
  NAND2_X1 U517 ( .A1(n376), .A2(n565), .ZN(n567) );
  XNOR2_X1 U518 ( .A(n376), .B(KEYINPUT38), .ZN(n639) );
  NAND2_X1 U519 ( .A1(n564), .A2(n376), .ZN(n690) );
  OR2_X1 U520 ( .A1(n586), .A2(n376), .ZN(n375) );
  XNOR2_X1 U521 ( .A(n538), .B(n509), .ZN(n510) );
  XNOR2_X2 U522 ( .A(G104), .B(G122), .ZN(n378) );
  OR2_X2 U523 ( .A1(n587), .A2(n381), .ZN(n589) );
  NAND2_X1 U524 ( .A1(n577), .A2(n382), .ZN(n385) );
  XNOR2_X2 U525 ( .A(n494), .B(n423), .ZN(n577) );
  NAND2_X1 U526 ( .A1(n723), .A2(G472), .ZN(n628) );
  NOR2_X4 U527 ( .A1(n627), .A2(n626), .ZN(n723) );
  XNOR2_X1 U528 ( .A(n628), .B(n629), .ZN(n630) );
  INV_X1 U529 ( .A(n657), .ZN(n615) );
  AND2_X1 U530 ( .A1(n657), .A2(n389), .ZN(n552) );
  XNOR2_X2 U531 ( .A(n437), .B(G472), .ZN(n657) );
  NOR2_X1 U532 ( .A1(n725), .A2(G902), .ZN(n505) );
  XNOR2_X2 U533 ( .A(n530), .B(n392), .ZN(n517) );
  XNOR2_X1 U534 ( .A(n394), .B(n500), .ZN(n501) );
  XNOR2_X1 U535 ( .A(n498), .B(n401), .ZN(n394) );
  XNOR2_X1 U536 ( .A(n579), .B(KEYINPUT109), .ZN(n751) );
  NOR2_X2 U537 ( .A1(n607), .A2(n399), .ZN(n583) );
  NAND2_X1 U538 ( .A1(n622), .A2(n734), .ZN(n624) );
  NOR2_X2 U539 ( .A1(n568), .A2(n590), .ZN(n692) );
  NAND2_X1 U540 ( .A1(n553), .A2(n577), .ZN(n568) );
  NAND2_X1 U541 ( .A1(n636), .A2(n397), .ZN(n638) );
  XNOR2_X2 U542 ( .A(KEYINPUT1), .B(n577), .ZN(n650) );
  XOR2_X2 U543 ( .A(G143), .B(G128), .Z(n530) );
  XNOR2_X2 U544 ( .A(n400), .B(KEYINPUT39), .ZN(n546) );
  NAND2_X1 U545 ( .A1(n523), .A2(n559), .ZN(n400) );
  XNOR2_X1 U546 ( .A(n497), .B(n351), .ZN(n401) );
  NAND2_X1 U547 ( .A1(n422), .A2(n421), .ZN(n420) );
  XNOR2_X2 U548 ( .A(G902), .B(KEYINPUT15), .ZN(n626) );
  NAND2_X1 U549 ( .A1(n403), .A2(n610), .ZN(n611) );
  XNOR2_X1 U550 ( .A(n609), .B(KEYINPUT34), .ZN(n403) );
  NOR2_X2 U551 ( .A1(n704), .A2(n727), .ZN(n706) );
  NAND2_X1 U552 ( .A1(n580), .A2(n353), .ZN(n427) );
  NAND2_X1 U553 ( .A1(n644), .A2(n641), .ZN(n408) );
  XNOR2_X1 U554 ( .A(n409), .B(KEYINPUT122), .ZN(G63) );
  NOR2_X2 U555 ( .A1(n722), .A2(n727), .ZN(n409) );
  XNOR2_X1 U556 ( .A(n410), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U557 ( .A1(n717), .A2(n727), .ZN(n410) );
  NAND2_X1 U558 ( .A1(n424), .A2(n416), .ZN(n415) );
  OR2_X1 U559 ( .A1(n756), .A2(n557), .ZN(n416) );
  NAND2_X1 U560 ( .A1(n420), .A2(n418), .ZN(n417) );
  NAND2_X1 U561 ( .A1(n755), .A2(n419), .ZN(n418) );
  INV_X1 U562 ( .A(n557), .ZN(n421) );
  INV_X1 U563 ( .A(n755), .ZN(n422) );
  XNOR2_X2 U564 ( .A(n436), .B(n362), .ZN(n755) );
  XNOR2_X2 U565 ( .A(n430), .B(n428), .ZN(n714) );
  XNOR2_X2 U566 ( .A(n432), .B(n431), .ZN(n430) );
  XNOR2_X2 U567 ( .A(n539), .B(n433), .ZN(n432) );
  XNOR2_X2 U568 ( .A(n536), .B(KEYINPUT12), .ZN(n433) );
  XNOR2_X1 U569 ( .A(n476), .B(n472), .ZN(n438) );
  NAND2_X1 U570 ( .A1(n446), .A2(n728), .ZN(n439) );
  NAND2_X1 U571 ( .A1(n440), .A2(n445), .ZN(n444) );
  NAND2_X1 U572 ( .A1(n447), .A2(n518), .ZN(n440) );
  INV_X1 U573 ( .A(n516), .ZN(n447) );
  NAND2_X1 U574 ( .A1(n516), .A2(n517), .ZN(n445) );
  NAND2_X1 U575 ( .A1(n442), .A2(n441), .ZN(n446) );
  NAND2_X1 U576 ( .A1(n447), .A2(n517), .ZN(n441) );
  NAND2_X1 U577 ( .A1(n516), .A2(n518), .ZN(n442) );
  INV_X1 U578 ( .A(n728), .ZN(n443) );
  NAND2_X1 U579 ( .A1(n590), .A2(KEYINPUT0), .ZN(n461) );
  AND2_X1 U580 ( .A1(n461), .A2(n459), .ZN(n451) );
  NOR2_X1 U581 ( .A1(n598), .A2(n455), .ZN(n454) );
  INV_X1 U582 ( .A(n459), .ZN(n455) );
  INV_X1 U583 ( .A(n590), .ZN(n458) );
  NAND2_X1 U584 ( .A1(n462), .A2(n468), .ZN(n466) );
  AND2_X1 U585 ( .A1(n685), .A2(n754), .ZN(n462) );
  AND2_X1 U586 ( .A1(n685), .A2(n754), .ZN(n463) );
  INV_X1 U587 ( .A(n750), .ZN(n468) );
  XNOR2_X2 U588 ( .A(n624), .B(n623), .ZN(n633) );
  NOR2_X2 U589 ( .A1(n630), .A2(n727), .ZN(n632) );
  XNOR2_X1 U590 ( .A(n716), .B(n715), .ZN(n717) );
  XNOR2_X1 U591 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U592 ( .A(n709), .B(n364), .ZN(n710) );
  AND2_X1 U593 ( .A1(n615), .A2(n653), .ZN(n469) );
  XNOR2_X1 U594 ( .A(n556), .B(KEYINPUT84), .ZN(n557) );
  INV_X1 U595 ( .A(KEYINPUT44), .ZN(n612) );
  INV_X1 U596 ( .A(KEYINPUT75), .ZN(n623) );
  XNOR2_X1 U597 ( .A(KEYINPUT41), .B(KEYINPUT108), .ZN(n548) );
  XNOR2_X1 U598 ( .A(n475), .B(n509), .ZN(n476) );
  XNOR2_X1 U599 ( .A(n531), .B(G134), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n540), .B(G475), .ZN(n541) );
  INV_X1 U601 ( .A(KEYINPUT121), .ZN(n718) );
  XNOR2_X1 U602 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U603 ( .A(KEYINPUT63), .B(KEYINPUT87), .ZN(n631) );
  XNOR2_X1 U604 ( .A(n677), .B(n676), .ZN(G75) );
  XOR2_X1 U605 ( .A(KEYINPUT5), .B(KEYINPUT99), .Z(n471) );
  XNOR2_X1 U606 ( .A(n471), .B(n470), .ZN(n472) );
  XOR2_X1 U607 ( .A(KEYINPUT74), .B(KEYINPUT98), .Z(n474) );
  NAND2_X1 U608 ( .A1(n535), .A2(G210), .ZN(n473) );
  XNOR2_X1 U609 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U610 ( .A(n477), .B(KEYINPUT73), .ZN(n519) );
  NAND2_X1 U611 ( .A1(n519), .A2(G214), .ZN(n478) );
  XOR2_X1 U612 ( .A(KEYINPUT90), .B(n478), .Z(n640) );
  XOR2_X1 U613 ( .A(KEYINPUT91), .B(KEYINPUT14), .Z(n482) );
  XNOR2_X1 U614 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U615 ( .A(KEYINPUT72), .B(n483), .ZN(n484) );
  NAND2_X1 U616 ( .A1(G952), .A2(n484), .ZN(n670) );
  NOR2_X1 U617 ( .A1(G953), .A2(n670), .ZN(n594) );
  AND2_X1 U618 ( .A1(n484), .A2(G953), .ZN(n485) );
  NAND2_X1 U619 ( .A1(G902), .A2(n485), .ZN(n591) );
  NOR2_X1 U620 ( .A1(G900), .A2(n591), .ZN(n486) );
  NOR2_X1 U621 ( .A1(n594), .A2(n486), .ZN(n549) );
  XNOR2_X1 U622 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U623 ( .A(G110), .B(n489), .Z(n492) );
  NAND2_X1 U624 ( .A1(G227), .A2(n490), .ZN(n491) );
  XNOR2_X1 U625 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U626 ( .A(G137), .B(G128), .Z(n496) );
  XNOR2_X1 U627 ( .A(G119), .B(G110), .ZN(n495) );
  XNOR2_X1 U628 ( .A(n496), .B(n495), .ZN(n498) );
  XOR2_X1 U629 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n497) );
  NAND2_X1 U630 ( .A1(n490), .A2(G234), .ZN(n499) );
  XOR2_X1 U631 ( .A(KEYINPUT8), .B(n499), .Z(n524) );
  NAND2_X1 U632 ( .A1(G221), .A2(n524), .ZN(n500) );
  XNOR2_X1 U633 ( .A(n501), .B(n739), .ZN(n725) );
  NAND2_X1 U634 ( .A1(G234), .A2(n626), .ZN(n502) );
  NAND2_X1 U635 ( .A1(G217), .A2(n506), .ZN(n504) );
  NAND2_X1 U636 ( .A1(n506), .A2(G221), .ZN(n507) );
  XOR2_X1 U637 ( .A(KEYINPUT21), .B(n507), .Z(n597) );
  INV_X1 U638 ( .A(n597), .ZN(n652) );
  XOR2_X1 U639 ( .A(KEYINPUT77), .B(KEYINPUT89), .Z(n513) );
  XNOR2_X1 U640 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n512) );
  XNOR2_X1 U641 ( .A(n513), .B(n512), .ZN(n514) );
  INV_X1 U642 ( .A(n517), .ZN(n518) );
  AND2_X1 U643 ( .A1(G210), .A2(n519), .ZN(n520) );
  INV_X1 U644 ( .A(n639), .ZN(n522) );
  NAND2_X1 U645 ( .A1(G217), .A2(n524), .ZN(n526) );
  XNOR2_X1 U646 ( .A(G122), .B(n527), .ZN(n528) );
  INV_X1 U647 ( .A(n530), .ZN(n531) );
  NOR2_X1 U648 ( .A1(n719), .A2(G902), .ZN(n533) );
  INV_X1 U649 ( .A(n561), .ZN(n542) );
  XOR2_X1 U650 ( .A(G143), .B(KEYINPUT11), .Z(n537) );
  NAND2_X1 U651 ( .A1(n535), .A2(G214), .ZN(n536) );
  INV_X1 U652 ( .A(n538), .ZN(n539) );
  XNOR2_X1 U653 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n540) );
  NAND2_X1 U654 ( .A1(n542), .A2(n544), .ZN(n696) );
  INV_X1 U655 ( .A(n696), .ZN(n686) );
  NAND2_X1 U656 ( .A1(n546), .A2(n686), .ZN(n699) );
  NAND2_X1 U657 ( .A1(KEYINPUT2), .A2(n699), .ZN(n543) );
  XNOR2_X1 U658 ( .A(KEYINPUT79), .B(n543), .ZN(n588) );
  NAND2_X2 U659 ( .A1(n545), .A2(n561), .ZN(n694) );
  INV_X1 U660 ( .A(n694), .ZN(n691) );
  XNOR2_X1 U661 ( .A(n547), .B(KEYINPUT104), .ZN(n641) );
  NOR2_X1 U662 ( .A1(n639), .A2(n640), .ZN(n644) );
  INV_X1 U663 ( .A(n663), .ZN(n554) );
  NOR2_X1 U664 ( .A1(n549), .A2(n652), .ZN(n550) );
  XNOR2_X1 U665 ( .A(KEYINPUT106), .B(KEYINPUT28), .ZN(n551) );
  XNOR2_X1 U666 ( .A(n552), .B(n551), .ZN(n553) );
  INV_X1 U667 ( .A(KEYINPUT46), .ZN(n556) );
  NAND2_X1 U668 ( .A1(n559), .A2(n558), .ZN(n563) );
  NOR2_X1 U669 ( .A1(n561), .A2(n560), .ZN(n610) );
  INV_X1 U670 ( .A(n610), .ZN(n562) );
  NOR2_X1 U671 ( .A1(n563), .A2(n562), .ZN(n564) );
  INV_X1 U672 ( .A(n640), .ZN(n565) );
  XNOR2_X2 U673 ( .A(n567), .B(n566), .ZN(n574) );
  XNOR2_X2 U674 ( .A(n574), .B(KEYINPUT19), .ZN(n590) );
  NAND2_X1 U675 ( .A1(n696), .A2(n694), .ZN(n643) );
  NAND2_X1 U676 ( .A1(n692), .A2(n643), .ZN(n569) );
  NAND2_X1 U677 ( .A1(KEYINPUT47), .A2(n569), .ZN(n570) );
  NAND2_X1 U678 ( .A1(n571), .A2(n692), .ZN(n572) );
  XNOR2_X1 U679 ( .A(n657), .B(KEYINPUT6), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n583), .A2(n574), .ZN(n576) );
  XNOR2_X1 U681 ( .A(KEYINPUT36), .B(KEYINPUT85), .ZN(n575) );
  XNOR2_X1 U682 ( .A(n576), .B(n575), .ZN(n578) );
  NAND2_X1 U683 ( .A1(n578), .A2(n650), .ZN(n579) );
  INV_X1 U684 ( .A(n751), .ZN(n580) );
  XNOR2_X1 U685 ( .A(n582), .B(n581), .ZN(n587) );
  INV_X1 U686 ( .A(n650), .ZN(n599) );
  NAND2_X1 U687 ( .A1(n599), .A2(n583), .ZN(n584) );
  NOR2_X1 U688 ( .A1(n640), .A2(n584), .ZN(n585) );
  XNOR2_X1 U689 ( .A(n585), .B(KEYINPUT43), .ZN(n586) );
  XNOR2_X1 U690 ( .A(n589), .B(KEYINPUT83), .ZN(n622) );
  NOR2_X1 U691 ( .A1(G898), .A2(n591), .ZN(n592) );
  XNOR2_X1 U692 ( .A(n592), .B(KEYINPUT92), .ZN(n593) );
  NOR2_X1 U693 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U694 ( .A(KEYINPUT93), .B(n595), .ZN(n596) );
  NAND2_X1 U695 ( .A1(n641), .A2(n597), .ZN(n598) );
  NAND2_X1 U696 ( .A1(n650), .A2(n607), .ZN(n600) );
  NOR2_X1 U697 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U698 ( .A(KEYINPUT78), .B(n602), .ZN(n603) );
  XNOR2_X1 U699 ( .A(KEYINPUT32), .B(n604), .ZN(n754) );
  XNOR2_X1 U700 ( .A(n605), .B(KEYINPUT105), .ZN(n606) );
  NAND2_X1 U701 ( .A1(n606), .A2(n469), .ZN(n685) );
  NAND2_X1 U702 ( .A1(n649), .A2(n650), .ZN(n614) );
  NOR2_X1 U703 ( .A1(n614), .A2(n607), .ZN(n608) );
  XNOR2_X1 U704 ( .A(n608), .B(KEYINPUT33), .ZN(n637) );
  NOR2_X1 U705 ( .A1(n657), .A2(n616), .ZN(n613) );
  NAND2_X1 U706 ( .A1(n354), .A2(n613), .ZN(n680) );
  OR2_X1 U707 ( .A1(n615), .A2(n614), .ZN(n660) );
  NOR2_X1 U708 ( .A1(n616), .A2(n660), .ZN(n618) );
  XNOR2_X1 U709 ( .A(KEYINPUT100), .B(KEYINPUT31), .ZN(n617) );
  XNOR2_X1 U710 ( .A(n618), .B(n617), .ZN(n697) );
  NAND2_X1 U711 ( .A1(n680), .A2(n697), .ZN(n620) );
  NAND2_X1 U712 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U713 ( .A1(n633), .A2(n625), .ZN(n627) );
  XNOR2_X1 U714 ( .A(n632), .B(n631), .ZN(G57) );
  INV_X1 U715 ( .A(KEYINPUT116), .ZN(n673) );
  AND2_X1 U716 ( .A1(n633), .A2(n634), .ZN(n636) );
  INV_X1 U717 ( .A(n637), .ZN(n648) );
  XNOR2_X1 U718 ( .A(KEYINPUT115), .B(KEYINPUT52), .ZN(n668) );
  NAND2_X1 U719 ( .A1(n640), .A2(n639), .ZN(n642) );
  NAND2_X1 U720 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U721 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U722 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U723 ( .A1(n648), .A2(n647), .ZN(n666) );
  OR2_X1 U724 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U725 ( .A(n651), .B(KEYINPUT50), .ZN(n659) );
  XOR2_X1 U726 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n655) );
  NAND2_X1 U727 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U728 ( .A(n655), .B(n654), .Z(n656) );
  NOR2_X1 U729 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U730 ( .A1(n659), .A2(n658), .ZN(n661) );
  NAND2_X1 U731 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U732 ( .A(KEYINPUT51), .B(n662), .Z(n664) );
  NAND2_X1 U733 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U734 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U735 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X1 U736 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U737 ( .A(n673), .B(n672), .ZN(n674) );
  INV_X1 U738 ( .A(KEYINPUT117), .ZN(n675) );
  XNOR2_X1 U739 ( .A(n675), .B(KEYINPUT53), .ZN(n676) );
  XOR2_X1 U740 ( .A(G101), .B(n465), .Z(G3) );
  NOR2_X1 U741 ( .A1(n694), .A2(n680), .ZN(n678) );
  XOR2_X1 U742 ( .A(KEYINPUT110), .B(n678), .Z(n679) );
  XNOR2_X1 U743 ( .A(G104), .B(n679), .ZN(G6) );
  NOR2_X1 U744 ( .A1(n680), .A2(n696), .ZN(n684) );
  XOR2_X1 U745 ( .A(KEYINPUT111), .B(KEYINPUT26), .Z(n682) );
  XNOR2_X1 U746 ( .A(G107), .B(KEYINPUT27), .ZN(n681) );
  XNOR2_X1 U747 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U748 ( .A(n684), .B(n683), .ZN(G9) );
  XNOR2_X1 U749 ( .A(n685), .B(G110), .ZN(G12) );
  XOR2_X1 U750 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n688) );
  NAND2_X1 U751 ( .A1(n692), .A2(n686), .ZN(n687) );
  XNOR2_X1 U752 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U753 ( .A(G128), .B(n689), .ZN(G30) );
  XNOR2_X1 U754 ( .A(G143), .B(n690), .ZN(G45) );
  NAND2_X1 U755 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U756 ( .A(n693), .B(G146), .ZN(G48) );
  NOR2_X1 U757 ( .A1(n697), .A2(n694), .ZN(n695) );
  XOR2_X1 U758 ( .A(G113), .B(n695), .Z(G15) );
  NOR2_X1 U759 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U760 ( .A(G116), .B(n698), .Z(G18) );
  XNOR2_X1 U761 ( .A(G134), .B(n699), .ZN(G36) );
  XOR2_X1 U762 ( .A(G140), .B(n700), .Z(G42) );
  NAND2_X1 U763 ( .A1(n723), .A2(G210), .ZN(n703) );
  XNOR2_X1 U764 ( .A(KEYINPUT56), .B(KEYINPUT118), .ZN(n705) );
  XNOR2_X1 U765 ( .A(n706), .B(n705), .ZN(G51) );
  NAND2_X1 U766 ( .A1(n723), .A2(G469), .ZN(n711) );
  XOR2_X1 U767 ( .A(KEYINPUT120), .B(KEYINPUT119), .Z(n708) );
  XNOR2_X1 U768 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n707) );
  XNOR2_X1 U769 ( .A(n711), .B(n710), .ZN(n712) );
  NOR2_X1 U770 ( .A1(n727), .A2(n712), .ZN(G54) );
  NAND2_X1 U771 ( .A1(n723), .A2(G475), .ZN(n716) );
  XOR2_X1 U772 ( .A(KEYINPUT59), .B(KEYINPUT88), .Z(n713) );
  XNOR2_X1 U773 ( .A(n714), .B(n713), .ZN(n715) );
  NAND2_X1 U774 ( .A1(n723), .A2(G478), .ZN(n721) );
  NAND2_X1 U775 ( .A1(G217), .A2(n723), .ZN(n724) );
  XNOR2_X1 U776 ( .A(n725), .B(n724), .ZN(n726) );
  NOR2_X1 U777 ( .A1(n727), .A2(n726), .ZN(G66) );
  NOR2_X1 U778 ( .A1(G898), .A2(n490), .ZN(n730) );
  XOR2_X1 U779 ( .A(n728), .B(KEYINPUT124), .Z(n729) );
  NOR2_X1 U780 ( .A1(n730), .A2(n729), .ZN(n738) );
  XOR2_X1 U781 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n732) );
  NAND2_X1 U782 ( .A1(G224), .A2(G953), .ZN(n731) );
  XNOR2_X1 U783 ( .A(n732), .B(n731), .ZN(n733) );
  NAND2_X1 U784 ( .A1(n733), .A2(G898), .ZN(n736) );
  NAND2_X1 U785 ( .A1(n734), .A2(n490), .ZN(n735) );
  NAND2_X1 U786 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U787 ( .A(n738), .B(n737), .ZN(G69) );
  XNOR2_X1 U788 ( .A(n739), .B(KEYINPUT125), .ZN(n741) );
  XOR2_X1 U789 ( .A(n741), .B(n740), .Z(n745) );
  XOR2_X1 U790 ( .A(n745), .B(n742), .Z(n743) );
  NAND2_X1 U791 ( .A1(n743), .A2(n490), .ZN(n744) );
  XNOR2_X1 U792 ( .A(n744), .B(KEYINPUT126), .ZN(n749) );
  XNOR2_X1 U793 ( .A(G227), .B(n745), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n746), .A2(G900), .ZN(n747) );
  NAND2_X1 U795 ( .A1(n747), .A2(G953), .ZN(n748) );
  NAND2_X1 U796 ( .A1(n749), .A2(n748), .ZN(G72) );
  XOR2_X1 U797 ( .A(n750), .B(G122), .Z(G24) );
  XOR2_X1 U798 ( .A(KEYINPUT113), .B(KEYINPUT37), .Z(n753) );
  XNOR2_X1 U799 ( .A(n751), .B(G125), .ZN(n752) );
  XNOR2_X1 U800 ( .A(n753), .B(n752), .ZN(G27) );
  XNOR2_X1 U801 ( .A(G119), .B(n754), .ZN(G21) );
  XNOR2_X1 U802 ( .A(G131), .B(n755), .ZN(G33) );
  XOR2_X1 U803 ( .A(G137), .B(n756), .Z(n757) );
  XNOR2_X1 U804 ( .A(KEYINPUT127), .B(n757), .ZN(G39) );
endmodule

