//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 0 1 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1274, new_n1275, new_n1276, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1342, new_n1343, new_n1344;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G107), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  INV_X1    g0023(.A(G97), .ZN(new_n224));
  INV_X1    g0024(.A(G257), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n222), .B1(new_n202), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n206), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n209), .B(new_n215), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(new_n223), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XOR2_X1   g0038(.A(G50), .B(G58), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  NAND3_X1  g0044(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n245));
  AND2_X1   g0045(.A1(new_n245), .A2(new_n212), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT8), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G58), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n213), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n250), .A2(new_n252), .B1(G150), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n246), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G13), .A3(G20), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n246), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(G20), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G50), .ZN(new_n261));
  OAI22_X1  g0061(.A1(new_n259), .A2(new_n261), .B1(G50), .B2(new_n258), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(G1), .A3(G13), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT65), .ZN(new_n266));
  AND2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT3), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n272), .A2(KEYINPUT65), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G77), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n269), .A2(new_n274), .A3(G223), .A4(G1698), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n269), .A2(new_n274), .A3(G222), .A4(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n276), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n265), .B1(new_n280), .B2(KEYINPUT66), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT66), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n276), .A2(new_n282), .A3(new_n277), .A4(new_n279), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT64), .ZN(new_n285));
  AND2_X1   g0085(.A1(G33), .A2(G41), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n285), .B1(new_n286), .B2(new_n212), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n264), .A2(KEYINPUT64), .A3(G1), .A4(G13), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n287), .A2(new_n289), .A3(G274), .A4(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n287), .A2(new_n290), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(new_n289), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n292), .B1(G226), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n284), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G169), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n263), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G179), .ZN(new_n299));
  INV_X1    g0099(.A(new_n295), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n300), .B1(new_n281), .B2(new_n283), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n298), .A2(KEYINPUT67), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n302), .B1(KEYINPUT67), .B2(new_n298), .ZN(new_n303));
  INV_X1    g0103(.A(G68), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G20), .ZN(new_n305));
  INV_X1    g0105(.A(new_n253), .ZN(new_n306));
  OAI221_X1 g0106(.A(new_n305), .B1(new_n251), .B2(new_n217), .C1(new_n306), .C2(new_n201), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n245), .A2(new_n212), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT11), .ZN(new_n310));
  INV_X1    g0110(.A(G13), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n311), .A2(G1), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT70), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n312), .A2(new_n313), .A3(G20), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n258), .A2(KEYINPUT70), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT12), .B1(new_n316), .B2(G68), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT12), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n317), .B1(new_n305), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n308), .B1(new_n314), .B2(new_n315), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n321), .A2(G68), .A3(new_n260), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n310), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT14), .ZN(new_n324));
  NOR2_X1   g0124(.A1(G226), .A2(G1698), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n325), .B1(new_n223), .B2(G1698), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n269), .A2(new_n326), .A3(new_n274), .ZN(new_n327));
  NAND2_X1  g0127(.A1(G33), .A2(G97), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n265), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n287), .A2(G238), .A3(new_n290), .A4(new_n288), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n291), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT13), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n329), .A2(new_n331), .A3(KEYINPUT13), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n324), .B(G169), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n329), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT13), .ZN(new_n337));
  INV_X1    g0137(.A(new_n331), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n339), .A2(G179), .A3(new_n332), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n339), .A2(new_n332), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n324), .B1(new_n342), .B2(G169), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n323), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G190), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n346), .A2(new_n323), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n342), .A2(G200), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n250), .A2(new_n253), .B1(G20), .B2(G77), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT15), .B(G87), .ZN(new_n351));
  OAI21_X1  g0151(.A(KEYINPUT69), .B1(new_n351), .B2(new_n251), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n351), .A2(KEYINPUT69), .A3(new_n251), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n308), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n217), .B1(new_n257), .B2(G20), .ZN(new_n356));
  XNOR2_X1  g0156(.A(new_n258), .B(new_n313), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n321), .A2(new_n356), .B1(new_n357), .B2(new_n217), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n292), .B1(G244), .B2(new_n294), .ZN(new_n360));
  OR2_X1    g0160(.A1(KEYINPUT68), .A2(G107), .ZN(new_n361));
  NAND2_X1  g0161(.A1(KEYINPUT68), .A2(G107), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n265), .B1(new_n275), .B2(new_n364), .ZN(new_n365));
  MUX2_X1   g0165(.A(G232), .B(G238), .S(G1698), .Z(new_n366));
  OAI21_X1  g0166(.A(new_n365), .B1(new_n275), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n360), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n359), .B1(new_n297), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(G179), .B2(new_n368), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(G200), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n371), .B(new_n359), .C1(new_n345), .C2(new_n368), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n303), .A2(new_n344), .A3(new_n349), .A4(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n259), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n250), .A2(new_n260), .ZN(new_n376));
  INV_X1    g0176(.A(new_n258), .ZN(new_n377));
  INV_X1    g0177(.A(new_n250), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n375), .A2(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OR2_X1    g0179(.A1(G223), .A2(G1698), .ZN(new_n380));
  INV_X1    g0180(.A(G226), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(G1698), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n380), .B(new_n382), .C1(new_n267), .C2(new_n268), .ZN(new_n383));
  NAND2_X1  g0183(.A1(G33), .A2(G87), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n265), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n385), .A2(G190), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT74), .ZN(new_n387));
  NOR2_X1   g0187(.A1(G41), .A2(G45), .ZN(new_n388));
  OAI21_X1  g0188(.A(G232), .B1(new_n388), .B2(G1), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n257), .B(G274), .C1(G41), .C2(G45), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n387), .B1(new_n391), .B2(new_n293), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n389), .A2(new_n390), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n393), .A2(KEYINPUT74), .A3(new_n287), .A4(new_n290), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n386), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G200), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n391), .A2(new_n293), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n396), .B1(new_n397), .B2(new_n385), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  XOR2_X1   g0199(.A(KEYINPUT72), .B(KEYINPUT16), .Z(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT7), .B1(new_n275), .B2(new_n213), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n272), .A2(KEYINPUT7), .A3(new_n213), .A4(new_n273), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT73), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n267), .A2(new_n268), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT73), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT7), .A4(new_n213), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(G68), .B1(new_n402), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n202), .A2(new_n304), .ZN(new_n410));
  NOR2_X1   g0210(.A1(G58), .A2(G68), .ZN(new_n411));
  OAI21_X1  g0211(.A(G20), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n253), .A2(G159), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n401), .B1(new_n409), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT7), .B1(new_n405), .B2(new_n213), .ZN(new_n417));
  INV_X1    g0217(.A(new_n403), .ZN(new_n418));
  OAI21_X1  g0218(.A(G68), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n419), .A2(KEYINPUT16), .A3(new_n415), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n308), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n379), .B(new_n399), .C1(new_n416), .C2(new_n421), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n422), .B(KEYINPUT17), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n383), .A2(new_n384), .ZN(new_n424));
  INV_X1    g0224(.A(new_n265), .ZN(new_n425));
  AOI21_X1  g0225(.A(G179), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n426), .A2(new_n392), .A3(new_n394), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT75), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT75), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n426), .A2(new_n392), .A3(new_n429), .A4(new_n394), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n297), .B1(new_n397), .B2(new_n385), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT76), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT76), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n428), .A2(new_n434), .A3(new_n430), .A4(new_n431), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n379), .B1(new_n416), .B2(new_n421), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n433), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT18), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT18), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n433), .A2(new_n439), .A3(new_n435), .A4(new_n436), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n423), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n296), .A2(G200), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n284), .A2(G190), .A3(new_n295), .ZN(new_n443));
  XNOR2_X1  g0243(.A(new_n263), .B(KEYINPUT9), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT10), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(KEYINPUT71), .A3(new_n443), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n444), .B1(G190), .B2(new_n301), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n450), .B(new_n442), .C1(KEYINPUT71), .C2(KEYINPUT10), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n374), .A2(new_n441), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(G116), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n454), .B1(new_n257), .B2(G33), .ZN(new_n455));
  OAI22_X1  g0255(.A1(new_n321), .A2(new_n454), .B1(new_n357), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G283), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n457), .B(new_n213), .C1(G33), .C2(new_n224), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n454), .A2(G20), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(new_n308), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT20), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n458), .A2(KEYINPUT20), .A3(new_n308), .A4(new_n459), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n456), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT79), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT79), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n456), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  XOR2_X1   g0269(.A(KEYINPUT78), .B(G303), .Z(new_n470));
  AOI21_X1  g0270(.A(new_n470), .B1(new_n269), .B2(new_n274), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n220), .A2(G1698), .ZN(new_n472));
  OAI221_X1 g0272(.A(new_n472), .B1(G257), .B2(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n425), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(G45), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(G1), .ZN(new_n477));
  AND2_X1   g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  NOR2_X1   g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n480), .A2(new_n287), .A3(G270), .A4(new_n290), .ZN(new_n481));
  XNOR2_X1  g0281(.A(KEYINPUT5), .B(G41), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n257), .A2(G45), .A3(G274), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n287), .A2(new_n482), .A3(new_n484), .A4(new_n290), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n297), .B1(new_n475), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n469), .A2(KEYINPUT21), .A3(new_n487), .ZN(new_n488));
  AND3_X1   g0288(.A1(new_n456), .A2(new_n464), .A3(new_n467), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n467), .B1(new_n456), .B2(new_n464), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT21), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n475), .A2(G179), .A3(new_n486), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n469), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n475), .A2(new_n486), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G200), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n475), .A2(new_n486), .A3(G190), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n497), .A2(new_n466), .A3(new_n468), .A4(new_n498), .ZN(new_n499));
  AND4_X1   g0299(.A1(new_n488), .A2(new_n493), .A3(new_n495), .A4(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT22), .ZN(new_n501));
  INV_X1    g0301(.A(G87), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n501), .B1(new_n275), .B2(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(KEYINPUT22), .B(G87), .C1(new_n267), .C2(new_n268), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G116), .ZN(new_n505));
  AOI21_X1  g0305(.A(G20), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n361), .A2(G20), .A3(new_n362), .ZN(new_n508));
  OAI21_X1  g0308(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n508), .A2(KEYINPUT23), .B1(G20), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n503), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(KEYINPUT24), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT24), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n508), .A2(KEYINPUT23), .ZN(new_n514));
  INV_X1    g0314(.A(new_n509), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n514), .B1(new_n213), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n516), .A2(new_n506), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n513), .B1(new_n517), .B2(new_n503), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n308), .B1(new_n512), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n377), .A2(new_n219), .ZN(new_n520));
  XNOR2_X1  g0320(.A(new_n520), .B(KEYINPUT25), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n246), .B(new_n258), .C1(G1), .C2(new_n271), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n522), .A2(new_n219), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n480), .A2(new_n287), .A3(G264), .A4(new_n290), .ZN(new_n525));
  NOR2_X1   g0325(.A1(G250), .A2(G1698), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n526), .B1(new_n225), .B2(G1698), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n272), .A2(new_n273), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n527), .A2(new_n528), .B1(G33), .B2(G294), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n485), .B(new_n525), .C1(new_n529), .C2(new_n265), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n396), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(G190), .B2(new_n530), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n519), .A2(new_n524), .A3(new_n532), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n480), .A2(new_n287), .A3(new_n290), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n225), .A2(G1698), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(G250), .B2(G1698), .ZN(new_n536));
  INV_X1    g0336(.A(G294), .ZN(new_n537));
  OAI22_X1  g0337(.A1(new_n536), .A2(new_n405), .B1(new_n271), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n534), .A2(G264), .B1(new_n538), .B2(new_n425), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n539), .A2(KEYINPUT80), .A3(G179), .A4(new_n485), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT80), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n541), .B1(new_n530), .B2(G169), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n530), .A2(new_n299), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n511), .A2(KEYINPUT24), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n517), .A2(new_n513), .A3(new_n503), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n246), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n524), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n544), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n533), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(G250), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n483), .B1(new_n477), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n552), .A2(new_n287), .A3(new_n290), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT77), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n218), .A2(G1698), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(G238), .B2(G1698), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n505), .B1(new_n557), .B2(new_n405), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n425), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n552), .A2(KEYINPUT77), .A3(new_n287), .A4(new_n290), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n555), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G200), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n304), .A2(G20), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT19), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n213), .A2(G33), .A3(G97), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n528), .A2(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n213), .B1(new_n328), .B2(new_n564), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n502), .A2(new_n224), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n567), .B1(new_n363), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n246), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n522), .A2(new_n502), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n314), .A2(new_n315), .A3(new_n351), .ZN(new_n572));
  NOR3_X1   g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n554), .A2(new_n553), .B1(new_n558), .B2(new_n425), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n574), .A2(G190), .A3(new_n560), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n562), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n561), .A2(new_n297), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n574), .A2(new_n299), .A3(new_n560), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n566), .A2(new_n569), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n308), .ZN(new_n580));
  OR2_X1    g0380(.A1(new_n522), .A2(new_n351), .ZN(new_n581));
  INV_X1    g0381(.A(new_n572), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n577), .A2(new_n578), .A3(new_n583), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n576), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT7), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n269), .A2(new_n274), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n586), .B1(new_n587), .B2(G20), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n404), .A2(new_n407), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n364), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT6), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n591), .A2(new_n224), .A3(G107), .ZN(new_n592));
  XNOR2_X1  g0392(.A(G97), .B(G107), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n592), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  OAI22_X1  g0394(.A1(new_n594), .A2(new_n213), .B1(new_n217), .B2(new_n306), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n308), .B1(new_n590), .B2(new_n595), .ZN(new_n596));
  MUX2_X1   g0396(.A(new_n258), .B(new_n522), .S(G97), .Z(new_n597));
  NAND4_X1  g0397(.A1(new_n480), .A2(new_n287), .A3(G257), .A4(new_n290), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n485), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n269), .A2(new_n274), .A3(G250), .A4(G1698), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT4), .ZN(new_n601));
  NOR3_X1   g0401(.A1(new_n601), .A2(new_n218), .A3(G1698), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n269), .A2(new_n274), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n278), .A2(G244), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n601), .B1(new_n405), .B2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n600), .A2(new_n603), .A3(new_n457), .A4(new_n605), .ZN(new_n606));
  AOI211_X1 g0406(.A(G190), .B(new_n599), .C1(new_n606), .C2(new_n425), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n425), .ZN(new_n608));
  INV_X1    g0408(.A(new_n599), .ZN(new_n609));
  AOI21_X1  g0409(.A(G200), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n596), .B(new_n597), .C1(new_n607), .C2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(G20), .B1(new_n269), .B2(new_n274), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n404), .B(new_n407), .C1(new_n612), .C2(KEYINPUT7), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n595), .B1(new_n613), .B2(new_n363), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n597), .B1(new_n614), .B2(new_n246), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n608), .A2(new_n609), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n297), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n599), .B1(new_n606), .B2(new_n425), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n299), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n615), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n585), .A2(new_n611), .A3(new_n620), .ZN(new_n621));
  AND4_X1   g0421(.A1(new_n453), .A2(new_n500), .A3(new_n550), .A4(new_n621), .ZN(G372));
  INV_X1    g0422(.A(KEYINPUT84), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n452), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n449), .A2(new_n451), .A3(KEYINPUT84), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n370), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n349), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n344), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n629), .A2(new_n423), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n436), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n632), .B(new_n439), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n626), .B1(new_n630), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n303), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n585), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n638), .A2(new_n639), .A3(new_n620), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n620), .A2(KEYINPUT83), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT83), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n615), .A2(new_n617), .A3(new_n643), .A4(new_n619), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n396), .B1(new_n574), .B2(new_n560), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n522), .A2(new_n502), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n580), .A2(new_n647), .A3(new_n582), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT81), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT81), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n562), .A2(new_n573), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n649), .A2(new_n575), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(KEYINPUT82), .B1(new_n652), .B2(new_n584), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n652), .A2(KEYINPUT82), .A3(new_n584), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n645), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n641), .B1(new_n656), .B2(KEYINPUT26), .ZN(new_n657));
  INV_X1    g0457(.A(new_n584), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n533), .A2(new_n611), .A3(new_n620), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n493), .A2(new_n488), .A3(new_n495), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n549), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n654), .A2(new_n655), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n658), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n657), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n453), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n637), .A2(new_n665), .ZN(G369));
  NAND2_X1  g0466(.A1(new_n312), .A2(new_n213), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G213), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G343), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n469), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g0473(.A(new_n673), .B(KEYINPUT85), .Z(new_n674));
  INV_X1    g0474(.A(new_n660), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT86), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n674), .A2(new_n675), .A3(KEYINPUT86), .ZN(new_n679));
  INV_X1    g0479(.A(new_n500), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n678), .B(new_n679), .C1(new_n680), .C2(new_n674), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n672), .B1(new_n547), .B2(new_n548), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n550), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n549), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n672), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n681), .A2(G330), .A3(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n660), .A2(new_n672), .ZN(new_n688));
  INV_X1    g0488(.A(new_n672), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n688), .A2(new_n550), .B1(new_n684), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n687), .A2(new_n690), .ZN(G399));
  NOR3_X1   g0491(.A1(new_n363), .A2(G116), .A3(new_n568), .ZN(new_n692));
  XOR2_X1   g0492(.A(new_n692), .B(KEYINPUT87), .Z(new_n693));
  INV_X1    g0493(.A(new_n207), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G41), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G1), .ZN(new_n697));
  OAI22_X1  g0497(.A1(new_n693), .A2(new_n697), .B1(new_n210), .B2(new_n696), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n672), .B1(new_n657), .B2(new_n663), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n533), .A2(new_n611), .A3(new_n620), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n549), .A2(new_n493), .A3(new_n488), .A4(new_n495), .ZN(new_n704));
  INV_X1    g0504(.A(new_n655), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n703), .B(new_n704), .C1(new_n705), .C2(new_n653), .ZN(new_n706));
  OR3_X1    g0506(.A1(new_n620), .A2(new_n638), .A3(KEYINPUT26), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(new_n584), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n645), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n639), .B1(new_n662), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n689), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT29), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n702), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n500), .A2(new_n621), .A3(new_n550), .A4(new_n689), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT88), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n525), .B1(new_n529), .B2(new_n265), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n715), .B1(new_n561), .B2(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n539), .A2(new_n574), .A3(KEYINPUT88), .A4(new_n560), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n717), .A2(new_n494), .A3(new_n718), .A4(new_n618), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n475), .A2(new_n486), .A3(G179), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n616), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(KEYINPUT30), .A3(new_n718), .A4(new_n717), .ZN(new_n724));
  AOI21_X1  g0524(.A(G179), .B1(new_n475), .B2(new_n486), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n616), .A2(new_n725), .A3(new_n530), .A4(new_n561), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n721), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n672), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT31), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n727), .A2(KEYINPUT31), .A3(new_n672), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n714), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n713), .B1(G330), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n699), .B1(new_n733), .B2(G1), .ZN(G364));
  NOR2_X1   g0534(.A1(new_n311), .A2(G20), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G45), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n736), .A2(KEYINPUT89), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n257), .B1(new_n736), .B2(KEYINPUT89), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n695), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n740), .B1(new_n681), .B2(G330), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(G330), .B2(new_n681), .ZN(new_n742));
  INV_X1    g0542(.A(new_n740), .ZN(new_n743));
  NOR4_X1   g0543(.A1(new_n213), .A2(new_n299), .A3(new_n345), .A4(new_n396), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n213), .A2(G179), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(G190), .A3(G200), .ZN(new_n747));
  OAI22_X1  g0547(.A1(new_n745), .A2(new_n201), .B1(new_n747), .B2(new_n502), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n213), .A2(new_n299), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(new_n345), .A3(G200), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n748), .B1(G68), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n746), .A2(new_n345), .A3(G200), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n753), .A2(KEYINPUT95), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(KEYINPUT95), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G107), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n299), .A2(new_n396), .A3(G190), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT96), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n752), .B(new_n758), .C1(new_n224), .C2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G190), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n746), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G159), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g0567(.A(KEYINPUT94), .B(KEYINPUT32), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n749), .A2(G190), .A3(new_n396), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n275), .B1(G58), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n749), .A2(new_n764), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT93), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n773), .A2(new_n774), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n769), .B(new_n772), .C1(new_n779), .C2(new_n217), .ZN(new_n780));
  INV_X1    g0580(.A(G311), .ZN(new_n781));
  INV_X1    g0581(.A(G329), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n773), .A2(new_n781), .B1(new_n765), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(G322), .B2(new_n771), .ZN(new_n784));
  INV_X1    g0584(.A(new_n747), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n587), .B1(G303), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G317), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(KEYINPUT33), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n787), .A2(KEYINPUT33), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n751), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n744), .A2(G326), .B1(G294), .B2(new_n760), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n784), .A2(new_n786), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G283), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n756), .A2(new_n793), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n763), .A2(new_n780), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n212), .B1(G20), .B2(new_n297), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n743), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n275), .A2(new_n694), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n798), .A2(G355), .B1(new_n454), .B2(new_n694), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n240), .A2(G45), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT90), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n694), .A2(new_n528), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(G45), .B2(new_n210), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n799), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT91), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NOR2_X1   g0607(.A1(G13), .A2(G33), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT92), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(G20), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(new_n796), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n810), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n797), .B1(new_n806), .B2(new_n812), .C1(new_n681), .C2(new_n813), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n742), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(G396));
  NAND2_X1  g0616(.A1(new_n627), .A2(new_n689), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n372), .B1(new_n359), .B2(new_n689), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n370), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n700), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n732), .A2(G330), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n740), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n823), .B2(new_n822), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n796), .A2(new_n808), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n743), .B1(new_n217), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n796), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n771), .A2(G143), .B1(new_n744), .B2(G137), .ZN(new_n829));
  INV_X1    g0629(.A(G150), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n829), .B1(new_n830), .B2(new_n750), .C1(new_n779), .C2(new_n766), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT34), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n757), .A2(G68), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n747), .A2(new_n201), .ZN(new_n835));
  INV_X1    g0635(.A(G132), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n528), .B1(new_n765), .B2(new_n836), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n835), .B(new_n837), .C1(G58), .C2(new_n760), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(new_n831), .B2(new_n832), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n275), .B1(new_n781), .B2(new_n765), .C1(new_n537), .C2(new_n770), .ZN(new_n841));
  AOI22_X1  g0641(.A1(G283), .A2(new_n751), .B1(new_n785), .B2(G107), .ZN(new_n842));
  INV_X1    g0642(.A(G303), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n842), .B1(new_n843), .B2(new_n745), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n841), .B(new_n844), .C1(G116), .C2(new_n778), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n757), .A2(G87), .B1(G97), .B2(new_n761), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n833), .A2(new_n840), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n827), .B1(new_n828), .B2(new_n847), .C1(new_n821), .C2(new_n809), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n825), .A2(new_n848), .ZN(G384));
  INV_X1    g0649(.A(new_n594), .ZN(new_n850));
  OR2_X1    g0650(.A1(new_n850), .A2(KEYINPUT35), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(KEYINPUT35), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n851), .A2(G116), .A3(new_n214), .A4(new_n852), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n853), .B(KEYINPUT36), .Z(new_n854));
  OAI211_X1 g0654(.A(new_n211), .B(G77), .C1(new_n202), .C2(new_n304), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n201), .A2(G68), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n257), .B(G13), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  INV_X1    g0659(.A(new_n670), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n436), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n437), .A2(new_n859), .A3(new_n422), .A4(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n419), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n400), .B1(new_n863), .B2(new_n414), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n864), .A2(new_n420), .A3(new_n308), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n432), .A2(new_n670), .B1(new_n865), .B2(new_n379), .ZN(new_n866));
  INV_X1    g0666(.A(new_n422), .ZN(new_n867));
  OAI21_X1  g0667(.A(KEYINPUT37), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n862), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT98), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n670), .B1(new_n865), .B2(new_n379), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n441), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n862), .A2(KEYINPUT98), .A3(new_n868), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n871), .A2(new_n873), .A3(KEYINPUT38), .A4(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n861), .B1(new_n633), .B2(new_n423), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n437), .A2(new_n859), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n861), .A2(new_n422), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n632), .A2(new_n861), .A3(new_n422), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n878), .A2(new_n879), .B1(KEYINPUT37), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n876), .B1(new_n877), .B2(new_n881), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n875), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT100), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n732), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n714), .A2(new_n730), .A3(KEYINPUT100), .A4(new_n731), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT97), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n344), .A2(new_n887), .ZN(new_n888));
  OAI211_X1 g0688(.A(KEYINPUT97), .B(new_n323), .C1(new_n341), .C2(new_n343), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n323), .A2(new_n672), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(new_n347), .B2(new_n348), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n890), .B1(new_n341), .B2(new_n343), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n820), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n885), .A2(new_n886), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT40), .B1(new_n883), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n876), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n875), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n885), .A2(new_n886), .A3(new_n894), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT40), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n896), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n453), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n885), .A2(new_n886), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n903), .A2(new_n906), .ZN(new_n908));
  INV_X1    g0708(.A(G330), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n875), .A2(new_n882), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT39), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n898), .A2(KEYINPUT39), .A3(new_n875), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n888), .A2(new_n889), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n689), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT99), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT99), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n915), .A2(new_n918), .A3(new_n689), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n913), .A2(new_n914), .A3(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n642), .B(new_n644), .C1(new_n705), .C2(new_n653), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n640), .B1(new_n922), .B2(new_n639), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n706), .A2(new_n584), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n689), .B(new_n821), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n817), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n892), .A2(new_n893), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n926), .A2(new_n899), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n634), .A2(new_n670), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n921), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n904), .B1(new_n702), .B2(new_n712), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n931), .A2(new_n636), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n930), .B(new_n932), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n910), .A2(new_n933), .B1(new_n257), .B2(new_n735), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n910), .A2(new_n933), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n858), .B1(new_n934), .B2(new_n935), .ZN(G367));
  INV_X1    g0736(.A(KEYINPUT105), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT101), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT42), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n688), .A2(new_n550), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n620), .A2(new_n689), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n615), .A2(new_n672), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n611), .A2(new_n620), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n939), .B1(new_n940), .B2(new_n945), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n688), .A2(KEYINPUT42), .A3(new_n550), .A4(new_n944), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n620), .B1(new_n943), .B2(new_n549), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n946), .A2(new_n947), .B1(new_n689), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n662), .B1(new_n573), .B2(new_n689), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n658), .A2(new_n648), .A3(new_n672), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n938), .B1(new_n950), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n949), .A2(KEYINPUT101), .A3(new_n954), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n687), .A2(new_n945), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n950), .A2(new_n955), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n958), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(KEYINPUT102), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT102), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n958), .A2(new_n964), .A3(new_n959), .A4(new_n961), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n958), .A2(new_n961), .ZN(new_n967));
  INV_X1    g0767(.A(new_n959), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT104), .ZN(new_n971));
  XNOR2_X1  g0771(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n690), .B2(new_n944), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(KEYINPUT45), .B1(new_n690), .B2(new_n944), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n690), .A2(KEYINPUT45), .A3(new_n944), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n971), .A2(new_n974), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n690), .ZN(new_n979));
  INV_X1    g0779(.A(new_n972), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n979), .A2(new_n945), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n981), .A2(new_n973), .A3(KEYINPUT104), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n978), .A2(new_n687), .A3(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n687), .ZN(new_n984));
  AND3_X1   g0784(.A1(new_n981), .A2(new_n973), .A3(KEYINPUT104), .ZN(new_n985));
  INV_X1    g0785(.A(new_n977), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n986), .A2(new_n975), .B1(new_n973), .B2(KEYINPUT104), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n984), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n983), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n681), .A2(G330), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n940), .B1(new_n686), .B2(new_n688), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n990), .B(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n733), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n695), .B(KEYINPUT41), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n739), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n937), .B1(new_n970), .B2(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n963), .A2(new_n965), .B1(new_n968), .B2(new_n967), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n993), .A2(new_n994), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n997), .B(KEYINPUT105), .C1(new_n998), .C2(new_n739), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n802), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n811), .B1(new_n207), .B2(new_n351), .C1(new_n236), .C2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT106), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n743), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n778), .A2(G283), .B1(new_n363), .B2(new_n760), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT107), .Z(new_n1006));
  NAND2_X1  g0806(.A1(new_n757), .A2(G97), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n785), .A2(G116), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT46), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n405), .B1(new_n765), .B2(new_n787), .C1(new_n770), .C2(new_n470), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n751), .A2(G294), .B1(new_n744), .B2(G311), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1007), .A2(new_n1009), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1006), .A2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT108), .ZN(new_n1015));
  XOR2_X1   g0815(.A(KEYINPUT109), .B(G137), .Z(new_n1016));
  OAI221_X1 g0816(.A(new_n587), .B1(new_n830), .B2(new_n770), .C1(new_n765), .C2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(G50), .B2(new_n778), .ZN(new_n1018));
  INV_X1    g0818(.A(G143), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n745), .A2(new_n1019), .B1(new_n766), .B2(new_n750), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G58), .B2(new_n785), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n757), .A2(G77), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n761), .A2(G68), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1018), .A2(new_n1021), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1015), .A2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT47), .Z(new_n1026));
  OAI221_X1 g0826(.A(new_n1004), .B1(new_n1003), .B2(new_n1002), .C1(new_n1026), .C2(new_n828), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n953), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1027), .B1(new_n810), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1000), .A2(new_n1030), .ZN(G387));
  INV_X1    g0831(.A(new_n992), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n739), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n233), .A2(new_n476), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n1034), .A2(new_n802), .B1(new_n693), .B2(new_n798), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n250), .A2(new_n201), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT50), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n476), .B1(new_n304), .B2(new_n217), .ZN(new_n1038));
  NOR3_X1   g0838(.A1(new_n693), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n1035), .A2(new_n1039), .B1(G107), .B2(new_n207), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n743), .B1(new_n1040), .B2(new_n811), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n762), .A2(new_n351), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n770), .A2(new_n201), .B1(new_n773), .B2(new_n304), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n765), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n405), .B(new_n1044), .C1(G150), .C2(new_n1045), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n745), .A2(new_n766), .B1(new_n747), .B2(new_n217), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n250), .B2(new_n751), .ZN(new_n1048));
  AND4_X1   g0848(.A1(new_n1007), .A2(new_n1043), .A3(new_n1046), .A4(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n785), .A2(G294), .B1(new_n760), .B2(G283), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT110), .Z(new_n1051));
  AOI22_X1  g0851(.A1(G311), .A2(new_n751), .B1(new_n771), .B2(G317), .ZN(new_n1052));
  INV_X1    g0852(.A(G322), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1052), .B1(new_n1053), .B2(new_n745), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n470), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1054), .B1(new_n1055), .B2(new_n778), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1051), .B1(new_n1056), .B2(KEYINPUT48), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT111), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1056), .A2(KEYINPUT48), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1060), .A2(KEYINPUT49), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n528), .B1(new_n1045), .B2(G326), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n756), .B2(new_n454), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n1060), .B2(KEYINPUT49), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1049), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1041), .B1(new_n686), .B2(new_n813), .C1(new_n1065), .C2(new_n828), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1033), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1032), .A2(new_n733), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n695), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1032), .A2(new_n733), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1067), .B1(new_n1069), .B2(new_n1070), .ZN(G393));
  NAND2_X1  g0871(.A1(new_n983), .A2(KEYINPUT112), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT112), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n978), .A2(new_n1073), .A3(new_n687), .A4(new_n982), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1072), .A2(new_n988), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n739), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n811), .B1(new_n224), .B2(new_n207), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n243), .A2(new_n1001), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n740), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n745), .A2(new_n787), .B1(new_n781), .B2(new_n770), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT52), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n760), .A2(G116), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n793), .B2(new_n747), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n1055), .B2(new_n751), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n773), .A2(new_n537), .B1(new_n765), .B2(new_n1053), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1086), .A2(new_n587), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1082), .A2(new_n1085), .A3(new_n758), .A4(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n778), .A2(new_n250), .B1(G50), .B2(new_n751), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1090), .A2(KEYINPUT113), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(KEYINPUT113), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n528), .B1(new_n765), .B2(new_n1019), .C1(new_n304), .C2(new_n747), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n757), .B2(G87), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1091), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n745), .A2(new_n830), .B1(new_n766), .B2(new_n770), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT51), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n761), .A2(G77), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1088), .B1(new_n1095), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1080), .B1(new_n1102), .B2(new_n796), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n944), .B2(new_n813), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1075), .A2(new_n1068), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n695), .B1(new_n1068), .B2(new_n989), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1077), .B(new_n1104), .C1(new_n1105), .C2(new_n1106), .ZN(G390));
  NOR3_X1   g0907(.A1(new_n904), .A2(new_n909), .A3(new_n905), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n931), .A2(new_n1108), .A3(new_n636), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT114), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n927), .B(new_n1110), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n885), .A2(G330), .A3(new_n821), .A4(new_n886), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n689), .B(new_n819), .C1(new_n708), .C2(new_n710), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1114), .A2(new_n817), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n927), .A2(new_n732), .A3(G330), .A4(new_n821), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1113), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n927), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n823), .B2(new_n820), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n885), .A2(G330), .A3(new_n886), .A4(new_n894), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n926), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1117), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1109), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT115), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1114), .A2(new_n817), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n927), .B(KEYINPUT114), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n920), .B1(new_n875), .B2(new_n882), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n913), .A2(new_n914), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n920), .B1(new_n926), .B2(new_n927), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1131), .B(new_n1116), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n905), .A2(new_n909), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1135), .A2(new_n894), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1126), .A2(new_n1134), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n920), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n817), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n700), .B2(new_n821), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1139), .B1(new_n1141), .B2(new_n1118), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n913), .A2(new_n914), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1142), .A2(new_n1143), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1144), .A2(new_n1120), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1134), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1125), .B(new_n1124), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1138), .A2(new_n1147), .A3(new_n695), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1137), .A2(new_n739), .A3(new_n1134), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n743), .B1(new_n378), .B2(new_n826), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n275), .B1(new_n537), .B2(new_n765), .C1(new_n454), .C2(new_n770), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n778), .B2(G97), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n745), .A2(new_n793), .B1(new_n747), .B2(new_n502), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n363), .B2(new_n751), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1152), .A2(new_n1154), .A3(new_n834), .A4(new_n1099), .ZN(new_n1155));
  INV_X1    g0955(.A(G128), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n745), .A2(new_n1156), .B1(new_n750), .B2(new_n1016), .ZN(new_n1157));
  INV_X1    g0957(.A(G125), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n770), .A2(new_n836), .B1(new_n765), .B2(new_n1158), .ZN(new_n1159));
  NOR3_X1   g0959(.A1(new_n1157), .A2(new_n275), .A3(new_n1159), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n1160), .B1(new_n201), .B2(new_n756), .C1(new_n766), .C2(new_n762), .ZN(new_n1161));
  OR3_X1    g0961(.A1(new_n747), .A2(KEYINPUT53), .A3(new_n830), .ZN(new_n1162));
  OAI21_X1  g0962(.A(KEYINPUT53), .B1(new_n747), .B2(new_n830), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT54), .B(G143), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1162), .B(new_n1163), .C1(new_n779), .C2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1155), .B1(new_n1161), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT116), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n796), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1150), .B1(new_n1168), .B2(new_n1170), .C1(new_n1132), .C2(new_n809), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1149), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1148), .A2(new_n1172), .ZN(G378));
  NAND2_X1  g0973(.A1(new_n626), .A2(new_n303), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n263), .A2(new_n670), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  XOR2_X1   g0976(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1177));
  INV_X1    g0977(.A(new_n1175), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n625), .ZN(new_n1179));
  AOI21_X1  g0979(.A(KEYINPUT84), .B1(new_n449), .B2(new_n451), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n303), .B(new_n1178), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1176), .A2(new_n1177), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1177), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1181), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1178), .B1(new_n626), .B2(new_n303), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1183), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1182), .A2(new_n1186), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n903), .A2(G330), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1187), .B1(new_n903), .B2(G330), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n930), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1182), .A2(new_n1186), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n911), .A2(new_n885), .A3(new_n886), .A4(new_n894), .ZN(new_n1192));
  AOI21_X1  g0992(.A(KEYINPUT40), .B1(new_n898), .B2(new_n875), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1192), .A2(KEYINPUT40), .B1(new_n1193), .B2(new_n900), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1191), .B1(new_n1194), .B2(new_n909), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n930), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n903), .A2(G330), .A3(new_n1187), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1190), .A2(new_n739), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n757), .A2(G58), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n765), .A2(new_n793), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n528), .A2(G41), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(G107), .C2(new_n771), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G77), .A2(new_n785), .B1(new_n744), .B2(G116), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1200), .A2(new_n1203), .A3(new_n1023), .A4(new_n1204), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n750), .A2(new_n224), .B1(new_n773), .B2(new_n351), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT117), .Z(new_n1207));
  NOR2_X1   g1007(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n1209));
  XOR2_X1   g1009(.A(new_n1208), .B(new_n1209), .Z(new_n1210));
  OAI211_X1 g1010(.A(new_n1202), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1211));
  INV_X1    g1011(.A(G137), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n770), .A2(new_n1156), .B1(new_n773), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1164), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1213), .B1(new_n785), .B2(new_n1214), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n751), .A2(G132), .B1(new_n744), .B2(G125), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(new_n830), .C2(new_n762), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(KEYINPUT59), .ZN(new_n1218));
  AOI211_X1 g1018(.A(G33), .B(G41), .C1(new_n1045), .C2(G124), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(new_n766), .C2(new_n756), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1217), .A2(KEYINPUT59), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1211), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n796), .B1(new_n1210), .B2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n743), .B1(new_n201), .B2(new_n826), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(new_n1191), .C2(new_n809), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1199), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1190), .A2(KEYINPUT57), .A3(new_n1198), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1134), .B(new_n1123), .C1(new_n1144), .C2(new_n1120), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1229), .A2(new_n1109), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n695), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1196), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1229), .A2(new_n1109), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT57), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1227), .B1(new_n1231), .B2(new_n1236), .ZN(G375));
  AND2_X1   g1037(.A1(new_n1117), .A2(new_n1122), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n931), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1108), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1239), .A2(new_n1240), .A3(new_n637), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1238), .A2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1242), .A2(new_n1124), .A3(new_n994), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT119), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n743), .B1(new_n304), .B2(new_n826), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1200), .A2(new_n528), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT120), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1045), .A2(G128), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n1249), .B1(new_n830), .B2(new_n773), .C1(new_n770), .C2(new_n1016), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n751), .A2(new_n1214), .B1(new_n744), .B2(G132), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n766), .B2(new_n747), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1250), .B(new_n1252), .C1(G50), .C2(new_n761), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n275), .B1(new_n843), .B2(new_n765), .C1(new_n793), .C2(new_n770), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(G116), .A2(new_n751), .B1(new_n785), .B2(G97), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n537), .B2(new_n745), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1254), .B(new_n1256), .C1(new_n363), .C2(new_n778), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1042), .B1(G77), .B2(new_n757), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1248), .A2(new_n1253), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n808), .ZN(new_n1260));
  OAI221_X1 g1060(.A(new_n1246), .B1(new_n828), .B2(new_n1259), .C1(new_n1128), .C2(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1261), .B1(new_n1238), .B2(new_n1076), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1262), .B(KEYINPUT121), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1245), .A2(new_n1263), .A3(new_n1264), .ZN(G381));
  INV_X1    g1065(.A(G390), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1000), .A2(new_n1030), .A3(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(G378), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1067), .B(new_n815), .C1(new_n1070), .C2(new_n1069), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(G381), .A2(G384), .A3(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1268), .A2(new_n1269), .A3(new_n1271), .ZN(new_n1272));
  OR2_X1    g1072(.A1(new_n1272), .A2(G375), .ZN(G407));
  NAND2_X1  g1073(.A1(new_n671), .A2(G213), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1269), .A2(new_n1275), .ZN(new_n1276));
  OAI211_X1 g1076(.A(G407), .B(G213), .C1(G375), .C2(new_n1276), .ZN(G409));
  AOI21_X1  g1077(.A(new_n1266), .B1(new_n1000), .B2(new_n1030), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT127), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G393), .A2(G396), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1279), .B1(new_n1280), .B2(new_n1270), .ZN(new_n1281));
  NOR3_X1   g1081(.A1(new_n1268), .A2(new_n1278), .A3(new_n1281), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1280), .A2(new_n1279), .A3(new_n1270), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1283), .A2(new_n1281), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(G387), .A2(G390), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1284), .B1(new_n1285), .B2(new_n1267), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1282), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT124), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT122), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1190), .A2(new_n994), .A3(new_n1198), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1289), .B1(new_n1290), .B2(new_n1230), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1234), .A2(KEYINPUT122), .A3(new_n994), .A4(new_n1235), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT123), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1226), .A2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1199), .A2(KEYINPUT123), .A3(new_n1225), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(G378), .B1(new_n1293), .B2(new_n1297), .ZN(new_n1298));
  OAI211_X1 g1098(.A(G378), .B(new_n1227), .C1(new_n1231), .C2(new_n1236), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1288), .B1(new_n1298), .B2(new_n1300), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1199), .A2(KEYINPUT123), .A3(new_n1225), .ZN(new_n1302));
  AOI21_X1  g1102(.A(KEYINPUT123), .B1(new_n1199), .B2(new_n1225), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1269), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1306), .A2(KEYINPUT124), .A3(new_n1299), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT125), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT60), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1308), .B1(new_n1242), .B2(new_n1309), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1238), .A2(new_n1241), .A3(KEYINPUT125), .A4(KEYINPUT60), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1242), .A2(new_n1309), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n696), .B1(new_n1109), .B2(new_n1123), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1310), .A2(new_n1311), .A3(new_n1312), .A4(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1263), .A2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1315), .A2(new_n825), .A3(new_n848), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1263), .A2(new_n1314), .A3(G384), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1301), .A2(new_n1274), .A3(new_n1307), .A4(new_n1319), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1320), .A2(KEYINPUT62), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1274), .B1(new_n1298), .B2(new_n1300), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1275), .A2(G2897), .ZN(new_n1323));
  XOR2_X1   g1123(.A(new_n1323), .B(KEYINPUT126), .Z(new_n1324));
  INV_X1    g1124(.A(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1318), .A2(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1316), .A2(new_n1317), .A3(new_n1324), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT61), .B1(new_n1322), .B2(new_n1328), .ZN(new_n1329));
  OAI211_X1 g1129(.A(new_n1274), .B(new_n1319), .C1(new_n1298), .C2(new_n1300), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(KEYINPUT62), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1329), .A2(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1287), .B1(new_n1321), .B2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT63), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1320), .A2(new_n1334), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1287), .A2(KEYINPUT61), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1301), .A2(new_n1274), .A3(new_n1307), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(new_n1328), .ZN(new_n1338));
  OR2_X1    g1138(.A1(new_n1330), .A2(new_n1334), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1335), .A2(new_n1336), .A3(new_n1338), .A4(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1333), .A2(new_n1340), .ZN(G405));
  AND2_X1   g1141(.A1(G375), .A2(new_n1269), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1342), .A2(new_n1300), .ZN(new_n1343));
  XNOR2_X1  g1143(.A(new_n1343), .B(new_n1318), .ZN(new_n1344));
  XNOR2_X1  g1144(.A(new_n1344), .B(new_n1287), .ZN(G402));
endmodule


