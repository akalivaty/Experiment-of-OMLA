//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n803, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1015, new_n1016;
  XNOR2_X1  g000(.A(KEYINPUT0), .B(G57gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G85gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G1gat), .B(G29gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G127gat), .B(G134gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT68), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(G127gat), .A2(G134gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(G127gat), .A2(G134gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(KEYINPUT68), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G120gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G113gat), .ZN(new_n215));
  INV_X1    g014(.A(G113gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G120gat), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n215), .A2(new_n217), .A3(KEYINPUT69), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT69), .B1(new_n215), .B2(new_n217), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT1), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n213), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n215), .A2(new_n217), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n223), .A2(new_n207), .A3(new_n221), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT70), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT70), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n223), .A2(new_n207), .A3(new_n226), .A4(new_n221), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G155gat), .B(G162gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(G141gat), .B(G148gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT2), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n230), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n230), .ZN(new_n235));
  OR2_X1    g034(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n236));
  INV_X1    g035(.A(G162gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT80), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT80), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G162gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n236), .A2(new_n238), .A3(new_n240), .A4(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT2), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n235), .B1(new_n243), .B2(KEYINPUT81), .ZN(new_n244));
  AND2_X1   g043(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT80), .B(G162gat), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n233), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT81), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n231), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n234), .B1(new_n244), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT82), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n229), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n234), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n230), .B1(new_n249), .B2(new_n250), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n242), .A2(new_n250), .A3(KEYINPUT2), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(new_n232), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n255), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NOR3_X1   g058(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT1), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n225), .B(new_n227), .C1(new_n260), .C2(new_n213), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT82), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n254), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n259), .A2(new_n261), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT4), .ZN(new_n266));
  NAND2_X1  g065(.A1(G225gat), .A2(G233gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT3), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n270), .A3(new_n261), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n264), .A2(new_n266), .A3(new_n267), .A4(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT5), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT83), .B1(new_n229), .B2(new_n252), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT83), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n275), .A3(new_n261), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n274), .A2(new_n262), .A3(new_n254), .A4(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n267), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT84), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n277), .A2(KEYINPUT84), .A3(new_n278), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n273), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n265), .A2(new_n263), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT85), .ZN(new_n285));
  NOR4_X1   g084(.A1(new_n259), .A2(new_n261), .A3(KEYINPUT85), .A4(KEYINPUT4), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n254), .A2(new_n262), .A3(KEYINPUT4), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n285), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  AND4_X1   g088(.A1(new_n283), .A2(new_n289), .A3(new_n267), .A4(new_n271), .ZN(new_n290));
  OAI211_X1 g089(.A(KEYINPUT6), .B(new_n206), .C1(new_n282), .C2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n206), .B1(new_n282), .B2(new_n290), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n293));
  INV_X1    g092(.A(new_n271), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT85), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n295), .B1(new_n265), .B2(new_n263), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n296), .A2(new_n286), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n294), .B1(new_n297), .B2(new_n288), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n298), .A2(new_n283), .A3(new_n267), .ZN(new_n299));
  INV_X1    g098(.A(new_n281), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n300), .A2(new_n279), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n299), .B(new_n205), .C1(new_n301), .C2(new_n273), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n292), .A2(new_n293), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT74), .ZN(new_n304));
  NAND2_X1  g103(.A1(G197gat), .A2(G204gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(G197gat), .A2(G204gat), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G197gat), .ZN(new_n309));
  INV_X1    g108(.A(G204gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n311), .A2(KEYINPUT74), .A3(new_n305), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT22), .ZN(new_n314));
  XOR2_X1   g113(.A(G211gat), .B(G218gat), .Z(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n317));
  INV_X1    g116(.A(G211gat), .ZN(new_n318));
  INV_X1    g117(.A(G218gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(new_n319), .A3(KEYINPUT22), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(new_n318), .B2(new_n319), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n313), .A2(new_n317), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n317), .B1(new_n313), .B2(new_n321), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n316), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT25), .ZN(new_n325));
  AND2_X1   g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n326), .A2(KEYINPUT64), .A3(KEYINPUT24), .ZN(new_n327));
  NAND3_X1  g126(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n328), .B1(G183gat), .B2(G190gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT64), .ZN(new_n330));
  NAND2_X1  g129(.A1(G183gat), .A2(G190gat), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT24), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n327), .A2(new_n329), .A3(new_n333), .ZN(new_n334));
  AND2_X1   g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT23), .ZN(new_n336));
  INV_X1    g135(.A(G169gat), .ZN(new_n337));
  INV_X1    g136(.A(G176gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n335), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n325), .B1(new_n334), .B2(new_n342), .ZN(new_n343));
  AND3_X1   g142(.A1(new_n331), .A2(KEYINPUT65), .A3(new_n332), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT65), .B1(new_n331), .B2(new_n332), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n344), .A2(new_n329), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n335), .ZN(new_n347));
  INV_X1    g146(.A(new_n340), .ZN(new_n348));
  NOR3_X1   g147(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n349));
  OAI211_X1 g148(.A(KEYINPUT25), .B(new_n347), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT66), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  AOI211_X1 g150(.A(new_n325), .B(new_n335), .C1(new_n339), .C2(new_n340), .ZN(new_n352));
  NOR2_X1   g151(.A1(G183gat), .A2(G190gat), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n353), .B1(new_n326), .B2(KEYINPUT24), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n331), .A2(new_n332), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT65), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT65), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n354), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT66), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n352), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n343), .A2(new_n351), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n337), .A2(new_n338), .ZN(new_n364));
  OR3_X1    g163(.A1(new_n364), .A2(KEYINPUT67), .A3(KEYINPUT26), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT26), .B1(new_n364), .B2(KEYINPUT67), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n365), .A2(new_n347), .A3(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT27), .B(G183gat), .ZN(new_n368));
  INV_X1    g167(.A(G190gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(KEYINPUT28), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT28), .B1(new_n368), .B2(new_n369), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n367), .B(new_n331), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n363), .A2(KEYINPUT76), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT76), .B1(new_n363), .B2(new_n373), .ZN(new_n375));
  INV_X1    g174(.A(G226gat), .ZN(new_n376));
  INV_X1    g175(.A(G233gat), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NOR3_X1   g178(.A1(new_n374), .A2(new_n375), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n373), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n378), .A2(KEYINPUT29), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n324), .B1(new_n380), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT77), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n381), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n378), .ZN(new_n389));
  NOR3_X1   g188(.A1(new_n306), .A2(new_n307), .A3(new_n304), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT74), .B1(new_n311), .B2(new_n305), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n321), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT75), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n313), .A2(new_n317), .A3(new_n321), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n393), .A2(new_n394), .B1(new_n314), .B2(new_n315), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n374), .A2(new_n375), .ZN(new_n396));
  INV_X1    g195(.A(new_n382), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n389), .B(new_n395), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT76), .ZN(new_n399));
  NOR3_X1   g198(.A1(new_n346), .A2(KEYINPUT66), .A3(new_n350), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n361), .B1(new_n352), .B2(new_n360), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n355), .A2(KEYINPUT64), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n358), .A2(new_n330), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n354), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT25), .B1(new_n404), .B2(new_n341), .ZN(new_n405));
  NOR3_X1   g204(.A1(new_n400), .A2(new_n401), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n373), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n399), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n363), .A2(KEYINPUT76), .A3(new_n373), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n378), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n383), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n411), .A2(KEYINPUT77), .A3(new_n324), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n387), .A2(new_n398), .A3(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G8gat), .B(G36gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(G92gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(KEYINPUT78), .ZN(new_n416));
  INV_X1    g215(.A(G64gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n413), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n387), .A2(new_n398), .A3(new_n412), .A4(new_n418), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(KEYINPUT30), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT77), .B1(new_n411), .B2(new_n324), .ZN(new_n423));
  AOI211_X1 g222(.A(new_n386), .B(new_n395), .C1(new_n410), .C2(new_n383), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT30), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n425), .A2(new_n426), .A3(new_n398), .A4(new_n418), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n291), .A2(new_n303), .B1(new_n422), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n393), .A2(new_n394), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT29), .B1(new_n429), .B2(new_n316), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n259), .ZN(new_n431));
  NAND2_X1  g230(.A1(G228gat), .A2(G233gat), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n431), .A2(new_n270), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT29), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n324), .B1(new_n269), .B2(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT87), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT86), .B1(new_n395), .B2(KEYINPUT29), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT86), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n324), .A2(new_n440), .A3(new_n435), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n439), .A2(new_n268), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n436), .B1(new_n442), .B2(new_n259), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n438), .B1(new_n443), .B2(new_n433), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT3), .B1(new_n430), .B2(new_n440), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n252), .B1(new_n445), .B2(new_n439), .ZN(new_n446));
  OAI211_X1 g245(.A(KEYINPUT87), .B(new_n432), .C1(new_n446), .C2(new_n436), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n437), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(G22gat), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT88), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(G78gat), .B(G106gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT31), .B(G50gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n448), .A2(new_n449), .ZN(new_n455));
  AOI211_X1 g254(.A(G22gat), .B(new_n437), .C1(new_n444), .C2(new_n447), .ZN(new_n456));
  OAI22_X1  g255(.A1(new_n450), .A2(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n444), .A2(new_n447), .ZN(new_n458));
  INV_X1    g257(.A(new_n437), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(G22gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n448), .A2(new_n449), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n461), .A2(KEYINPUT88), .A3(new_n462), .A4(new_n453), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n381), .A2(new_n261), .ZN(new_n465));
  NAND2_X1  g264(.A1(G227gat), .A2(G233gat), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n229), .A2(new_n363), .A3(new_n373), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(KEYINPUT34), .ZN(new_n469));
  INV_X1    g268(.A(new_n466), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n229), .A2(new_n363), .A3(new_n373), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n229), .B1(new_n373), .B2(new_n363), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT71), .B(G71gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(G99gat), .ZN(new_n475));
  XOR2_X1   g274(.A(G15gat), .B(G43gat), .Z(new_n476));
  XNOR2_X1  g275(.A(new_n475), .B(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT33), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n473), .A2(KEYINPUT32), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT72), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n473), .A2(KEYINPUT72), .A3(KEYINPUT32), .A4(new_n478), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT33), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n473), .B1(KEYINPUT32), .B2(new_n483), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n481), .A2(new_n482), .B1(new_n477), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n469), .B1(new_n485), .B2(KEYINPUT73), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n477), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT32), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n465), .A2(new_n467), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n488), .B1(new_n489), .B2(new_n470), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT72), .B1(new_n490), .B2(new_n478), .ZN(new_n491));
  INV_X1    g290(.A(new_n482), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n487), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT73), .ZN(new_n494));
  INV_X1    g293(.A(new_n469), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n486), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n428), .A2(new_n464), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT35), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n303), .A2(new_n291), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n422), .A2(new_n427), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT35), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n493), .A2(new_n469), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n485), .A2(new_n495), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n506), .B1(new_n457), .B2(new_n463), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT36), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n509), .B1(new_n486), .B2(new_n496), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT36), .B1(new_n504), .B2(new_n505), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n457), .A2(new_n463), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n500), .A2(new_n501), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OR2_X1    g314(.A1(new_n277), .A2(new_n278), .ZN(new_n516));
  OAI211_X1 g315(.A(KEYINPUT39), .B(new_n516), .C1(new_n298), .C2(new_n267), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n289), .A2(new_n271), .ZN(new_n518));
  XOR2_X1   g317(.A(KEYINPUT89), .B(KEYINPUT39), .Z(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n278), .A3(new_n519), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n517), .A2(KEYINPUT40), .A3(new_n205), .A4(new_n520), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n521), .A2(new_n292), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n517), .A2(new_n205), .A3(new_n520), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT40), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n522), .A2(new_n427), .A3(new_n422), .A4(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT90), .B(KEYINPUT38), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(KEYINPUT37), .B1(new_n425), .B2(new_n398), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n411), .A2(new_n324), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT37), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n382), .B1(new_n374), .B2(new_n375), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n395), .B1(new_n532), .B2(new_n389), .ZN(new_n533));
  NOR3_X1   g332(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n419), .B(new_n528), .C1(new_n529), .C2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n535), .A2(new_n291), .A3(new_n303), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n413), .A2(new_n531), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n387), .A2(KEYINPUT37), .A3(new_n398), .A4(new_n412), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n418), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n421), .B1(new_n539), .B2(new_n528), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n464), .B(new_n526), .C1(new_n536), .C2(new_n540), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n499), .A2(new_n508), .B1(new_n515), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(G43gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(G50gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT92), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT15), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(G50gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(G43gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(new_n544), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(new_n549), .ZN(new_n551));
  INV_X1    g350(.A(G29gat), .ZN(new_n552));
  INV_X1    g351(.A(G36gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT14), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT14), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(G29gat), .B2(G36gat), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G29gat), .A2(G36gat), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n550), .A2(new_n551), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n549), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n554), .A2(new_n556), .A3(KEYINPUT91), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n558), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT91), .B1(new_n554), .B2(new_n556), .ZN(new_n563));
  OAI211_X1 g362(.A(KEYINPUT15), .B(new_n560), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(KEYINPUT93), .B(KEYINPUT17), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(G15gat), .B(G22gat), .Z(new_n569));
  INV_X1    g368(.A(G1gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G15gat), .B(G22gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT16), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n572), .B1(new_n573), .B2(G1gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n571), .A2(new_n574), .A3(KEYINPUT94), .ZN(new_n575));
  INV_X1    g374(.A(G8gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n559), .A2(new_n564), .A3(KEYINPUT17), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n568), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n575), .B(G8gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(new_n565), .ZN(new_n581));
  NAND2_X1  g380(.A1(G229gat), .A2(G233gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT18), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n577), .A2(new_n559), .A3(new_n564), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(new_n581), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n582), .B(KEYINPUT13), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n579), .A2(KEYINPUT18), .A3(new_n581), .A4(new_n582), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n585), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(KEYINPUT11), .B(G169gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(G197gat), .ZN(new_n594));
  XOR2_X1   g393(.A(G113gat), .B(G141gat), .Z(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT12), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n592), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n585), .A2(new_n590), .A3(new_n597), .A4(new_n591), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(KEYINPUT95), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT95), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n592), .A2(new_n602), .A3(new_n598), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT96), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n601), .A2(new_n603), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT96), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n542), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G134gat), .B(G162gat), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT101), .ZN(new_n614));
  INV_X1    g413(.A(G85gat), .ZN(new_n615));
  INV_X1    g414(.A(G92gat), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(KEYINPUT101), .A2(G85gat), .A3(G92gat), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n617), .A2(KEYINPUT7), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G99gat), .A2(G106gat), .ZN(new_n620));
  AOI22_X1  g419(.A1(KEYINPUT8), .A2(new_n620), .B1(new_n615), .B2(new_n616), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT7), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n614), .B(new_n622), .C1(new_n615), .C2(new_n616), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n619), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g423(.A(G99gat), .B(G106gat), .Z(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n625), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n627), .A2(new_n621), .A3(new_n619), .A4(new_n623), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G232gat), .A2(G233gat), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n631), .B(KEYINPUT100), .Z(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  AOI22_X1  g432(.A1(new_n630), .A2(new_n565), .B1(KEYINPUT41), .B2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT102), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n568), .A2(new_n629), .A3(new_n578), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n633), .A2(KEYINPUT41), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G190gat), .B(G218gat), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n635), .B(new_n636), .C1(KEYINPUT41), .C2(new_n633), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n639), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n641), .B1(new_n639), .B2(new_n642), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n613), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n645), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n647), .A2(new_n612), .A3(new_n643), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n650));
  XNOR2_X1  g449(.A(G183gat), .B(G211gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT21), .ZN(new_n654));
  INV_X1    g453(.A(G57gat), .ZN(new_n655));
  OR3_X1    g454(.A1(new_n655), .A2(new_n417), .A3(KEYINPUT98), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n417), .B1(new_n655), .B2(KEYINPUT98), .ZN(new_n657));
  INV_X1    g456(.A(G71gat), .ZN(new_n658));
  INV_X1    g457(.A(G78gat), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n658), .A2(new_n659), .A3(KEYINPUT9), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n656), .B(new_n657), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n655), .A2(new_n417), .ZN(new_n663));
  NAND2_X1  g462(.A1(G57gat), .A2(G64gat), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(KEYINPUT9), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n660), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT97), .B1(G71gat), .B2(G78gat), .ZN(new_n667));
  OR3_X1    g466(.A1(KEYINPUT97), .A2(G71gat), .A3(G78gat), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n665), .A2(new_n666), .A3(new_n667), .A4(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n662), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n577), .B1(new_n654), .B2(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT99), .ZN(new_n672));
  AND2_X1   g471(.A1(G231gat), .A2(G233gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n662), .A2(new_n669), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(KEYINPUT21), .ZN(new_n676));
  XOR2_X1   g475(.A(G127gat), .B(G155gat), .Z(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n674), .A2(new_n679), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n653), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n682), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n684), .A2(new_n652), .A3(new_n680), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n649), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n629), .A2(new_n670), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT10), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n675), .A2(new_n626), .A3(new_n628), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n630), .A2(KEYINPUT10), .A3(new_n675), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(new_n692), .A3(KEYINPUT103), .ZN(new_n693));
  NAND2_X1  g492(.A1(G230gat), .A2(G233gat), .ZN(new_n694));
  OR3_X1    g493(.A1(new_n690), .A2(KEYINPUT103), .A3(new_n689), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n688), .A2(new_n690), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n697), .A2(G230gat), .A3(G233gat), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(G120gat), .B(G148gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(new_n338), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(new_n310), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n702), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n696), .A2(new_n698), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n687), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n611), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(new_n500), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(new_n570), .ZN(G1324gat));
  NOR2_X1   g509(.A1(new_n708), .A2(new_n501), .ZN(new_n711));
  NAND2_X1  g510(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n573), .A2(new_n576), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n714), .A2(KEYINPUT42), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(KEYINPUT42), .ZN(new_n716));
  OAI211_X1 g515(.A(new_n715), .B(new_n716), .C1(new_n576), .C2(new_n711), .ZN(G1325gat));
  INV_X1    g516(.A(G15gat), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n485), .A2(KEYINPUT73), .A3(new_n469), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n495), .B1(new_n493), .B2(new_n494), .ZN(new_n720));
  OAI21_X1  g519(.A(KEYINPUT36), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n506), .A2(new_n509), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n708), .A2(new_n718), .A3(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n506), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n611), .A2(new_n707), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n724), .B1(new_n718), .B2(new_n726), .ZN(G1326gat));
  NOR2_X1   g526(.A1(new_n708), .A2(new_n464), .ZN(new_n728));
  XOR2_X1   g527(.A(KEYINPUT43), .B(G22gat), .Z(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1327gat));
  NAND2_X1  g529(.A1(new_n499), .A2(new_n508), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n515), .A2(new_n541), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n649), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n686), .A2(new_n706), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n733), .A2(new_n609), .A3(new_n734), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n303), .A2(new_n291), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n735), .A2(new_n552), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT45), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(new_n542), .B2(new_n649), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n646), .A2(new_n648), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n723), .B1(new_n428), .B2(new_n464), .ZN(new_n742));
  OR2_X1    g541(.A1(new_n536), .A2(new_n540), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n526), .A2(new_n464), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AOI22_X1  g544(.A1(new_n498), .A2(KEYINPUT35), .B1(new_n503), .B2(new_n507), .ZN(new_n746));
  OAI211_X1 g545(.A(KEYINPUT44), .B(new_n741), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n740), .A2(new_n604), .A3(new_n747), .A4(new_n734), .ZN(new_n748));
  OAI21_X1  g547(.A(G29gat), .B1(new_n748), .B2(new_n500), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n738), .A2(new_n749), .ZN(G1328gat));
  INV_X1    g549(.A(new_n501), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n553), .A3(new_n751), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n752), .A2(KEYINPUT104), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(KEYINPUT104), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT46), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(G36gat), .B1(new_n748), .B2(new_n501), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n753), .A2(KEYINPUT46), .A3(new_n754), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(G1329gat));
  OAI21_X1  g559(.A(G43gat), .B1(new_n748), .B2(new_n723), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n735), .A2(new_n543), .A3(new_n725), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT105), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT47), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n763), .B(new_n765), .ZN(G1330gat));
  NOR3_X1   g565(.A1(new_n748), .A2(new_n547), .A3(new_n464), .ZN(new_n767));
  AOI21_X1  g566(.A(G50gat), .B1(new_n735), .B2(new_n513), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n769), .B(KEYINPUT48), .Z(G1331gat));
  INV_X1    g569(.A(new_n541), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n507), .A2(new_n502), .A3(new_n428), .ZN(new_n772));
  AOI22_X1  g571(.A1(new_n457), .A2(new_n463), .B1(new_n496), .B2(new_n486), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n502), .B1(new_n773), .B2(new_n428), .ZN(new_n774));
  OAI22_X1  g573(.A1(new_n771), .A2(new_n742), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n687), .A2(new_n604), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n775), .A2(new_n706), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT106), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n775), .A2(KEYINPUT106), .A3(new_n706), .A4(new_n776), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(new_n500), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(new_n655), .ZN(G1332gat));
  INV_X1    g582(.A(KEYINPUT49), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n751), .B1(new_n784), .B2(new_n417), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT107), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n779), .A2(new_n780), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n784), .A2(new_n417), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n787), .B(new_n788), .ZN(G1333gat));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n779), .A2(new_n725), .A3(new_n780), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n658), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT108), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n779), .A2(G71gat), .A3(new_n512), .A4(new_n780), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n793), .B1(new_n792), .B2(new_n794), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n790), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n792), .A2(new_n794), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT108), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(KEYINPUT50), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n797), .A2(new_n801), .ZN(G1334gat));
  NOR2_X1   g601(.A1(new_n781), .A2(new_n464), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(new_n659), .ZN(G1335gat));
  NOR2_X1   g603(.A1(new_n686), .A2(new_n604), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n733), .A2(new_n805), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n806), .A2(KEYINPUT51), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n806), .A2(KEYINPUT51), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n706), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n736), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n686), .A2(new_n810), .A3(new_n604), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n740), .A2(new_n747), .A3(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n814), .A2(G85gat), .ZN(new_n815));
  AOI22_X1  g614(.A1(new_n812), .A2(new_n615), .B1(new_n815), .B2(new_n736), .ZN(G1336gat));
  NOR2_X1   g615(.A1(new_n501), .A2(G92gat), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n706), .B(new_n817), .C1(new_n807), .C2(new_n808), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n740), .A2(new_n751), .A3(new_n747), .A4(new_n813), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(G92gat), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT109), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n820), .A2(KEYINPUT109), .A3(G92gat), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT110), .B1(KEYINPUT111), .B2(KEYINPUT51), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n827), .B1(new_n733), .B2(new_n805), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT110), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n775), .A2(new_n829), .A3(new_n741), .A4(new_n805), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT111), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n828), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n706), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT112), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT51), .B1(new_n830), .B2(KEYINPUT111), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT112), .ZN(new_n838));
  NOR4_X1   g637(.A1(new_n837), .A2(new_n828), .A3(new_n838), .A4(new_n834), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n826), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n822), .B1(new_n840), .B2(new_n819), .ZN(G1337gat));
  INV_X1    g640(.A(G99gat), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n811), .A2(new_n842), .A3(new_n725), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n814), .A2(new_n512), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n843), .B1(new_n842), .B2(new_n844), .ZN(G1338gat));
  NOR3_X1   g644(.A1(new_n464), .A2(G106gat), .A3(new_n810), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n833), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n740), .A2(new_n513), .A3(new_n747), .A4(new_n813), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(G106gat), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n848), .A2(KEYINPUT113), .A3(G106gat), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n847), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT53), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n846), .B1(new_n807), .B2(new_n808), .ZN(new_n855));
  XNOR2_X1  g654(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n855), .A2(new_n849), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n854), .A2(new_n857), .ZN(G1339gat));
  NOR2_X1   g657(.A1(new_n587), .A2(new_n589), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT115), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n582), .B1(new_n579), .B2(new_n581), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n596), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(new_n706), .A3(new_n600), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT55), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n694), .B1(new_n693), .B2(new_n695), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n702), .B1(new_n696), .B2(KEYINPUT54), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n864), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n869), .ZN(new_n871));
  INV_X1    g670(.A(new_n866), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(KEYINPUT54), .A3(new_n696), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n871), .A2(new_n873), .A3(KEYINPUT55), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n870), .A2(new_n874), .A3(new_n705), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n863), .B1(new_n875), .B2(new_n606), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n863), .B(KEYINPUT116), .C1(new_n875), .C2(new_n606), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n878), .A2(new_n649), .A3(new_n879), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n862), .A2(new_n600), .ZN(new_n881));
  INV_X1    g680(.A(new_n875), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n741), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n686), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n687), .A2(new_n706), .A3(new_n604), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n886), .A2(new_n500), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n773), .A2(new_n501), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XOR2_X1   g688(.A(new_n889), .B(KEYINPUT118), .Z(new_n890));
  NAND3_X1  g689(.A1(new_n890), .A2(new_n216), .A3(new_n604), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n892), .B1(new_n886), .B2(new_n513), .ZN(new_n893));
  OAI211_X1 g692(.A(KEYINPUT117), .B(new_n464), .C1(new_n884), .C2(new_n885), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n895), .A2(new_n736), .A3(new_n501), .A4(new_n725), .ZN(new_n896));
  OAI21_X1  g695(.A(G113gat), .B1(new_n896), .B2(new_n610), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n891), .A2(new_n897), .ZN(G1340gat));
  NAND3_X1  g697(.A1(new_n890), .A2(new_n214), .A3(new_n706), .ZN(new_n899));
  OAI21_X1  g698(.A(G120gat), .B1(new_n896), .B2(new_n810), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(G1341gat));
  INV_X1    g700(.A(new_n889), .ZN(new_n902));
  AOI21_X1  g701(.A(G127gat), .B1(new_n902), .B2(new_n686), .ZN(new_n903));
  INV_X1    g702(.A(new_n686), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n896), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n903), .B1(new_n905), .B2(G127gat), .ZN(G1342gat));
  NOR3_X1   g705(.A1(new_n889), .A2(G134gat), .A3(new_n649), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT56), .ZN(new_n908));
  OAI21_X1  g707(.A(G134gat), .B1(new_n896), .B2(new_n649), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1343gat));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n512), .A2(new_n751), .A3(new_n500), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT119), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n875), .B1(new_n605), .B2(new_n608), .ZN(new_n914));
  INV_X1    g713(.A(new_n863), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n649), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n686), .B1(new_n916), .B2(new_n883), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n513), .B1(new_n917), .B2(new_n885), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n913), .B1(new_n918), .B2(KEYINPUT57), .ZN(new_n919));
  INV_X1    g718(.A(new_n886), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT57), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n920), .A2(new_n921), .A3(new_n513), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n911), .B1(new_n923), .B2(new_n610), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n919), .A2(new_n922), .A3(KEYINPUT122), .A4(new_n609), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n924), .A2(G141gat), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n513), .A2(new_n723), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT121), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n887), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n501), .B1(new_n927), .B2(KEYINPUT121), .ZN(new_n930));
  NOR4_X1   g729(.A1(new_n929), .A2(G141gat), .A3(new_n610), .A4(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n931), .A2(KEYINPUT58), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n926), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT120), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n919), .A2(new_n922), .A3(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n934), .B1(new_n919), .B2(new_n922), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n604), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n931), .B1(new_n938), .B2(G141gat), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT58), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n933), .B1(new_n939), .B2(new_n940), .ZN(G1344gat));
  NOR2_X1   g740(.A1(new_n929), .A2(new_n930), .ZN(new_n942));
  INV_X1    g741(.A(G148gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n942), .A2(new_n943), .A3(new_n706), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n706), .B1(new_n936), .B2(new_n937), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT59), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n945), .A2(new_n946), .A3(G148gat), .ZN(new_n947));
  OAI21_X1  g746(.A(KEYINPUT57), .B1(new_n886), .B2(new_n464), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n687), .A2(new_n706), .A3(new_n609), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n921), .B(new_n513), .C1(new_n917), .C2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  OR3_X1    g750(.A1(new_n951), .A2(new_n810), .A3(new_n913), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n946), .B1(new_n952), .B2(G148gat), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n944), .B1(new_n947), .B2(new_n953), .ZN(G1345gat));
  AOI21_X1  g753(.A(new_n247), .B1(new_n942), .B2(new_n686), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n936), .A2(new_n937), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n956), .A2(new_n904), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n955), .B1(new_n957), .B2(new_n247), .ZN(G1346gat));
  AOI21_X1  g757(.A(new_n248), .B1(new_n942), .B2(new_n741), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n956), .A2(new_n649), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n959), .B1(new_n960), .B2(new_n248), .ZN(G1347gat));
  NOR2_X1   g760(.A1(new_n736), .A2(new_n501), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(new_n725), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n963), .B1(new_n893), .B2(new_n894), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(G169gat), .B1(new_n965), .B2(new_n610), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n920), .A2(new_n773), .A3(new_n962), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n968), .A2(new_n337), .A3(new_n604), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n966), .A2(new_n969), .ZN(G1348gat));
  AOI21_X1  g769(.A(G176gat), .B1(new_n968), .B2(new_n706), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n965), .A2(new_n810), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n971), .B1(new_n972), .B2(G176gat), .ZN(G1349gat));
  NAND2_X1  g772(.A1(new_n964), .A2(new_n686), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(G183gat), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n968), .A2(new_n686), .A3(new_n368), .ZN(new_n976));
  NAND2_X1  g775(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  NOR2_X1   g777(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n979), .B(KEYINPUT124), .ZN(new_n980));
  INV_X1    g779(.A(new_n980), .ZN(new_n981));
  XNOR2_X1  g780(.A(new_n978), .B(new_n981), .ZN(G1350gat));
  NAND3_X1  g781(.A1(new_n968), .A2(new_n369), .A3(new_n741), .ZN(new_n983));
  AOI211_X1 g782(.A(KEYINPUT61), .B(new_n369), .C1(new_n964), .C2(new_n741), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT61), .ZN(new_n985));
  INV_X1    g784(.A(new_n963), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n895), .A2(new_n741), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n985), .B1(new_n987), .B2(G190gat), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n983), .B1(new_n984), .B2(new_n988), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT125), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI211_X1 g790(.A(KEYINPUT125), .B(new_n983), .C1(new_n984), .C2(new_n988), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(new_n992), .ZN(G1351gat));
  NOR3_X1   g792(.A1(new_n512), .A2(new_n736), .A3(new_n501), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n920), .A2(new_n513), .A3(new_n994), .ZN(new_n995));
  INV_X1    g794(.A(new_n995), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n996), .A2(new_n309), .A3(new_n604), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n997), .B(KEYINPUT126), .ZN(new_n998));
  INV_X1    g797(.A(new_n951), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n999), .A2(new_n994), .ZN(new_n1000));
  OAI21_X1  g799(.A(G197gat), .B1(new_n1000), .B2(new_n610), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n998), .A2(new_n1001), .ZN(G1352gat));
  NAND3_X1  g801(.A1(new_n996), .A2(new_n310), .A3(new_n706), .ZN(new_n1003));
  OR3_X1    g802(.A1(new_n1003), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(KEYINPUT62), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n999), .A2(new_n706), .A3(new_n994), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1006), .A2(G204gat), .ZN(new_n1007));
  OAI21_X1  g806(.A(KEYINPUT127), .B1(new_n1003), .B2(KEYINPUT62), .ZN(new_n1008));
  NAND4_X1  g807(.A1(new_n1004), .A2(new_n1005), .A3(new_n1007), .A4(new_n1008), .ZN(G1353gat));
  NAND3_X1  g808(.A1(new_n996), .A2(new_n318), .A3(new_n686), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n999), .A2(new_n686), .A3(new_n994), .ZN(new_n1011));
  AND3_X1   g810(.A1(new_n1011), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1012));
  AOI21_X1  g811(.A(KEYINPUT63), .B1(new_n1011), .B2(G211gat), .ZN(new_n1013));
  OAI21_X1  g812(.A(new_n1010), .B1(new_n1012), .B2(new_n1013), .ZN(G1354gat));
  OAI21_X1  g813(.A(G218gat), .B1(new_n1000), .B2(new_n649), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n996), .A2(new_n319), .A3(new_n741), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1015), .A2(new_n1016), .ZN(G1355gat));
endmodule


