//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT67), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT68), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n452), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT69), .ZN(G319));
  XOR2_X1   g036(.A(KEYINPUT70), .B(G2104), .Z(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(G101), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  OR2_X1    g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(new_n464), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n475), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(new_n464), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT71), .ZN(G160));
  NAND2_X1  g054(.A1(new_n466), .A2(new_n468), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n480), .A2(new_n464), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT72), .Z(new_n487));
  NAND3_X1  g062(.A1(new_n482), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR4_X1   g065(.A1(new_n474), .A2(KEYINPUT4), .A3(new_n490), .A4(G2105), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n469), .A2(G138), .A3(new_n464), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(KEYINPUT4), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G114), .C2(new_n464), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n469), .A2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G126), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OR2_X1    g073(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT75), .B1(new_n503), .B2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT75), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(new_n501), .A3(G543), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n502), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT74), .A2(G651), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT73), .A2(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n516));
  AOI21_X1  g091(.A(KEYINPUT73), .B1(KEYINPUT74), .B2(G651), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n507), .A2(new_n518), .A3(G88), .ZN(new_n519));
  INV_X1    g094(.A(G50), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(G543), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n510), .A2(new_n522), .ZN(G166));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(new_n502), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n505), .B1(new_n501), .B2(G543), .ZN(new_n527));
  NOR3_X1   g102(.A1(new_n503), .A2(KEYINPUT75), .A3(KEYINPUT5), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(G63), .A2(G651), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n525), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n507), .A2(new_n518), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n531), .B1(G89), .B2(new_n533), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n518), .A2(KEYINPUT76), .A3(G543), .ZN(new_n535));
  AOI21_X1  g110(.A(KEYINPUT76), .B1(new_n518), .B2(G543), .ZN(new_n536));
  OAI21_X1  g111(.A(G51), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(G168));
  INV_X1    g113(.A(G52), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT76), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n521), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n518), .A2(KEYINPUT76), .A3(G543), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n539), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n507), .A2(new_n518), .A3(G90), .ZN(new_n544));
  NAND2_X1  g119(.A1(G77), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n546), .B1(new_n507), .B2(G64), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n544), .B1(new_n547), .B2(new_n509), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT77), .ZN(new_n549));
  NOR3_X1   g124(.A1(new_n543), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  OAI211_X1 g125(.A(G64), .B(new_n526), .C1(new_n527), .C2(new_n528), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n509), .B1(new_n551), .B2(new_n545), .ZN(new_n552));
  AND3_X1   g127(.A1(new_n507), .A2(new_n518), .A3(G90), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g129(.A(G52), .B1(new_n535), .B2(new_n536), .ZN(new_n555));
  AOI21_X1  g130(.A(KEYINPUT77), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n550), .A2(new_n556), .ZN(G301));
  INV_X1    g132(.A(G301), .ZN(G171));
  INV_X1    g133(.A(G43), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n559), .B1(new_n541), .B2(new_n542), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G81), .ZN(new_n562));
  OAI22_X1  g137(.A1(new_n561), .A2(new_n509), .B1(new_n562), .B2(new_n532), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  AOI22_X1  g144(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n570), .A2(new_n509), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(G91), .B2(new_n533), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n518), .A2(G53), .A3(G543), .ZN(new_n573));
  AND2_X1   g148(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n572), .A2(new_n576), .ZN(G299));
  NAND2_X1  g152(.A1(new_n534), .A2(new_n537), .ZN(G286));
  OR2_X1    g153(.A1(new_n510), .A2(new_n522), .ZN(G303));
  OAI21_X1  g154(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n507), .A2(new_n518), .A3(G87), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n518), .A2(G49), .A3(G543), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G288));
  NAND3_X1  g158(.A1(new_n518), .A2(G48), .A3(G543), .ZN(new_n584));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n507), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n586));
  OAI221_X1 g161(.A(new_n584), .B1(new_n532), .B2(new_n585), .C1(new_n586), .C2(new_n509), .ZN(G305));
  INV_X1    g162(.A(G47), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(new_n541), .B2(new_n542), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n590), .A2(new_n509), .B1(new_n591), .B2(new_n532), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G290));
  NAND3_X1  g169(.A1(new_n533), .A2(KEYINPUT10), .A3(G92), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n532), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n529), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n595), .A2(new_n598), .B1(G651), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n541), .A2(new_n542), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G54), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n605), .A2(G868), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g182(.A(new_n606), .B1(G171), .B2(G868), .ZN(G321));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n609), .A2(KEYINPUT78), .ZN(new_n610));
  AND2_X1   g185(.A1(new_n609), .A2(KEYINPUT78), .ZN(new_n611));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(G299), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n610), .B1(new_n611), .B2(new_n613), .ZN(G297));
  AOI21_X1  g189(.A(new_n610), .B1(new_n611), .B2(new_n613), .ZN(G280));
  INV_X1    g190(.A(new_n605), .ZN(new_n616));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G860), .ZN(G148));
  OR3_X1    g193(.A1(new_n605), .A2(KEYINPUT79), .A3(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(KEYINPUT79), .B1(new_n605), .B2(G559), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n621), .A2(new_n612), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n622), .B1(new_n612), .B2(new_n564), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n481), .A2(G135), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n483), .A2(G123), .ZN(new_n626));
  OR2_X1    g201(.A1(G99), .A2(G2105), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n627), .B(G2104), .C1(G111), .C2(new_n464), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(G2096), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n475), .A2(new_n463), .A3(new_n464), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT80), .B(G2100), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n632), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n629), .A2(G2096), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n630), .A2(new_n635), .A3(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT82), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2427), .B(G2430), .Z(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n644), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2451), .B(G2454), .Z(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n648), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT83), .Z(G401));
  XOR2_X1   g230(.A(KEYINPUT84), .B(KEYINPUT18), .Z(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g234(.A1(new_n659), .A2(KEYINPUT17), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n657), .A2(new_n658), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n656), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n659), .B2(new_n656), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n662), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2096), .B(G2100), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT85), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1961), .B(G1966), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT20), .Z(new_n676));
  NOR2_X1   g251(.A1(new_n669), .A2(new_n671), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n678), .A2(new_n674), .A3(new_n672), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n676), .B(new_n679), .C1(new_n674), .C2(new_n678), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT86), .ZN(new_n681));
  XOR2_X1   g256(.A(G1981), .B(G1986), .Z(new_n682));
  XNOR2_X1  g257(.A(G1991), .B(G1996), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n681), .B(new_n686), .ZN(G229));
  INV_X1    g262(.A(KEYINPUT101), .ZN(new_n688));
  INV_X1    g263(.A(G29), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G32), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n481), .A2(G141), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT94), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT95), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT26), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n463), .A2(G105), .A3(new_n464), .ZN(new_n697));
  INV_X1    g272(.A(G129), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n696), .B(new_n697), .C1(new_n496), .C2(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n693), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n690), .B1(new_n700), .B2(new_n689), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT96), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT27), .B(G1996), .Z(new_n703));
  OR3_X1    g278(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n702), .B1(new_n701), .B2(new_n703), .ZN(new_n705));
  NAND2_X1  g280(.A1(G160), .A2(G29), .ZN(new_n706));
  INV_X1    g281(.A(G34), .ZN(new_n707));
  AOI21_X1  g282(.A(G29), .B1(new_n707), .B2(KEYINPUT24), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(KEYINPUT24), .B2(new_n707), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  AOI22_X1  g286(.A1(new_n704), .A2(new_n705), .B1(new_n711), .B2(G2084), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT97), .ZN(new_n713));
  OR2_X1    g288(.A1(G29), .A2(G33), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT25), .Z(new_n716));
  INV_X1    g291(.A(G139), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(new_n470), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT93), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n464), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n714), .B1(new_n721), .B2(new_n689), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G2072), .ZN(new_n723));
  AND3_X1   g298(.A1(new_n712), .A2(new_n713), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n713), .B1(new_n712), .B2(new_n723), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n689), .A2(G27), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G164), .B2(new_n689), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT100), .ZN(new_n729));
  INV_X1    g304(.A(G2078), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G16), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G4), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n616), .B2(new_n732), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G1348), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n689), .A2(G26), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT28), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n481), .A2(G140), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n483), .A2(G128), .ZN(new_n740));
  OR2_X1    g315(.A1(G104), .A2(G2105), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n741), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n742));
  AND3_X1   g317(.A1(new_n739), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n738), .B1(new_n743), .B2(new_n689), .ZN(new_n744));
  INV_X1    g319(.A(G2067), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n732), .A2(G21), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G286), .B2(G16), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1966), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n732), .A2(G20), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT23), .ZN(new_n752));
  INV_X1    g327(.A(G299), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(new_n732), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1956), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n689), .A2(G35), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G162), .B2(new_n689), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT29), .B(G2090), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT31), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n760), .A2(G11), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(G11), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT30), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n763), .A2(G28), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n689), .B1(new_n763), .B2(G28), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n761), .B(new_n762), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n629), .A2(new_n689), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(KEYINPUT98), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(KEYINPUT98), .B2(new_n767), .ZN(new_n769));
  NOR4_X1   g344(.A1(new_n750), .A2(new_n755), .A3(new_n759), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n732), .A2(G5), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G171), .B2(new_n732), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n729), .A2(new_n730), .B1(G1961), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(G16), .A2(G19), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n564), .B2(G16), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT92), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(G1341), .Z(new_n777));
  AND4_X1   g352(.A1(new_n736), .A2(new_n770), .A3(new_n773), .A4(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G2084), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n710), .A2(new_n779), .B1(new_n701), .B2(new_n703), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G1961), .B2(new_n772), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT99), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n726), .A2(new_n778), .A3(new_n782), .ZN(new_n783));
  MUX2_X1   g358(.A(G6), .B(G305), .S(G16), .Z(new_n784));
  XOR2_X1   g359(.A(KEYINPUT32), .B(G1981), .Z(new_n785));
  XOR2_X1   g360(.A(new_n784), .B(new_n785), .Z(new_n786));
  NOR2_X1   g361(.A1(G16), .A2(G23), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT89), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G288), .B2(new_n732), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT33), .B(G1976), .Z(new_n790));
  XOR2_X1   g365(.A(new_n789), .B(new_n790), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n732), .A2(G22), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT90), .Z(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G166), .B2(new_n732), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1971), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n786), .A2(new_n791), .A3(new_n795), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT88), .B(KEYINPUT34), .Z(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n481), .A2(G131), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n483), .A2(G119), .ZN(new_n800));
  OR2_X1    g375(.A1(G95), .A2(G2105), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n801), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT87), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n799), .A2(new_n800), .A3(new_n803), .ZN(new_n804));
  MUX2_X1   g379(.A(G25), .B(new_n804), .S(G29), .Z(new_n805));
  XOR2_X1   g380(.A(KEYINPUT35), .B(G1991), .Z(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n805), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n732), .A2(G24), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n593), .B2(new_n732), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(G1986), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n810), .A2(G1986), .ZN(new_n812));
  NOR3_X1   g387(.A1(new_n808), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n796), .A2(new_n797), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n798), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT91), .B(KEYINPUT36), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n815), .B(new_n816), .Z(new_n817));
  OAI21_X1  g392(.A(new_n688), .B1(new_n783), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n782), .A2(new_n778), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n815), .B(new_n816), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n819), .A2(KEYINPUT101), .A3(new_n726), .A4(new_n820), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n818), .A2(new_n821), .ZN(G311));
  NAND3_X1  g397(.A1(new_n819), .A2(new_n726), .A3(new_n820), .ZN(G150));
  NAND2_X1  g398(.A1(new_n616), .A2(G559), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT38), .ZN(new_n825));
  INV_X1    g400(.A(G55), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(new_n541), .B2(new_n542), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n828));
  INV_X1    g403(.A(G93), .ZN(new_n829));
  OAI22_X1  g404(.A1(new_n828), .A2(new_n509), .B1(new_n829), .B2(new_n532), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n564), .A2(new_n831), .ZN(new_n832));
  OAI22_X1  g407(.A1(new_n560), .A2(new_n563), .B1(new_n827), .B2(new_n830), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n825), .B(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT39), .ZN(new_n836));
  AOI21_X1  g411(.A(G860), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n836), .B2(new_n835), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT102), .ZN(new_n839));
  OAI21_X1  g414(.A(G860), .B1(new_n827), .B2(new_n830), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT37), .Z(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n841), .ZN(G145));
  XNOR2_X1  g417(.A(G160), .B(G162), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n629), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n739), .A2(new_n740), .A3(new_n742), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n499), .B(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n721), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n847), .A2(new_n700), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n700), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n481), .A2(G142), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT103), .Z(new_n853));
  INV_X1    g428(.A(KEYINPUT104), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(new_n483), .B2(G130), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n483), .A2(new_n854), .A3(G130), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n464), .A2(G118), .ZN(new_n857));
  OAI21_X1  g432(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n858));
  OAI221_X1 g433(.A(new_n853), .B1(new_n855), .B2(new_n856), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n804), .B(new_n632), .Z(new_n860));
  XOR2_X1   g435(.A(new_n859), .B(new_n860), .Z(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n844), .B1(new_n851), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n849), .A2(new_n861), .A3(new_n850), .ZN(new_n864));
  AOI21_X1  g439(.A(G37), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n850), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n862), .B1(new_n866), .B2(new_n848), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n867), .A2(new_n864), .A3(KEYINPUT105), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT105), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n849), .A2(new_n869), .A3(new_n861), .A4(new_n850), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n844), .A3(new_n870), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n865), .A2(new_n871), .A3(KEYINPUT40), .ZN(new_n872));
  AOI21_X1  g447(.A(KEYINPUT40), .B1(new_n865), .B2(new_n871), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(G395));
  INV_X1    g449(.A(new_n834), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n621), .B(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT41), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n605), .A2(G299), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n605), .A2(G299), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n877), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n616), .A2(new_n753), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n882), .A2(KEYINPUT41), .A3(new_n878), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n876), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n879), .A2(new_n880), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n885), .B1(new_n886), .B2(new_n876), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT106), .ZN(new_n888));
  INV_X1    g463(.A(new_n592), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n603), .A2(G47), .ZN(new_n890));
  INV_X1    g465(.A(G288), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(G288), .B1(new_n589), .B2(new_n592), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n888), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n892), .A2(new_n888), .A3(new_n893), .ZN(new_n896));
  XNOR2_X1  g471(.A(G303), .B(G305), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(G166), .B(G305), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n894), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(KEYINPUT42), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT107), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n902), .B1(new_n898), .B2(new_n900), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n898), .A2(new_n902), .A3(new_n900), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n901), .B1(new_n906), .B2(KEYINPUT42), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n887), .B(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n908), .A2(new_n612), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n831), .A2(G868), .ZN(new_n910));
  OR3_X1    g485(.A1(new_n909), .A2(KEYINPUT108), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT108), .B1(new_n909), .B2(new_n910), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(G295));
  INV_X1    g488(.A(KEYINPUT109), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n908), .A2(new_n612), .ZN(new_n915));
  INV_X1    g490(.A(new_n910), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NOR3_X1   g492(.A1(new_n909), .A2(KEYINPUT109), .A3(new_n910), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(G331));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n920));
  OAI21_X1  g495(.A(G168), .B1(new_n550), .B2(new_n556), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n549), .B1(new_n543), .B2(new_n548), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n554), .A2(new_n555), .A3(KEYINPUT77), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(G286), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n875), .A2(new_n921), .A3(new_n924), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n925), .A2(new_n886), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n922), .A2(G286), .A3(new_n923), .ZN(new_n927));
  AOI21_X1  g502(.A(G286), .B1(new_n922), .B2(new_n923), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n834), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n905), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n931), .A2(new_n903), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT111), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n921), .A2(new_n924), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n934), .A2(new_n834), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n929), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n934), .A2(KEYINPUT110), .A3(new_n834), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n933), .B1(new_n939), .B2(new_n884), .ZN(new_n940));
  AOI221_X4 g515(.A(new_n936), .B1(new_n832), .B2(new_n833), .C1(new_n921), .C2(new_n924), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT110), .B1(new_n934), .B2(new_n834), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n925), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n881), .A2(new_n883), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(KEYINPUT111), .A3(new_n944), .ZN(new_n945));
  AOI211_X1 g520(.A(new_n930), .B(new_n932), .C1(new_n940), .C2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n947));
  INV_X1    g522(.A(G37), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n930), .B1(new_n940), .B2(new_n945), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n948), .B1(new_n949), .B2(new_n906), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n920), .B1(new_n947), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT113), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n949), .A2(new_n906), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n926), .B1(new_n942), .B2(new_n941), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n925), .A2(new_n929), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n955), .B1(new_n884), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(G37), .B1(new_n957), .B2(new_n932), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n953), .B1(new_n959), .B2(KEYINPUT43), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n961));
  AOI211_X1 g536(.A(KEYINPUT113), .B(new_n961), .C1(new_n954), .C2(new_n958), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n952), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT112), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT43), .B1(new_n950), .B2(new_n946), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n954), .A2(new_n958), .A3(new_n961), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n964), .B1(new_n967), .B2(new_n920), .ZN(new_n968));
  AOI211_X1 g543(.A(KEYINPUT112), .B(KEYINPUT44), .C1(new_n965), .C2(new_n966), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n963), .B1(new_n968), .B2(new_n969), .ZN(G397));
  INV_X1    g545(.A(G1384), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n971), .B1(new_n493), .B2(new_n498), .ZN(new_n972));
  INV_X1    g547(.A(G40), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n472), .A2(new_n973), .A3(new_n477), .ZN(new_n974));
  XOR2_X1   g549(.A(KEYINPUT114), .B(KEYINPUT45), .Z(new_n975));
  NAND3_X1  g550(.A1(new_n972), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  OR2_X1    g551(.A1(new_n976), .A2(G1996), .ZN(new_n977));
  INV_X1    g552(.A(new_n700), .ZN(new_n978));
  OR2_X1    g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n976), .A2(G1986), .A3(G290), .ZN(new_n980));
  INV_X1    g555(.A(new_n976), .ZN(new_n981));
  AND2_X1   g556(.A1(G290), .A2(G1986), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  XOR2_X1   g558(.A(new_n983), .B(KEYINPUT115), .Z(new_n984));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n845), .A2(G2067), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT116), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n981), .B1(new_n988), .B2(new_n978), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n988), .A2(G1996), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n804), .B(new_n806), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n992), .B(KEYINPUT117), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n981), .ZN(new_n994));
  AND4_X1   g569(.A1(new_n979), .A2(new_n984), .A3(new_n991), .A4(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n465), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n996), .B1(new_n481), .B2(G137), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n997), .B(G40), .C1(new_n464), .C2(new_n476), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n998), .B1(new_n972), .B2(KEYINPUT50), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT50), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n1000), .B(new_n971), .C1(new_n493), .C2(new_n498), .ZN(new_n1001));
  AOI21_X1  g576(.A(G1961), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n998), .B1(new_n972), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1005), .A2(G2078), .ZN(new_n1006));
  INV_X1    g581(.A(new_n975), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n971), .B(new_n1007), .C1(new_n493), .C2(new_n498), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n1004), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n972), .A2(new_n975), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT118), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g587(.A(KEYINPUT45), .B(new_n971), .C1(new_n493), .C2(new_n498), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n1013), .A2(new_n974), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n972), .A2(KEYINPUT118), .A3(new_n975), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1012), .A2(new_n1014), .A3(new_n730), .A4(new_n1015), .ZN(new_n1016));
  AOI211_X1 g591(.A(new_n1002), .B(new_n1009), .C1(new_n1005), .C2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT124), .B1(new_n1017), .B2(G301), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT124), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1016), .A2(new_n1005), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n972), .A2(KEYINPUT50), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n1021), .A2(new_n974), .A3(new_n1001), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1020), .B1(G1961), .B2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1019), .B(G171), .C1(new_n1023), .C2(new_n1009), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n997), .A2(G40), .A3(new_n1006), .ZN(new_n1025));
  INV_X1    g600(.A(new_n476), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1026), .A2(KEYINPUT125), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n464), .B1(new_n1026), .B2(KEYINPUT125), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n1010), .A2(new_n1029), .A3(new_n1013), .ZN(new_n1030));
  AOI211_X1 g605(.A(new_n1030), .B(new_n1002), .C1(new_n1016), .C2(new_n1005), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT54), .B1(new_n1031), .B2(G301), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1018), .A2(new_n1024), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(G171), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1034), .B(KEYINPUT54), .C1(G171), .C2(new_n1017), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(G8), .B1(new_n972), .B2(new_n998), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT121), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT121), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1039), .B(G8), .C1(new_n972), .C2(new_n998), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n891), .A2(G1976), .ZN(new_n1042));
  INV_X1    g617(.A(G1976), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT52), .B1(G288), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g620(.A(G305), .B(G1981), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1046), .B(KEYINPUT49), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1041), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  AOI22_X1  g624(.A1(new_n1038), .A2(new_n1040), .B1(G1976), .B2(new_n891), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G8), .ZN(new_n1054));
  NOR2_X1   g629(.A1(G166), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT55), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT119), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1055), .A2(new_n1058), .A3(KEYINPUT55), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1057), .A2(KEYINPUT120), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT120), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1055), .A2(KEYINPUT55), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1064));
  INV_X1    g639(.A(G1971), .ZN(new_n1065));
  INV_X1    g640(.A(G2090), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1064), .A2(new_n1065), .B1(new_n1022), .B2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1060), .B(new_n1063), .C1(new_n1067), .C2(new_n1054), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1063), .A2(new_n1060), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1015), .A2(new_n974), .A3(new_n1013), .ZN(new_n1070));
  AOI21_X1  g645(.A(G1971), .B1(new_n1070), .B2(new_n1012), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1021), .A2(new_n974), .A3(new_n1001), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1072), .A2(G2090), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1069), .B(G8), .C1(new_n1071), .C2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1053), .A2(new_n1068), .A3(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1072), .A2(G2084), .ZN(new_n1076));
  AOI21_X1  g651(.A(G1966), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1077));
  OAI21_X1  g652(.A(G286), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n972), .A2(new_n1003), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1079), .A2(new_n974), .A3(new_n1008), .ZN(new_n1080));
  INV_X1    g655(.A(G1966), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1082), .B(G168), .C1(G2084), .C2(new_n1072), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1078), .A2(new_n1083), .A3(G8), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT51), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1022), .A2(new_n779), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1054), .B1(new_n1086), .B2(G168), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT51), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1075), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT57), .B1(new_n576), .B2(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n753), .B(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT56), .B(G2072), .Z(new_n1095));
  XNOR2_X1  g670(.A(new_n1095), .B(KEYINPUT123), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .A4(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G1956), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1072), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1094), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G1348), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n972), .A2(new_n998), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1072), .A2(new_n1101), .B1(new_n745), .B2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(new_n605), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1097), .A2(new_n1094), .A3(new_n1099), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1100), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT58), .B(G1341), .ZN(new_n1107));
  OAI22_X1  g682(.A1(new_n1064), .A2(G1996), .B1(new_n1102), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n564), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n972), .A2(new_n998), .A3(G2067), .ZN(new_n1112));
  AOI211_X1 g687(.A(new_n616), .B(new_n1112), .C1(new_n1072), .C2(new_n1101), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT60), .B1(new_n1104), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT60), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1103), .A2(new_n1115), .A3(new_n616), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1108), .A2(KEYINPUT59), .A3(new_n564), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1111), .A2(new_n1114), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1100), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1119), .A2(KEYINPUT61), .A3(new_n1105), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT61), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1105), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1121), .B1(new_n1122), .B2(new_n1100), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1106), .B1(new_n1118), .B2(new_n1124), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1036), .A2(new_n1090), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1088), .B1(new_n1087), .B2(new_n1078), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1083), .A2(new_n1088), .A3(G8), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT62), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1018), .A2(new_n1024), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1052), .ZN(new_n1132));
  AND4_X1   g707(.A1(new_n1068), .A2(new_n1074), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT62), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1085), .A2(new_n1134), .A3(new_n1089), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1129), .A2(new_n1130), .A3(new_n1133), .A4(new_n1135), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1086), .A2(new_n1054), .A3(G286), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1053), .A2(new_n1068), .A3(new_n1074), .A4(new_n1137), .ZN(new_n1138));
  OR2_X1    g713(.A1(new_n1138), .A2(KEYINPUT63), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n891), .A2(new_n1043), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1140), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1141));
  NOR2_X1   g716(.A1(G305), .A2(G1981), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1041), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1045), .B(new_n1048), .C1(new_n1051), .C2(new_n1050), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1143), .B1(new_n1144), .B2(new_n1074), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1145), .B1(new_n1138), .B2(KEYINPUT63), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1136), .A2(new_n1139), .A3(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n995), .B1(new_n1126), .B2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n804), .A2(new_n807), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n991), .A2(new_n979), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n985), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n981), .ZN(new_n1152));
  XOR2_X1   g727(.A(new_n980), .B(KEYINPUT48), .Z(new_n1153));
  NAND4_X1  g728(.A1(new_n991), .A2(new_n979), .A3(new_n994), .A4(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n977), .B(KEYINPUT46), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n989), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1156), .A2(KEYINPUT47), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1156), .A2(KEYINPUT47), .ZN(new_n1158));
  OR2_X1    g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1152), .A2(KEYINPUT126), .A3(new_n1154), .A4(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT126), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1154), .B1(new_n1158), .B2(new_n1157), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n976), .B1(new_n1150), .B2(new_n985), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1160), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1148), .A2(new_n1165), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g741(.A1(new_n865), .A2(new_n871), .ZN(new_n1168));
  INV_X1    g742(.A(new_n654), .ZN(new_n1169));
  OR2_X1    g743(.A1(G227), .A2(new_n460), .ZN(new_n1170));
  NOR3_X1   g744(.A1(G229), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  XOR2_X1   g745(.A(new_n1171), .B(KEYINPUT127), .Z(new_n1172));
  NAND3_X1  g746(.A1(new_n1168), .A2(new_n1172), .A3(new_n967), .ZN(G225));
  INV_X1    g747(.A(G225), .ZN(G308));
endmodule


