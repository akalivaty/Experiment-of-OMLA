

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753;

  AND2_X1 U376 ( .A1(n533), .A2(n695), .ZN(n534) );
  INV_X2 U377 ( .A(G953), .ZN(n485) );
  XOR2_X1 U378 ( .A(KEYINPUT111), .B(KEYINPUT42), .Z(n354) );
  XOR2_X1 U379 ( .A(KEYINPUT74), .B(G110), .Z(n355) );
  XNOR2_X2 U380 ( .A(n514), .B(n513), .ZN(n560) );
  XNOR2_X2 U381 ( .A(G146), .B(G125), .ZN(n483) );
  XNOR2_X2 U382 ( .A(n484), .B(G134), .ZN(n447) );
  XNOR2_X2 U383 ( .A(n390), .B(G143), .ZN(n484) );
  NAND2_X2 U384 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X2 U385 ( .A(n522), .B(n368), .ZN(n586) );
  NAND2_X2 U386 ( .A1(n520), .A2(n401), .ZN(n522) );
  INV_X1 U387 ( .A(n525), .ZN(n697) );
  NOR2_X1 U388 ( .A1(n531), .A2(n698), .ZN(n532) );
  XNOR2_X1 U389 ( .A(n356), .B(n354), .ZN(n550) );
  OR2_X1 U390 ( .A1(n707), .A2(n566), .ZN(n356) );
  XNOR2_X1 U391 ( .A(n532), .B(KEYINPUT68), .ZN(n695) );
  NOR2_X2 U392 ( .A1(G902), .A2(n662), .ZN(n409) );
  INV_X1 U393 ( .A(G128), .ZN(n390) );
  INV_X1 U394 ( .A(G469), .ZN(n407) );
  INV_X1 U395 ( .A(KEYINPUT34), .ZN(n358) );
  NAND2_X1 U396 ( .A1(n624), .A2(n623), .ZN(n626) );
  NOR2_X2 U397 ( .A1(n629), .A2(n628), .ZN(n691) );
  INV_X1 U398 ( .A(n550), .ZN(n549) );
  AND2_X1 U399 ( .A1(n377), .A2(n375), .ZN(n374) );
  XNOR2_X1 U400 ( .A(n359), .B(n358), .ZN(n589) );
  OR2_X1 U401 ( .A1(n584), .A2(n583), .ZN(n585) );
  AND2_X1 U402 ( .A1(n379), .A2(n376), .ZN(n373) );
  AND2_X1 U403 ( .A1(n504), .A2(n715), .ZN(n716) );
  XNOR2_X1 U404 ( .A(n507), .B(n506), .ZN(n707) );
  XNOR2_X1 U405 ( .A(n391), .B(KEYINPUT109), .ZN(n504) );
  XNOR2_X1 U406 ( .A(n501), .B(n392), .ZN(n711) );
  INV_X1 U407 ( .A(n499), .ZN(n357) );
  XNOR2_X1 U408 ( .A(n447), .B(n432), .ZN(n740) );
  XNOR2_X1 U409 ( .A(n732), .B(n418), .ZN(n491) );
  XNOR2_X1 U410 ( .A(n355), .B(n402), .ZN(n732) );
  XNOR2_X1 U411 ( .A(G119), .B(G116), .ZN(n411) );
  XNOR2_X1 U412 ( .A(G104), .B(G107), .ZN(n402) );
  NAND2_X1 U413 ( .A1(n501), .A2(n710), .ZN(n514) );
  XNOR2_X2 U414 ( .A(n500), .B(n357), .ZN(n501) );
  NAND2_X1 U415 ( .A1(n686), .A2(n586), .ZN(n359) );
  XNOR2_X2 U416 ( .A(n585), .B(KEYINPUT33), .ZN(n686) );
  OR2_X1 U417 ( .A1(n389), .A2(n682), .ZN(n572) );
  NAND2_X1 U418 ( .A1(n711), .A2(n710), .ZN(n391) );
  INV_X1 U419 ( .A(KEYINPUT8), .ZN(n445) );
  XNOR2_X1 U420 ( .A(G116), .B(G107), .ZN(n443) );
  INV_X1 U421 ( .A(KEYINPUT64), .ZN(n625) );
  XNOR2_X1 U422 ( .A(n385), .B(KEYINPUT85), .ZN(n628) );
  NAND2_X1 U423 ( .A1(n388), .A2(n387), .ZN(n561) );
  NOR2_X1 U424 ( .A1(n508), .A2(n679), .ZN(n387) );
  XNOR2_X1 U425 ( .A(n452), .B(n451), .ZN(n538) );
  NAND2_X1 U426 ( .A1(n586), .A2(n365), .ZN(n524) );
  NAND2_X1 U427 ( .A1(n651), .A2(n596), .ZN(n609) );
  XNOR2_X1 U428 ( .A(KEYINPUT4), .B(G101), .ZN(n418) );
  INV_X1 U429 ( .A(KEYINPUT38), .ZN(n392) );
  XNOR2_X1 U430 ( .A(G128), .B(G110), .ZN(n456) );
  XNOR2_X1 U431 ( .A(n483), .B(KEYINPUT10), .ZN(n461) );
  XNOR2_X1 U432 ( .A(G113), .B(G104), .ZN(n428) );
  XNOR2_X1 U433 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n487) );
  BUF_X1 U434 ( .A(n692), .Z(n747) );
  AND2_X1 U435 ( .A1(n593), .A2(n583), .ZN(n379) );
  OR2_X1 U436 ( .A1(n379), .A2(n376), .ZN(n375) );
  XNOR2_X1 U437 ( .A(n382), .B(KEYINPUT75), .ZN(n558) );
  AND2_X1 U438 ( .A1(n695), .A2(n366), .ZN(n384) );
  XNOR2_X1 U439 ( .A(n543), .B(n369), .ZN(n383) );
  XNOR2_X1 U440 ( .A(n560), .B(n371), .ZN(n565) );
  INV_X1 U441 ( .A(KEYINPUT19), .ZN(n371) );
  XNOR2_X1 U442 ( .A(n439), .B(n438), .ZN(n554) );
  XNOR2_X1 U443 ( .A(n437), .B(G475), .ZN(n438) );
  INV_X1 U444 ( .A(G472), .ZN(n399) );
  XNOR2_X1 U445 ( .A(n448), .B(n447), .ZN(n449) );
  NOR2_X1 U446 ( .A1(n691), .A2(n400), .ZN(n393) );
  INV_X1 U447 ( .A(G475), .ZN(n400) );
  NOR2_X1 U448 ( .A1(n691), .A2(n398), .ZN(n397) );
  NOR2_X1 U449 ( .A1(n485), .A2(G952), .ZN(n666) );
  AND2_X1 U450 ( .A1(n563), .A2(n694), .ZN(n682) );
  AND2_X1 U451 ( .A1(n528), .A2(n583), .ZN(n594) );
  NAND2_X1 U452 ( .A1(n380), .A2(n364), .ZN(n726) );
  NAND2_X1 U453 ( .A1(n360), .A2(n381), .ZN(n380) );
  XNOR2_X1 U454 ( .A(n551), .B(G131), .ZN(G33) );
  XOR2_X1 U455 ( .A(n693), .B(KEYINPUT83), .Z(n360) );
  OR2_X1 U456 ( .A1(n688), .A2(G953), .ZN(n361) );
  AND2_X1 U457 ( .A1(n695), .A2(n541), .ZN(n362) );
  OR2_X1 U458 ( .A1(n567), .A2(n680), .ZN(n363) );
  NOR2_X1 U459 ( .A1(n725), .A2(n361), .ZN(n364) );
  AND2_X1 U460 ( .A1(n503), .A2(n530), .ZN(n365) );
  AND2_X1 U461 ( .A1(n541), .A2(n544), .ZN(n366) );
  AND2_X1 U462 ( .A1(n362), .A2(n599), .ZN(n367) );
  XOR2_X1 U463 ( .A(n521), .B(KEYINPUT0), .Z(n368) );
  XNOR2_X1 U464 ( .A(KEYINPUT30), .B(KEYINPUT107), .ZN(n369) );
  INV_X1 U465 ( .A(KEYINPUT2), .ZN(n386) );
  AND2_X1 U466 ( .A1(n586), .A2(n370), .ZN(n536) );
  INV_X1 U467 ( .A(n705), .ZN(n370) );
  NAND2_X1 U468 ( .A1(n586), .A2(n367), .ZN(n671) );
  INV_X1 U469 ( .A(n565), .ZN(n520) );
  NAND2_X1 U470 ( .A1(n374), .A2(n372), .ZN(n651) );
  NAND2_X1 U471 ( .A1(n528), .A2(n373), .ZN(n372) );
  INV_X1 U472 ( .A(n595), .ZN(n376) );
  NAND2_X1 U473 ( .A1(n378), .A2(n595), .ZN(n377) );
  INV_X1 U474 ( .A(n528), .ZN(n378) );
  NOR2_X1 U475 ( .A1(n690), .A2(n691), .ZN(n381) );
  XNOR2_X2 U476 ( .A(n548), .B(KEYINPUT40), .ZN(n551) );
  NAND2_X1 U477 ( .A1(n384), .A2(n383), .ZN(n382) );
  NOR2_X1 U478 ( .A1(n627), .A2(n386), .ZN(n385) );
  NOR2_X1 U479 ( .A1(n561), .A2(n560), .ZN(n562) );
  INV_X1 U480 ( .A(n583), .ZN(n388) );
  NAND2_X1 U481 ( .A1(n363), .A2(n753), .ZN(n389) );
  INV_X1 U482 ( .A(n501), .ZN(n556) );
  NAND2_X1 U483 ( .A1(n394), .A2(n393), .ZN(n639) );
  INV_X1 U484 ( .A(n630), .ZN(n394) );
  NOR2_X2 U485 ( .A1(n630), .A2(n691), .ZN(n661) );
  NAND2_X1 U486 ( .A1(n396), .A2(n395), .ZN(n633) );
  INV_X1 U487 ( .A(n630), .ZN(n395) );
  NOR2_X1 U488 ( .A1(n691), .A2(n399), .ZN(n396) );
  NAND2_X1 U489 ( .A1(n394), .A2(n397), .ZN(n648) );
  INV_X1 U490 ( .A(G210), .ZN(n398) );
  OR2_X1 U491 ( .A1(n519), .A2(n518), .ZN(n401) );
  XNOR2_X1 U492 ( .A(n446), .B(n445), .ZN(n453) );
  NAND2_X1 U493 ( .A1(n453), .A2(G221), .ZN(n455) );
  XNOR2_X1 U494 ( .A(n407), .B(KEYINPUT70), .ZN(n408) );
  XNOR2_X1 U495 ( .A(n450), .B(n449), .ZN(n657) );
  XOR2_X1 U496 ( .A(KEYINPUT69), .B(G131), .Z(n432) );
  XNOR2_X1 U497 ( .A(n740), .B(G146), .ZN(n423) );
  XOR2_X1 U498 ( .A(G137), .B(G140), .Z(n460) );
  XOR2_X1 U499 ( .A(n460), .B(KEYINPUT95), .Z(n404) );
  NAND2_X1 U500 ( .A1(G227), .A2(n485), .ZN(n403) );
  XNOR2_X1 U501 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U502 ( .A(n491), .B(n405), .ZN(n406) );
  XNOR2_X1 U503 ( .A(n423), .B(n406), .ZN(n662) );
  XNOR2_X2 U504 ( .A(n409), .B(n408), .ZN(n541) );
  XNOR2_X1 U505 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n410) );
  XNOR2_X1 U506 ( .A(n541), .B(n410), .ZN(n533) );
  BUF_X1 U507 ( .A(n533), .Z(n694) );
  XNOR2_X1 U508 ( .A(n411), .B(KEYINPUT3), .ZN(n413) );
  XNOR2_X1 U509 ( .A(G113), .B(KEYINPUT71), .ZN(n412) );
  XNOR2_X1 U510 ( .A(n413), .B(n412), .ZN(n493) );
  XOR2_X1 U511 ( .A(KEYINPUT5), .B(KEYINPUT98), .Z(n415) );
  NOR2_X1 U512 ( .A1(G953), .A2(G237), .ZN(n425) );
  NAND2_X1 U513 ( .A1(n425), .A2(G210), .ZN(n414) );
  XNOR2_X1 U514 ( .A(n415), .B(n414), .ZN(n420) );
  INV_X1 U515 ( .A(KEYINPUT97), .ZN(n416) );
  XNOR2_X1 U516 ( .A(n416), .B(G137), .ZN(n417) );
  XNOR2_X1 U517 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U518 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U519 ( .A(n493), .B(n421), .ZN(n422) );
  XNOR2_X1 U520 ( .A(n423), .B(n422), .ZN(n631) );
  INV_X1 U521 ( .A(G902), .ZN(n477) );
  NAND2_X1 U522 ( .A1(n631), .A2(n477), .ZN(n424) );
  XNOR2_X2 U523 ( .A(n424), .B(G472), .ZN(n542) );
  XNOR2_X1 U524 ( .A(n542), .B(KEYINPUT6), .ZN(n583) );
  NAND2_X1 U525 ( .A1(G214), .A2(n425), .ZN(n427) );
  XOR2_X1 U526 ( .A(KEYINPUT11), .B(G122), .Z(n426) );
  XNOR2_X1 U527 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U528 ( .A(KEYINPUT101), .B(KEYINPUT12), .Z(n429) );
  XNOR2_X1 U529 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U530 ( .A(n431), .B(n430), .Z(n434) );
  XNOR2_X1 U531 ( .A(n432), .B(G143), .ZN(n433) );
  XNOR2_X1 U532 ( .A(n434), .B(n433), .ZN(n436) );
  XOR2_X1 U533 ( .A(G140), .B(n461), .Z(n435) );
  XNOR2_X1 U534 ( .A(n436), .B(n435), .ZN(n637) );
  NOR2_X1 U535 ( .A1(G902), .A2(n637), .ZN(n439) );
  XNOR2_X1 U536 ( .A(KEYINPUT102), .B(KEYINPUT13), .ZN(n437) );
  XOR2_X1 U537 ( .A(KEYINPUT7), .B(KEYINPUT103), .Z(n441) );
  XNOR2_X1 U538 ( .A(G122), .B(KEYINPUT104), .ZN(n440) );
  XNOR2_X1 U539 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U540 ( .A(n442), .B(KEYINPUT9), .Z(n444) );
  XNOR2_X1 U541 ( .A(n444), .B(n443), .ZN(n450) );
  NAND2_X1 U542 ( .A1(G234), .A2(n485), .ZN(n446) );
  AND2_X1 U543 ( .A1(G217), .A2(n453), .ZN(n448) );
  NAND2_X1 U544 ( .A1(n657), .A2(n477), .ZN(n452) );
  INV_X1 U545 ( .A(G478), .ZN(n451) );
  NAND2_X1 U546 ( .A1(n554), .A2(n538), .ZN(n679) );
  XOR2_X1 U547 ( .A(G119), .B(KEYINPUT96), .Z(n454) );
  XNOR2_X1 U548 ( .A(n455), .B(n454), .ZN(n459) );
  XOR2_X1 U549 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n457) );
  XOR2_X1 U550 ( .A(n457), .B(n456), .Z(n458) );
  XNOR2_X1 U551 ( .A(n459), .B(n458), .ZN(n462) );
  XOR2_X1 U552 ( .A(n461), .B(n460), .Z(n739) );
  XNOR2_X1 U553 ( .A(n462), .B(n739), .ZN(n655) );
  NAND2_X1 U554 ( .A1(n655), .A2(n477), .ZN(n467) );
  XOR2_X1 U555 ( .A(KEYINPUT25), .B(KEYINPUT76), .Z(n465) );
  XNOR2_X1 U556 ( .A(G902), .B(KEYINPUT15), .ZN(n620) );
  NAND2_X1 U557 ( .A1(n620), .A2(G234), .ZN(n463) );
  XNOR2_X1 U558 ( .A(n463), .B(KEYINPUT20), .ZN(n473) );
  AND2_X1 U559 ( .A1(n473), .A2(G217), .ZN(n464) );
  XNOR2_X1 U560 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U561 ( .A(n467), .B(n466), .ZN(n531) );
  INV_X1 U562 ( .A(n531), .ZN(n525) );
  NAND2_X1 U563 ( .A1(G234), .A2(G237), .ZN(n468) );
  XNOR2_X1 U564 ( .A(n468), .B(KEYINPUT14), .ZN(n469) );
  NAND2_X1 U565 ( .A1(G952), .A2(n469), .ZN(n724) );
  NOR2_X1 U566 ( .A1(n724), .A2(G953), .ZN(n518) );
  NAND2_X1 U567 ( .A1(G902), .A2(n469), .ZN(n516) );
  OR2_X1 U568 ( .A1(n485), .A2(n516), .ZN(n470) );
  NOR2_X1 U569 ( .A1(G900), .A2(n470), .ZN(n471) );
  NOR2_X1 U570 ( .A1(n518), .A2(n471), .ZN(n472) );
  XOR2_X1 U571 ( .A(KEYINPUT80), .B(n472), .Z(n544) );
  AND2_X1 U572 ( .A1(n697), .A2(n544), .ZN(n475) );
  AND2_X1 U573 ( .A1(n473), .A2(G221), .ZN(n474) );
  XNOR2_X1 U574 ( .A(n474), .B(KEYINPUT21), .ZN(n530) );
  NAND2_X1 U575 ( .A1(n475), .A2(n530), .ZN(n508) );
  INV_X1 U576 ( .A(n561), .ZN(n478) );
  INV_X1 U577 ( .A(G237), .ZN(n476) );
  NAND2_X1 U578 ( .A1(n477), .A2(n476), .ZN(n495) );
  NAND2_X1 U579 ( .A1(n495), .A2(G214), .ZN(n710) );
  NAND2_X1 U580 ( .A1(n478), .A2(n710), .ZN(n479) );
  OR2_X1 U581 ( .A1(n694), .A2(n479), .ZN(n482) );
  XOR2_X1 U582 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n480) );
  XNOR2_X1 U583 ( .A(KEYINPUT105), .B(n480), .ZN(n481) );
  XNOR2_X1 U584 ( .A(n482), .B(n481), .ZN(n502) );
  XNOR2_X1 U585 ( .A(n484), .B(n483), .ZN(n489) );
  NAND2_X1 U586 ( .A1(n485), .A2(G224), .ZN(n486) );
  XNOR2_X1 U587 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U588 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U589 ( .A(n491), .B(n490), .ZN(n494) );
  XNOR2_X1 U590 ( .A(KEYINPUT16), .B(G122), .ZN(n492) );
  XNOR2_X1 U591 ( .A(n493), .B(n492), .ZN(n733) );
  XNOR2_X1 U592 ( .A(n494), .B(n733), .ZN(n642) );
  NAND2_X1 U593 ( .A1(n642), .A2(n620), .ZN(n500) );
  NAND2_X1 U594 ( .A1(n495), .A2(G210), .ZN(n496) );
  XNOR2_X1 U595 ( .A(n496), .B(KEYINPUT92), .ZN(n498) );
  XNOR2_X1 U596 ( .A(KEYINPUT79), .B(KEYINPUT91), .ZN(n497) );
  XNOR2_X1 U597 ( .A(n498), .B(n497), .ZN(n499) );
  NAND2_X1 U598 ( .A1(n502), .A2(n556), .ZN(n579) );
  XNOR2_X1 U599 ( .A(n579), .B(G140), .ZN(G42) );
  INV_X1 U600 ( .A(n538), .ZN(n555) );
  OR2_X1 U601 ( .A1(n554), .A2(n555), .ZN(n712) );
  INV_X1 U602 ( .A(n712), .ZN(n503) );
  NAND2_X1 U603 ( .A1(n504), .A2(n503), .ZN(n507) );
  INV_X1 U604 ( .A(KEYINPUT110), .ZN(n505) );
  XNOR2_X1 U605 ( .A(n505), .B(KEYINPUT41), .ZN(n506) );
  INV_X1 U606 ( .A(n508), .ZN(n509) );
  NAND2_X1 U607 ( .A1(n509), .A2(n542), .ZN(n511) );
  INV_X1 U608 ( .A(KEYINPUT28), .ZN(n510) );
  XNOR2_X1 U609 ( .A(n511), .B(n510), .ZN(n512) );
  NAND2_X1 U610 ( .A1(n512), .A2(n541), .ZN(n566) );
  XOR2_X1 U611 ( .A(n549), .B(G137), .Z(G39) );
  INV_X1 U612 ( .A(KEYINPUT87), .ZN(n513) );
  NOR2_X1 U613 ( .A1(G898), .A2(n485), .ZN(n515) );
  XNOR2_X1 U614 ( .A(KEYINPUT93), .B(n515), .ZN(n735) );
  NOR2_X1 U615 ( .A1(n516), .A2(n735), .ZN(n517) );
  XNOR2_X1 U616 ( .A(n517), .B(KEYINPUT94), .ZN(n519) );
  INV_X1 U617 ( .A(KEYINPUT89), .ZN(n521) );
  INV_X1 U618 ( .A(KEYINPUT22), .ZN(n523) );
  XNOR2_X2 U619 ( .A(n524), .B(n523), .ZN(n528) );
  OR2_X1 U620 ( .A1(n542), .A2(n525), .ZN(n526) );
  NOR2_X1 U621 ( .A1(n694), .A2(n526), .ZN(n527) );
  NAND2_X1 U622 ( .A1(n528), .A2(n527), .ZN(n596) );
  XNOR2_X1 U623 ( .A(n596), .B(G110), .ZN(G12) );
  NOR2_X1 U624 ( .A1(n694), .A2(n697), .ZN(n529) );
  NAND2_X1 U625 ( .A1(n594), .A2(n529), .ZN(n605) );
  XNOR2_X1 U626 ( .A(n605), .B(G101), .ZN(G3) );
  INV_X1 U627 ( .A(n530), .ZN(n698) );
  XNOR2_X1 U628 ( .A(n534), .B(KEYINPUT73), .ZN(n584) );
  INV_X1 U629 ( .A(n542), .ZN(n599) );
  OR2_X1 U630 ( .A1(n584), .A2(n599), .ZN(n705) );
  XNOR2_X1 U631 ( .A(KEYINPUT99), .B(KEYINPUT31), .ZN(n535) );
  XNOR2_X1 U632 ( .A(n536), .B(n535), .ZN(n601) );
  INV_X1 U633 ( .A(n679), .ZN(n547) );
  NAND2_X1 U634 ( .A1(n601), .A2(n547), .ZN(n537) );
  XNOR2_X1 U635 ( .A(n537), .B(G113), .ZN(G15) );
  XNOR2_X1 U636 ( .A(G116), .B(KEYINPUT115), .ZN(n540) );
  OR2_X1 U637 ( .A1(n554), .A2(n538), .ZN(n674) );
  INV_X1 U638 ( .A(n674), .ZN(n577) );
  NAND2_X1 U639 ( .A1(n601), .A2(n577), .ZN(n539) );
  XOR2_X1 U640 ( .A(n540), .B(n539), .Z(G18) );
  NAND2_X1 U641 ( .A1(n542), .A2(n710), .ZN(n543) );
  NAND2_X1 U642 ( .A1(n558), .A2(n711), .ZN(n546) );
  XNOR2_X1 U643 ( .A(KEYINPUT86), .B(KEYINPUT39), .ZN(n545) );
  XNOR2_X1 U644 ( .A(n546), .B(n545), .ZN(n578) );
  NAND2_X1 U645 ( .A1(n578), .A2(n547), .ZN(n548) );
  NAND2_X1 U646 ( .A1(n551), .A2(n550), .ZN(n553) );
  INV_X1 U647 ( .A(KEYINPUT46), .ZN(n552) );
  XNOR2_X1 U648 ( .A(n553), .B(n552), .ZN(n574) );
  NAND2_X1 U649 ( .A1(n555), .A2(n554), .ZN(n587) );
  NOR2_X1 U650 ( .A1(n587), .A2(n556), .ZN(n557) );
  NAND2_X1 U651 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U652 ( .A(n559), .B(KEYINPUT108), .ZN(n753) );
  XNOR2_X1 U653 ( .A(n562), .B(KEYINPUT36), .ZN(n563) );
  NAND2_X1 U654 ( .A1(n674), .A2(n679), .ZN(n715) );
  XNOR2_X1 U655 ( .A(n715), .B(KEYINPUT82), .ZN(n603) );
  XNOR2_X1 U656 ( .A(n603), .B(KEYINPUT72), .ZN(n564) );
  NAND2_X1 U657 ( .A1(n564), .A2(n569), .ZN(n567) );
  OR2_X1 U658 ( .A1(n566), .A2(n565), .ZN(n680) );
  NAND2_X1 U659 ( .A1(n715), .A2(KEYINPUT72), .ZN(n568) );
  NOR2_X1 U660 ( .A1(n680), .A2(n568), .ZN(n570) );
  INV_X1 U661 ( .A(KEYINPUT47), .ZN(n569) );
  NOR2_X1 U662 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U663 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U664 ( .A1(n574), .A2(n573), .ZN(n576) );
  INV_X1 U665 ( .A(KEYINPUT48), .ZN(n575) );
  XNOR2_X1 U666 ( .A(n576), .B(n575), .ZN(n582) );
  AND2_X1 U667 ( .A1(n578), .A2(n577), .ZN(n685) );
  INV_X1 U668 ( .A(n579), .ZN(n580) );
  NOR2_X1 U669 ( .A1(n685), .A2(n580), .ZN(n581) );
  NAND2_X1 U670 ( .A1(n582), .A2(n581), .ZN(n627) );
  XNOR2_X1 U671 ( .A(n627), .B(KEYINPUT84), .ZN(n692) );
  NOR2_X1 U672 ( .A1(n692), .A2(n620), .ZN(n619) );
  INV_X1 U673 ( .A(n587), .ZN(n588) );
  NAND2_X1 U674 ( .A1(n589), .A2(n588), .ZN(n591) );
  XNOR2_X1 U675 ( .A(KEYINPUT77), .B(KEYINPUT35), .ZN(n590) );
  XNOR2_X2 U676 ( .A(n591), .B(n590), .ZN(n653) );
  INV_X1 U677 ( .A(KEYINPUT44), .ZN(n612) );
  NAND2_X1 U678 ( .A1(n653), .A2(n612), .ZN(n592) );
  INV_X1 U679 ( .A(KEYINPUT65), .ZN(n613) );
  NAND2_X1 U680 ( .A1(n592), .A2(n613), .ZN(n598) );
  AND2_X1 U681 ( .A1(n694), .A2(n697), .ZN(n593) );
  XNOR2_X1 U682 ( .A(KEYINPUT78), .B(KEYINPUT32), .ZN(n595) );
  INV_X1 U683 ( .A(n609), .ZN(n597) );
  NAND2_X1 U684 ( .A1(n598), .A2(n597), .ZN(n608) );
  INV_X1 U685 ( .A(n671), .ZN(n600) );
  OR2_X1 U686 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U687 ( .A(n602), .B(KEYINPUT100), .ZN(n604) );
  NAND2_X1 U688 ( .A1(n604), .A2(n603), .ZN(n606) );
  AND2_X1 U689 ( .A1(n606), .A2(n605), .ZN(n607) );
  AND2_X2 U690 ( .A1(n608), .A2(n607), .ZN(n617) );
  NAND2_X1 U691 ( .A1(n609), .A2(n613), .ZN(n611) );
  AND2_X1 U692 ( .A1(n653), .A2(KEYINPUT44), .ZN(n610) );
  NAND2_X1 U693 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X2 U696 ( .A(n618), .B(KEYINPUT45), .ZN(n689) );
  NAND2_X1 U697 ( .A1(n619), .A2(n689), .ZN(n624) );
  INV_X1 U698 ( .A(n620), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n621), .A2(KEYINPUT2), .ZN(n622) );
  XOR2_X1 U700 ( .A(KEYINPUT67), .B(n622), .Z(n623) );
  XNOR2_X2 U701 ( .A(n626), .B(n625), .ZN(n630) );
  INV_X1 U702 ( .A(n689), .ZN(n629) );
  XOR2_X1 U703 ( .A(KEYINPUT62), .B(n631), .Z(n632) );
  XNOR2_X1 U704 ( .A(n633), .B(n632), .ZN(n634) );
  NOR2_X1 U705 ( .A1(n634), .A2(n666), .ZN(n636) );
  XOR2_X1 U706 ( .A(KEYINPUT90), .B(KEYINPUT63), .Z(n635) );
  XNOR2_X1 U707 ( .A(n636), .B(n635), .ZN(G57) );
  XOR2_X1 U708 ( .A(KEYINPUT59), .B(n637), .Z(n638) );
  XNOR2_X1 U709 ( .A(n639), .B(n638), .ZN(n640) );
  NOR2_X1 U710 ( .A1(n640), .A2(n666), .ZN(n641) );
  XNOR2_X1 U711 ( .A(n641), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U712 ( .A(KEYINPUT55), .B(KEYINPUT88), .Z(n645) );
  XNOR2_X1 U713 ( .A(KEYINPUT81), .B(KEYINPUT120), .ZN(n643) );
  XNOR2_X1 U714 ( .A(n643), .B(KEYINPUT54), .ZN(n644) );
  XNOR2_X1 U715 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U716 ( .A(n642), .B(n646), .ZN(n647) );
  XNOR2_X1 U717 ( .A(n648), .B(n647), .ZN(n649) );
  NOR2_X1 U718 ( .A1(n649), .A2(n666), .ZN(n650) );
  XNOR2_X1 U719 ( .A(n650), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U720 ( .A(n651), .B(G119), .ZN(G21) );
  XOR2_X1 U721 ( .A(G122), .B(KEYINPUT127), .Z(n652) );
  XNOR2_X1 U722 ( .A(n653), .B(n652), .ZN(G24) );
  NAND2_X1 U723 ( .A1(n661), .A2(G217), .ZN(n654) );
  XOR2_X1 U724 ( .A(n655), .B(n654), .Z(n656) );
  NOR2_X1 U725 ( .A1(n656), .A2(n666), .ZN(G66) );
  NAND2_X1 U726 ( .A1(n661), .A2(G478), .ZN(n659) );
  XNOR2_X1 U727 ( .A(n657), .B(KEYINPUT121), .ZN(n658) );
  XNOR2_X1 U728 ( .A(n659), .B(n658), .ZN(n660) );
  NOR2_X1 U729 ( .A1(n660), .A2(n666), .ZN(G63) );
  NAND2_X1 U730 ( .A1(n661), .A2(G469), .ZN(n665) );
  XOR2_X1 U731 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n663) );
  XNOR2_X1 U732 ( .A(n662), .B(n663), .ZN(n664) );
  XNOR2_X1 U733 ( .A(n665), .B(n664), .ZN(n667) );
  NOR2_X1 U734 ( .A1(n667), .A2(n666), .ZN(G54) );
  NOR2_X1 U735 ( .A1(n679), .A2(n671), .ZN(n668) );
  XOR2_X1 U736 ( .A(G104), .B(n668), .Z(G6) );
  XOR2_X1 U737 ( .A(KEYINPUT26), .B(KEYINPUT112), .Z(n670) );
  XNOR2_X1 U738 ( .A(G107), .B(KEYINPUT27), .ZN(n669) );
  XNOR2_X1 U739 ( .A(n670), .B(n669), .ZN(n673) );
  NOR2_X1 U740 ( .A1(n674), .A2(n671), .ZN(n672) );
  XOR2_X1 U741 ( .A(n673), .B(n672), .Z(G9) );
  NOR2_X1 U742 ( .A1(n680), .A2(n674), .ZN(n678) );
  XOR2_X1 U743 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n676) );
  XNOR2_X1 U744 ( .A(G128), .B(KEYINPUT114), .ZN(n675) );
  XNOR2_X1 U745 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U746 ( .A(n678), .B(n677), .ZN(G30) );
  NOR2_X1 U747 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U748 ( .A(G146), .B(n681), .Z(G48) );
  XNOR2_X1 U749 ( .A(n682), .B(KEYINPUT116), .ZN(n683) );
  XNOR2_X1 U750 ( .A(n683), .B(KEYINPUT37), .ZN(n684) );
  XNOR2_X1 U751 ( .A(G125), .B(n684), .ZN(G27) );
  XOR2_X1 U752 ( .A(G134), .B(n685), .Z(G36) );
  INV_X1 U753 ( .A(n686), .ZN(n687) );
  NOR2_X1 U754 ( .A1(n687), .A2(n707), .ZN(n688) );
  NOR2_X1 U755 ( .A1(n689), .A2(KEYINPUT2), .ZN(n690) );
  NAND2_X1 U756 ( .A1(n747), .A2(n386), .ZN(n693) );
  NOR2_X1 U757 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U758 ( .A(KEYINPUT50), .B(n696), .Z(n703) );
  XOR2_X1 U759 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n700) );
  NAND2_X1 U760 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U761 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U762 ( .A1(n701), .A2(n542), .ZN(n702) );
  NAND2_X1 U763 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U764 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U765 ( .A(KEYINPUT51), .B(n706), .Z(n709) );
  INV_X1 U766 ( .A(n707), .ZN(n708) );
  NAND2_X1 U767 ( .A1(n709), .A2(n708), .ZN(n721) );
  NOR2_X1 U768 ( .A1(n711), .A2(n710), .ZN(n713) );
  NOR2_X1 U769 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U770 ( .A(KEYINPUT118), .B(n714), .Z(n718) );
  XNOR2_X1 U771 ( .A(n716), .B(KEYINPUT119), .ZN(n717) );
  NAND2_X1 U772 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U773 ( .A1(n686), .A2(n719), .ZN(n720) );
  NAND2_X1 U774 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U775 ( .A(KEYINPUT52), .B(n722), .Z(n723) );
  NOR2_X1 U776 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U777 ( .A(KEYINPUT53), .B(n726), .Z(G75) );
  NAND2_X1 U778 ( .A1(n689), .A2(n485), .ZN(n727) );
  XNOR2_X1 U779 ( .A(n727), .B(KEYINPUT122), .ZN(n731) );
  NAND2_X1 U780 ( .A1(G953), .A2(G224), .ZN(n728) );
  XNOR2_X1 U781 ( .A(KEYINPUT61), .B(n728), .ZN(n729) );
  NAND2_X1 U782 ( .A1(n729), .A2(G898), .ZN(n730) );
  NAND2_X1 U783 ( .A1(n731), .A2(n730), .ZN(n738) );
  XOR2_X1 U784 ( .A(n732), .B(G101), .Z(n734) );
  XNOR2_X1 U785 ( .A(n734), .B(n733), .ZN(n736) );
  NAND2_X1 U786 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U787 ( .A(n738), .B(n737), .Z(G69) );
  XOR2_X1 U788 ( .A(KEYINPUT123), .B(n739), .Z(n742) );
  XNOR2_X1 U789 ( .A(n740), .B(KEYINPUT4), .ZN(n741) );
  XNOR2_X1 U790 ( .A(n742), .B(n741), .ZN(n748) );
  XNOR2_X1 U791 ( .A(n748), .B(G227), .ZN(n743) );
  XNOR2_X1 U792 ( .A(n743), .B(KEYINPUT124), .ZN(n744) );
  NAND2_X1 U793 ( .A1(n744), .A2(G900), .ZN(n745) );
  NAND2_X1 U794 ( .A1(G953), .A2(n745), .ZN(n746) );
  XNOR2_X1 U795 ( .A(n746), .B(KEYINPUT125), .ZN(n751) );
  XOR2_X1 U796 ( .A(n748), .B(n747), .Z(n749) );
  NOR2_X1 U797 ( .A1(n749), .A2(G953), .ZN(n750) );
  NOR2_X1 U798 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U799 ( .A(KEYINPUT126), .B(n752), .Z(G72) );
  XNOR2_X1 U800 ( .A(G143), .B(n753), .ZN(G45) );
endmodule

