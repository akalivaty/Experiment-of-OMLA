

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783;

  OR2_X1 U379 ( .A1(n690), .A2(n382), .ZN(n376) );
  NAND2_X1 U380 ( .A1(n634), .A2(n699), .ZN(n621) );
  NOR2_X1 U381 ( .A1(n618), .A2(n730), .ZN(n414) );
  BUF_X1 U382 ( .A(n601), .Z(n617) );
  NAND2_X2 U383 ( .A1(n553), .A2(n552), .ZN(n704) );
  XNOR2_X1 U384 ( .A(n519), .B(n518), .ZN(n530) );
  XNOR2_X1 U385 ( .A(n367), .B(n450), .ZN(n492) );
  XNOR2_X2 U386 ( .A(G119), .B(KEYINPUT3), .ZN(n448) );
  AND2_X2 U387 ( .A1(n712), .A2(n532), .ZN(n541) );
  NAND2_X1 U388 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U389 ( .A1(n387), .A2(n386), .ZN(n689) );
  BUF_X1 U390 ( .A(n530), .Z(n580) );
  XNOR2_X1 U391 ( .A(n469), .B(n468), .ZN(n601) );
  XNOR2_X1 U392 ( .A(n492), .B(n455), .ZN(n756) );
  XNOR2_X1 U393 ( .A(G140), .B(G137), .ZN(n508) );
  NOR2_X2 U394 ( .A1(n601), .A2(n622), .ZN(n405) );
  NOR2_X2 U395 ( .A1(n385), .A2(n358), .ZN(n394) );
  XNOR2_X2 U396 ( .A(n368), .B(KEYINPUT39), .ZN(n634) );
  AND2_X1 U397 ( .A1(n524), .A2(n522), .ZN(n523) );
  XNOR2_X2 U398 ( .A(KEYINPUT68), .B(G101), .ZN(n483) );
  XNOR2_X2 U399 ( .A(n533), .B(KEYINPUT33), .ZN(n746) );
  INV_X1 U400 ( .A(G237), .ZN(n465) );
  NAND2_X1 U401 ( .A1(n645), .A2(n503), .ZN(n391) );
  XNOR2_X1 U402 ( .A(n372), .B(n371), .ZN(n590) );
  INV_X1 U403 ( .A(KEYINPUT74), .ZN(n371) );
  NOR2_X1 U404 ( .A1(n573), .A2(n572), .ZN(n372) );
  NAND2_X1 U405 ( .A1(n357), .A2(n409), .ZN(n408) );
  NAND2_X1 U406 ( .A1(n636), .A2(KEYINPUT65), .ZN(n409) );
  AND2_X1 U407 ( .A1(n654), .A2(n382), .ZN(n379) );
  XNOR2_X1 U408 ( .A(G137), .B(G116), .ZN(n489) );
  XOR2_X1 U409 ( .A(KEYINPUT96), .B(KEYINPUT75), .Z(n487) );
  NOR2_X1 U410 ( .A1(G953), .A2(G237), .ZN(n485) );
  XNOR2_X1 U411 ( .A(G131), .B(G134), .ZN(n481) );
  NOR2_X1 U412 ( .A1(n738), .A2(n392), .ZN(n739) );
  NOR2_X1 U413 ( .A1(n735), .A2(n447), .ZN(n365) );
  INV_X1 U414 ( .A(KEYINPUT105), .ZN(n364) );
  XNOR2_X1 U415 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U416 ( .A(n403), .B(n478), .ZN(n547) );
  XNOR2_X1 U417 ( .A(n448), .B(KEYINPUT85), .ZN(n367) );
  INV_X1 U418 ( .A(KEYINPUT72), .ZN(n449) );
  XNOR2_X1 U419 ( .A(G116), .B(G107), .ZN(n453) );
  XNOR2_X1 U420 ( .A(n497), .B(n496), .ZN(n498) );
  INV_X1 U421 ( .A(G110), .ZN(n496) );
  NAND2_X1 U422 ( .A1(n407), .A2(n751), .ZN(n644) );
  XNOR2_X1 U423 ( .A(n583), .B(KEYINPUT109), .ZN(n625) );
  AND2_X1 U424 ( .A1(n722), .A2(n596), .ZN(n581) );
  BUF_X1 U425 ( .A(n772), .Z(n370) );
  NAND2_X1 U426 ( .A1(n401), .A2(n400), .ZN(n402) );
  NAND2_X1 U427 ( .A1(G234), .A2(G237), .ZN(n471) );
  AND2_X1 U428 ( .A1(n381), .A2(n383), .ZN(n380) );
  NOR2_X1 U429 ( .A1(n606), .A2(n698), .ZN(n383) );
  INV_X1 U430 ( .A(G902), .ZN(n503) );
  XNOR2_X1 U431 ( .A(G119), .B(KEYINPUT24), .ZN(n509) );
  XNOR2_X1 U432 ( .A(G128), .B(G110), .ZN(n510) );
  XNOR2_X1 U433 ( .A(KEYINPUT90), .B(KEYINPUT23), .ZN(n507) );
  NAND2_X1 U434 ( .A1(n396), .A2(n362), .ZN(n395) );
  XNOR2_X1 U435 ( .A(n501), .B(n494), .ZN(n645) );
  XNOR2_X1 U436 ( .A(G122), .B(KEYINPUT103), .ZN(n416) );
  XNOR2_X1 U437 ( .A(KEYINPUT9), .B(KEYINPUT101), .ZN(n417) );
  XOR2_X1 U438 ( .A(KEYINPUT7), .B(KEYINPUT102), .Z(n418) );
  XNOR2_X1 U439 ( .A(G113), .B(G143), .ZN(n437) );
  XOR2_X1 U440 ( .A(KEYINPUT99), .B(G140), .Z(n432) );
  INV_X1 U441 ( .A(KEYINPUT4), .ZN(n461) );
  XNOR2_X1 U442 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n458) );
  XNOR2_X1 U443 ( .A(n410), .B(KEYINPUT83), .ZN(n711) );
  INV_X2 U444 ( .A(G953), .ZN(n772) );
  XNOR2_X1 U445 ( .A(n480), .B(n479), .ZN(n524) );
  NAND2_X1 U446 ( .A1(n547), .A2(n366), .ZN(n480) );
  XNOR2_X1 U447 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U448 ( .A(n444), .B(n443), .ZN(n554) );
  XNOR2_X1 U449 ( .A(n442), .B(n441), .ZN(n443) );
  INV_X1 U450 ( .A(G475), .ZN(n441) );
  INV_X1 U451 ( .A(KEYINPUT94), .ZN(n406) );
  BUF_X1 U452 ( .A(n524), .Z(n560) );
  XNOR2_X1 U453 ( .A(n501), .B(n502), .ZN(n658) );
  XNOR2_X1 U454 ( .A(G104), .B(G107), .ZN(n499) );
  XNOR2_X1 U455 ( .A(n768), .B(n498), .ZN(n500) );
  XNOR2_X1 U456 ( .A(n626), .B(KEYINPUT42), .ZN(n654) );
  AND2_X1 U457 ( .A1(n389), .A2(n388), .ZN(n387) );
  XNOR2_X1 U458 ( .A(n681), .B(n680), .ZN(n682) );
  XOR2_X1 U459 ( .A(n638), .B(KEYINPUT67), .Z(n357) );
  AND2_X1 U460 ( .A1(n361), .A2(n408), .ZN(n358) );
  OR2_X1 U461 ( .A1(n537), .A2(n540), .ZN(n359) );
  NAND2_X1 U462 ( .A1(n568), .A2(n567), .ZN(n360) );
  INV_X1 U463 ( .A(n358), .ZN(n396) );
  OR2_X1 U464 ( .A1(n357), .A2(n411), .ZN(n361) );
  INV_X1 U465 ( .A(KEYINPUT65), .ZN(n411) );
  NAND2_X1 U466 ( .A1(n357), .A2(KEYINPUT65), .ZN(n362) );
  AND2_X1 U467 ( .A1(n637), .A2(n411), .ZN(n363) );
  INV_X1 U468 ( .A(KEYINPUT46), .ZN(n382) );
  NAND2_X1 U469 ( .A1(n393), .A2(n395), .ZN(n397) );
  NAND2_X1 U470 ( .A1(n505), .A2(G221), .ZN(n506) );
  XNOR2_X1 U471 ( .A(n421), .B(n422), .ZN(n505) );
  XNOR2_X1 U472 ( .A(n523), .B(KEYINPUT32), .ZN(n687) );
  XNOR2_X1 U473 ( .A(n756), .B(n464), .ZN(n674) );
  NAND2_X1 U474 ( .A1(n619), .A2(n414), .ZN(n368) );
  NAND2_X1 U475 ( .A1(n712), .A2(n582), .ZN(n548) );
  XNOR2_X2 U476 ( .A(n504), .B(G469), .ZN(n582) );
  NAND2_X1 U477 ( .A1(n369), .A2(n582), .ZN(n583) );
  XNOR2_X1 U478 ( .A(n581), .B(KEYINPUT28), .ZN(n369) );
  NAND2_X1 U479 ( .A1(n642), .A2(n711), .ZN(n751) );
  NAND2_X1 U480 ( .A1(n375), .A2(KEYINPUT46), .ZN(n374) );
  NAND2_X1 U481 ( .A1(n399), .A2(n363), .ZN(n398) );
  NOR2_X1 U482 ( .A1(n663), .A2(G902), .ZN(n428) );
  XNOR2_X1 U483 ( .A(n426), .B(n425), .ZN(n663) );
  XNOR2_X2 U484 ( .A(n771), .B(n484), .ZN(n501) );
  XNOR2_X2 U485 ( .A(n482), .B(n481), .ZN(n771) );
  XNOR2_X2 U486 ( .A(n462), .B(n461), .ZN(n482) );
  NOR2_X2 U487 ( .A1(n377), .A2(n373), .ZN(n627) );
  NAND2_X1 U488 ( .A1(n376), .A2(n374), .ZN(n373) );
  INV_X1 U489 ( .A(n654), .ZN(n375) );
  NAND2_X1 U490 ( .A1(n380), .A2(n378), .ZN(n377) );
  NAND2_X1 U491 ( .A1(n379), .A2(n690), .ZN(n378) );
  AND2_X1 U492 ( .A1(n595), .A2(n594), .ZN(n381) );
  XNOR2_X2 U493 ( .A(n621), .B(n620), .ZN(n690) );
  NAND2_X1 U494 ( .A1(n384), .A2(n641), .ZN(n709) );
  INV_X1 U495 ( .A(n385), .ZN(n384) );
  XNOR2_X1 U496 ( .A(n385), .B(n774), .ZN(n773) );
  NAND2_X2 U497 ( .A1(n640), .A2(n707), .ZN(n385) );
  NAND2_X1 U498 ( .A1(n642), .A2(n370), .ZN(n759) );
  OR2_X1 U499 ( .A1(n538), .A2(n359), .ZN(n386) );
  NAND2_X1 U500 ( .A1(n537), .A2(n540), .ZN(n388) );
  NAND2_X1 U501 ( .A1(n538), .A2(n540), .ZN(n389) );
  AND2_X1 U502 ( .A1(n390), .A2(n562), .ZN(n563) );
  NAND2_X1 U503 ( .A1(n689), .A2(KEYINPUT44), .ZN(n390) );
  XNOR2_X2 U504 ( .A(n525), .B(n495), .ZN(n599) );
  XNOR2_X2 U505 ( .A(n391), .B(G472), .ZN(n525) );
  INV_X1 U506 ( .A(n746), .ZN(n392) );
  NAND2_X1 U507 ( .A1(n394), .A2(n641), .ZN(n393) );
  NAND2_X1 U508 ( .A1(n398), .A2(n397), .ZN(n407) );
  INV_X1 U509 ( .A(n709), .ZN(n399) );
  INV_X1 U510 ( .A(n652), .ZN(n400) );
  INV_X1 U511 ( .A(n687), .ZN(n401) );
  NOR2_X1 U512 ( .A1(n402), .A2(KEYINPUT44), .ZN(n568) );
  NAND2_X1 U513 ( .A1(n402), .A2(KEYINPUT44), .ZN(n528) );
  NAND2_X1 U514 ( .A1(n584), .A2(n477), .ZN(n403) );
  XNOR2_X1 U515 ( .A(n405), .B(n404), .ZN(n584) );
  INV_X1 U516 ( .A(KEYINPUT19), .ZN(n404) );
  NAND2_X1 U517 ( .A1(n543), .A2(n609), .ZN(n549) );
  XNOR2_X2 U518 ( .A(n548), .B(n406), .ZN(n609) );
  NAND2_X1 U519 ( .A1(n640), .A2(n413), .ZN(n410) );
  NOR2_X1 U520 ( .A1(n370), .A2(G952), .ZN(n684) );
  AND2_X1 U521 ( .A1(n515), .A2(G221), .ZN(n412) );
  XOR2_X1 U522 ( .A(n639), .B(KEYINPUT80), .Z(n413) );
  INV_X1 U523 ( .A(KEYINPUT84), .ZN(n565) );
  INV_X1 U524 ( .A(KEYINPUT5), .ZN(n488) );
  INV_X1 U525 ( .A(n596), .ZN(n597) );
  XNOR2_X1 U526 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U527 ( .A(n491), .B(n490), .ZN(n493) );
  XNOR2_X1 U528 ( .A(n462), .B(n416), .ZN(n420) );
  BUF_X1 U529 ( .A(n547), .Z(n543) );
  BUF_X1 U530 ( .A(n668), .Z(n669) );
  INV_X2 U531 ( .A(G143), .ZN(n415) );
  XNOR2_X2 U532 ( .A(n415), .B(G128), .ZN(n462) );
  XNOR2_X1 U533 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U534 ( .A(n420), .B(n419), .Z(n426) );
  NAND2_X1 U535 ( .A1(n772), .A2(G234), .ZN(n422) );
  XNOR2_X1 U536 ( .A(KEYINPUT71), .B(KEYINPUT8), .ZN(n421) );
  NAND2_X1 U537 ( .A1(n505), .A2(G217), .ZN(n424) );
  XOR2_X1 U538 ( .A(G134), .B(n453), .Z(n423) );
  XNOR2_X1 U539 ( .A(n424), .B(n423), .ZN(n425) );
  INV_X1 U540 ( .A(G478), .ZN(n427) );
  XNOR2_X1 U541 ( .A(n428), .B(n427), .ZN(n430) );
  INV_X1 U542 ( .A(KEYINPUT104), .ZN(n429) );
  XNOR2_X1 U543 ( .A(n430), .B(n429), .ZN(n555) );
  NAND2_X1 U544 ( .A1(G214), .A2(n485), .ZN(n431) );
  XNOR2_X1 U545 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U546 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n434) );
  XNOR2_X1 U547 ( .A(G131), .B(KEYINPUT100), .ZN(n433) );
  XNOR2_X1 U548 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U549 ( .A(n436), .B(n435), .ZN(n440) );
  XNOR2_X2 U550 ( .A(G146), .B(G125), .ZN(n456) );
  XNOR2_X1 U551 ( .A(n456), .B(KEYINPUT10), .ZN(n769) );
  XNOR2_X2 U552 ( .A(G122), .B(G104), .ZN(n452) );
  XNOR2_X1 U553 ( .A(n452), .B(n437), .ZN(n438) );
  XNOR2_X1 U554 ( .A(n769), .B(n438), .ZN(n439) );
  XNOR2_X1 U555 ( .A(n440), .B(n439), .ZN(n681) );
  NOR2_X1 U556 ( .A1(G902), .A2(n681), .ZN(n444) );
  INV_X1 U557 ( .A(KEYINPUT13), .ZN(n442) );
  INV_X1 U558 ( .A(n554), .ZN(n552) );
  NAND2_X1 U559 ( .A1(n555), .A2(n552), .ZN(n735) );
  XOR2_X1 U560 ( .A(KEYINPUT92), .B(KEYINPUT21), .Z(n446) );
  XNOR2_X1 U561 ( .A(G902), .B(KEYINPUT15), .ZN(n636) );
  NAND2_X1 U562 ( .A1(n636), .A2(G234), .ZN(n445) );
  XNOR2_X1 U563 ( .A(n445), .B(KEYINPUT20), .ZN(n515) );
  XNOR2_X1 U564 ( .A(n446), .B(n412), .ZN(n715) );
  XNOR2_X1 U565 ( .A(n715), .B(KEYINPUT93), .ZN(n529) );
  INV_X1 U566 ( .A(n529), .ZN(n447) );
  XNOR2_X1 U567 ( .A(n449), .B(G113), .ZN(n450) );
  XNOR2_X1 U568 ( .A(G110), .B(KEYINPUT16), .ZN(n451) );
  XNOR2_X1 U569 ( .A(n452), .B(n451), .ZN(n454) );
  XNOR2_X1 U570 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U571 ( .A(n456), .B(n483), .ZN(n460) );
  NAND2_X1 U572 ( .A1(n772), .A2(G224), .ZN(n457) );
  XNOR2_X1 U573 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U574 ( .A(n460), .B(n459), .ZN(n463) );
  XNOR2_X1 U575 ( .A(n482), .B(n463), .ZN(n464) );
  INV_X1 U576 ( .A(n636), .ZN(n637) );
  OR2_X2 U577 ( .A1(n674), .A2(n637), .ZN(n469) );
  NAND2_X1 U578 ( .A1(n503), .A2(n465), .ZN(n470) );
  NAND2_X1 U579 ( .A1(n470), .A2(G210), .ZN(n467) );
  INV_X1 U580 ( .A(KEYINPUT79), .ZN(n466) );
  AND2_X1 U581 ( .A1(n470), .A2(G214), .ZN(n622) );
  XNOR2_X1 U582 ( .A(n471), .B(KEYINPUT86), .ZN(n472) );
  XNOR2_X1 U583 ( .A(KEYINPUT14), .B(n472), .ZN(n474) );
  NAND2_X1 U584 ( .A1(n474), .A2(G902), .ZN(n473) );
  XOR2_X1 U585 ( .A(KEYINPUT88), .B(n473), .Z(n574) );
  NOR2_X1 U586 ( .A1(G898), .A2(n370), .ZN(n757) );
  NAND2_X1 U587 ( .A1(n574), .A2(n757), .ZN(n476) );
  NAND2_X1 U588 ( .A1(n474), .A2(G952), .ZN(n475) );
  XNOR2_X1 U589 ( .A(n475), .B(KEYINPUT87), .ZN(n743) );
  NAND2_X1 U590 ( .A1(n743), .A2(n370), .ZN(n578) );
  NAND2_X1 U591 ( .A1(n476), .A2(n578), .ZN(n477) );
  INV_X1 U592 ( .A(KEYINPUT0), .ZN(n478) );
  INV_X1 U593 ( .A(KEYINPUT22), .ZN(n479) );
  XNOR2_X1 U594 ( .A(n483), .B(G146), .ZN(n484) );
  NAND2_X1 U595 ( .A1(n485), .A2(G210), .ZN(n486) );
  XNOR2_X1 U596 ( .A(n487), .B(n486), .ZN(n491) );
  XNOR2_X1 U597 ( .A(n492), .B(n493), .ZN(n494) );
  INV_X1 U598 ( .A(KEYINPUT6), .ZN(n495) );
  XNOR2_X1 U599 ( .A(n599), .B(KEYINPUT78), .ZN(n521) );
  XNOR2_X1 U600 ( .A(n508), .B(KEYINPUT89), .ZN(n768) );
  NAND2_X1 U601 ( .A1(G227), .A2(n772), .ZN(n497) );
  XNOR2_X1 U602 ( .A(n500), .B(n499), .ZN(n502) );
  NAND2_X1 U603 ( .A1(n658), .A2(n503), .ZN(n504) );
  XNOR2_X1 U604 ( .A(n582), .B(KEYINPUT1), .ZN(n532) );
  BUF_X1 U605 ( .A(n532), .Z(n713) );
  XNOR2_X1 U606 ( .A(n769), .B(n506), .ZN(n514) );
  XNOR2_X1 U607 ( .A(n508), .B(n507), .ZN(n512) );
  XNOR2_X1 U608 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U609 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U610 ( .A(n514), .B(n513), .ZN(n668) );
  OR2_X2 U611 ( .A1(n668), .A2(G902), .ZN(n519) );
  NAND2_X1 U612 ( .A1(n515), .A2(G217), .ZN(n517) );
  XNOR2_X1 U613 ( .A(KEYINPUT91), .B(KEYINPUT25), .ZN(n516) );
  XNOR2_X1 U614 ( .A(n517), .B(n516), .ZN(n518) );
  INV_X1 U615 ( .A(n580), .ZN(n716) );
  NAND2_X1 U616 ( .A1(n713), .A2(n716), .ZN(n520) );
  NOR2_X1 U617 ( .A1(n521), .A2(n520), .ZN(n522) );
  BUF_X2 U618 ( .A(n525), .Z(n722) );
  OR2_X1 U619 ( .A1(n722), .A2(n580), .ZN(n526) );
  NOR2_X1 U620 ( .A1(n713), .A2(n526), .ZN(n527) );
  AND2_X1 U621 ( .A1(n560), .A2(n527), .ZN(n652) );
  XNOR2_X1 U622 ( .A(n528), .B(KEYINPUT66), .ZN(n564) );
  XNOR2_X2 U623 ( .A(n531), .B(KEYINPUT69), .ZN(n712) );
  NAND2_X1 U624 ( .A1(n541), .A2(n599), .ZN(n533) );
  NAND2_X1 U625 ( .A1(n746), .A2(n543), .ZN(n534) );
  XNOR2_X1 U626 ( .A(n534), .B(KEYINPUT34), .ZN(n538) );
  INV_X1 U627 ( .A(n555), .ZN(n553) );
  NAND2_X1 U628 ( .A1(n553), .A2(n554), .ZN(n536) );
  INV_X1 U629 ( .A(KEYINPUT106), .ZN(n535) );
  XNOR2_X1 U630 ( .A(n536), .B(n535), .ZN(n612) );
  INV_X1 U631 ( .A(n612), .ZN(n537) );
  INV_X1 U632 ( .A(KEYINPUT77), .ZN(n539) );
  XNOR2_X1 U633 ( .A(n539), .B(KEYINPUT35), .ZN(n540) );
  NAND2_X1 U634 ( .A1(n541), .A2(n722), .ZN(n542) );
  XNOR2_X1 U635 ( .A(n542), .B(KEYINPUT97), .ZN(n724) );
  NAND2_X1 U636 ( .A1(n724), .A2(n543), .ZN(n546) );
  INV_X1 U637 ( .A(KEYINPUT98), .ZN(n544) );
  XNOR2_X1 U638 ( .A(n544), .B(KEYINPUT31), .ZN(n545) );
  XNOR2_X1 U639 ( .A(n546), .B(n545), .ZN(n705) );
  XNOR2_X1 U640 ( .A(n549), .B(KEYINPUT95), .ZN(n551) );
  INV_X1 U641 ( .A(n722), .ZN(n550) );
  NAND2_X1 U642 ( .A1(n551), .A2(n550), .ZN(n691) );
  NAND2_X1 U643 ( .A1(n705), .A2(n691), .ZN(n557) );
  NAND2_X1 U644 ( .A1(n555), .A2(n554), .ZN(n702) );
  NAND2_X1 U645 ( .A1(n704), .A2(n702), .ZN(n729) );
  XNOR2_X1 U646 ( .A(n729), .B(KEYINPUT81), .ZN(n573) );
  INV_X1 U647 ( .A(n573), .ZN(n556) );
  NAND2_X1 U648 ( .A1(n557), .A2(n556), .ZN(n561) );
  OR2_X1 U649 ( .A1(n713), .A2(n716), .ZN(n558) );
  NOR2_X1 U650 ( .A1(n558), .A2(n599), .ZN(n559) );
  NAND2_X1 U651 ( .A1(n560), .A2(n559), .ZN(n651) );
  AND2_X1 U652 ( .A1(n561), .A2(n651), .ZN(n562) );
  NAND2_X1 U653 ( .A1(n564), .A2(n563), .ZN(n566) );
  XNOR2_X1 U654 ( .A(n566), .B(n565), .ZN(n569) );
  INV_X1 U655 ( .A(n689), .ZN(n567) );
  NAND2_X1 U656 ( .A1(n569), .A2(n360), .ZN(n571) );
  XNOR2_X1 U657 ( .A(KEYINPUT82), .B(KEYINPUT45), .ZN(n570) );
  XNOR2_X2 U658 ( .A(n571), .B(n570), .ZN(n641) );
  XNOR2_X1 U659 ( .A(KEYINPUT70), .B(KEYINPUT47), .ZN(n572) );
  OR2_X1 U660 ( .A1(n590), .A2(KEYINPUT73), .ZN(n585) );
  INV_X1 U661 ( .A(G900), .ZN(n576) );
  AND2_X1 U662 ( .A1(G953), .A2(n574), .ZN(n575) );
  NAND2_X1 U663 ( .A1(n576), .A2(n575), .ZN(n577) );
  AND2_X1 U664 ( .A1(n578), .A2(n577), .ZN(n607) );
  OR2_X1 U665 ( .A1(n607), .A2(n715), .ZN(n579) );
  NOR2_X1 U666 ( .A1(n580), .A2(n579), .ZN(n596) );
  AND2_X1 U667 ( .A1(n584), .A2(n625), .ZN(n700) );
  NAND2_X1 U668 ( .A1(n585), .A2(n700), .ZN(n589) );
  INV_X1 U669 ( .A(n700), .ZN(n587) );
  NOR2_X1 U670 ( .A1(KEYINPUT73), .A2(KEYINPUT47), .ZN(n586) );
  NAND2_X1 U671 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U672 ( .A1(n589), .A2(n588), .ZN(n595) );
  AND2_X1 U673 ( .A1(n590), .A2(KEYINPUT73), .ZN(n593) );
  INV_X1 U674 ( .A(KEYINPUT47), .ZN(n591) );
  NOR2_X1 U675 ( .A1(n729), .A2(n591), .ZN(n592) );
  NOR2_X1 U676 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U677 ( .A1(n702), .A2(n597), .ZN(n598) );
  AND2_X1 U678 ( .A1(n599), .A2(n598), .ZN(n600) );
  INV_X1 U679 ( .A(n622), .ZN(n732) );
  NAND2_X1 U680 ( .A1(n600), .A2(n732), .ZN(n628) );
  NOR2_X2 U681 ( .A1(n628), .A2(n617), .ZN(n602) );
  XNOR2_X1 U682 ( .A(n602), .B(KEYINPUT36), .ZN(n603) );
  NAND2_X1 U683 ( .A1(n603), .A2(n713), .ZN(n605) );
  INV_X1 U684 ( .A(KEYINPUT111), .ZN(n604) );
  XNOR2_X2 U685 ( .A(n605), .B(n604), .ZN(n782) );
  INV_X1 U686 ( .A(n782), .ZN(n606) );
  INV_X1 U687 ( .A(n607), .ZN(n608) );
  NAND2_X1 U688 ( .A1(n609), .A2(n608), .ZN(n611) );
  INV_X1 U689 ( .A(KEYINPUT76), .ZN(n610) );
  XNOR2_X1 U690 ( .A(n611), .B(n610), .ZN(n619) );
  INV_X1 U691 ( .A(n617), .ZN(n630) );
  NAND2_X1 U692 ( .A1(n612), .A2(n630), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n722), .A2(n732), .ZN(n614) );
  XNOR2_X1 U694 ( .A(KEYINPUT108), .B(KEYINPUT30), .ZN(n613) );
  XNOR2_X1 U695 ( .A(n614), .B(n613), .ZN(n618) );
  NOR2_X1 U696 ( .A1(n615), .A2(n618), .ZN(n616) );
  AND2_X1 U697 ( .A1(n619), .A2(n616), .ZN(n698) );
  XNOR2_X1 U698 ( .A(n617), .B(KEYINPUT38), .ZN(n733) );
  INV_X1 U699 ( .A(n733), .ZN(n730) );
  INV_X1 U700 ( .A(n702), .ZN(n699) );
  XNOR2_X1 U701 ( .A(KEYINPUT110), .B(KEYINPUT40), .ZN(n620) );
  NOR2_X1 U702 ( .A1(n735), .A2(n622), .ZN(n623) );
  NAND2_X1 U703 ( .A1(n623), .A2(n733), .ZN(n624) );
  XNOR2_X1 U704 ( .A(n624), .B(KEYINPUT41), .ZN(n745) );
  NAND2_X1 U705 ( .A1(n625), .A2(n745), .ZN(n626) );
  XNOR2_X1 U706 ( .A(n627), .B(KEYINPUT48), .ZN(n633) );
  NOR2_X1 U707 ( .A1(n713), .A2(n628), .ZN(n629) );
  XNOR2_X1 U708 ( .A(n629), .B(KEYINPUT43), .ZN(n631) );
  NOR2_X1 U709 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U710 ( .A(n632), .B(KEYINPUT107), .ZN(n780) );
  AND2_X2 U711 ( .A1(n633), .A2(n780), .ZN(n640) );
  INV_X1 U712 ( .A(n634), .ZN(n635) );
  OR2_X1 U713 ( .A1(n635), .A2(n704), .ZN(n707) );
  NAND2_X1 U714 ( .A1(n637), .A2(KEYINPUT2), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n707), .A2(KEYINPUT2), .ZN(n639) );
  BUF_X1 U716 ( .A(n641), .Z(n642) );
  INV_X1 U717 ( .A(KEYINPUT64), .ZN(n643) );
  XNOR2_X2 U718 ( .A(n644), .B(n643), .ZN(n679) );
  NAND2_X1 U719 ( .A1(n679), .A2(G472), .ZN(n647) );
  XOR2_X1 U720 ( .A(KEYINPUT62), .B(n645), .Z(n646) );
  XNOR2_X1 U721 ( .A(n647), .B(n646), .ZN(n648) );
  NOR2_X2 U722 ( .A1(n648), .A2(n684), .ZN(n650) );
  INV_X1 U723 ( .A(KEYINPUT63), .ZN(n649) );
  XNOR2_X1 U724 ( .A(n650), .B(n649), .ZN(G57) );
  XNOR2_X1 U725 ( .A(n651), .B(G101), .ZN(G3) );
  XOR2_X1 U726 ( .A(G110), .B(n652), .Z(G12) );
  NOR2_X1 U727 ( .A1(n691), .A2(n702), .ZN(n653) );
  XOR2_X1 U728 ( .A(G104), .B(n653), .Z(G6) );
  XNOR2_X1 U729 ( .A(n654), .B(G137), .ZN(G39) );
  BUF_X1 U730 ( .A(n679), .Z(n667) );
  NAND2_X1 U731 ( .A1(n667), .A2(G469), .ZN(n660) );
  XOR2_X1 U732 ( .A(KEYINPUT119), .B(KEYINPUT57), .Z(n656) );
  XNOR2_X1 U733 ( .A(KEYINPUT58), .B(KEYINPUT118), .ZN(n655) );
  XNOR2_X1 U734 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U735 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U736 ( .A(n660), .B(n659), .ZN(n661) );
  NOR2_X1 U737 ( .A1(n661), .A2(n684), .ZN(G54) );
  NAND2_X1 U738 ( .A1(n667), .A2(G478), .ZN(n665) );
  XOR2_X1 U739 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n662) );
  XNOR2_X1 U740 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U741 ( .A(n665), .B(n664), .ZN(n666) );
  NOR2_X1 U742 ( .A1(n666), .A2(n684), .ZN(G63) );
  NAND2_X1 U743 ( .A1(n667), .A2(G217), .ZN(n671) );
  XOR2_X1 U744 ( .A(KEYINPUT123), .B(n669), .Z(n670) );
  XNOR2_X1 U745 ( .A(n671), .B(n670), .ZN(n672) );
  NOR2_X1 U746 ( .A1(n672), .A2(n684), .ZN(G66) );
  NAND2_X1 U747 ( .A1(n679), .A2(G210), .ZN(n676) );
  XOR2_X1 U748 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n673) );
  XNOR2_X1 U749 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U750 ( .A(n676), .B(n675), .ZN(n677) );
  NOR2_X2 U751 ( .A1(n677), .A2(n684), .ZN(n678) );
  XNOR2_X1 U752 ( .A(n678), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U753 ( .A1(n679), .A2(G475), .ZN(n683) );
  XOR2_X1 U754 ( .A(KEYINPUT120), .B(KEYINPUT59), .Z(n680) );
  XNOR2_X1 U755 ( .A(n683), .B(n682), .ZN(n685) );
  NOR2_X2 U756 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U757 ( .A(n686), .B(KEYINPUT60), .ZN(G60) );
  BUF_X1 U758 ( .A(n687), .Z(n688) );
  XOR2_X1 U759 ( .A(G119), .B(n688), .Z(G21) );
  XOR2_X1 U760 ( .A(G122), .B(n689), .Z(G24) );
  XNOR2_X1 U761 ( .A(n690), .B(G131), .ZN(G33) );
  NOR2_X1 U762 ( .A1(n691), .A2(n704), .ZN(n693) );
  XNOR2_X1 U763 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n692) );
  XNOR2_X1 U764 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U765 ( .A(G107), .B(n694), .ZN(G9) );
  XOR2_X1 U766 ( .A(G128), .B(KEYINPUT29), .Z(n697) );
  INV_X1 U767 ( .A(n704), .ZN(n695) );
  NAND2_X1 U768 ( .A1(n700), .A2(n695), .ZN(n696) );
  XNOR2_X1 U769 ( .A(n697), .B(n696), .ZN(G30) );
  XOR2_X1 U770 ( .A(G143), .B(n698), .Z(G45) );
  NAND2_X1 U771 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U772 ( .A(n701), .B(G146), .ZN(G48) );
  NOR2_X1 U773 ( .A1(n705), .A2(n702), .ZN(n703) );
  XOR2_X1 U774 ( .A(G113), .B(n703), .Z(G15) );
  NOR2_X1 U775 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U776 ( .A(G116), .B(n706), .Z(G18) );
  XOR2_X1 U777 ( .A(n707), .B(G134), .Z(n708) );
  XNOR2_X1 U778 ( .A(n708), .B(KEYINPUT113), .ZN(G36) );
  BUF_X1 U779 ( .A(n709), .Z(n710) );
  NOR2_X1 U780 ( .A1(n711), .A2(n710), .ZN(n750) );
  NOR2_X1 U781 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U782 ( .A(KEYINPUT50), .B(n714), .Z(n720) );
  XNOR2_X1 U783 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n718) );
  NAND2_X1 U784 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U785 ( .A(n718), .B(n717), .Z(n719) );
  NAND2_X1 U786 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U787 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U788 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U789 ( .A(n725), .B(KEYINPUT51), .Z(n726) );
  XNOR2_X1 U790 ( .A(KEYINPUT115), .B(n726), .ZN(n727) );
  NAND2_X1 U791 ( .A1(n727), .A2(n745), .ZN(n728) );
  XOR2_X1 U792 ( .A(n728), .B(KEYINPUT116), .Z(n740) );
  NAND2_X1 U793 ( .A1(n729), .A2(n732), .ZN(n731) );
  NOR2_X1 U794 ( .A1(n731), .A2(n730), .ZN(n737) );
  NOR2_X1 U795 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U796 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U797 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U798 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U799 ( .A(n741), .B(KEYINPUT117), .ZN(n742) );
  XNOR2_X1 U800 ( .A(n742), .B(KEYINPUT52), .ZN(n744) );
  NAND2_X1 U801 ( .A1(n744), .A2(n743), .ZN(n748) );
  NAND2_X1 U802 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U803 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U804 ( .A1(n750), .A2(n749), .ZN(n753) );
  NAND2_X1 U805 ( .A1(n751), .A2(KEYINPUT2), .ZN(n752) );
  AND2_X1 U806 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U807 ( .A1(n370), .A2(n754), .ZN(n755) );
  XOR2_X1 U808 ( .A(KEYINPUT53), .B(n755), .Z(G75) );
  XNOR2_X1 U809 ( .A(n756), .B(G101), .ZN(n758) );
  NOR2_X1 U810 ( .A1(n758), .A2(n757), .ZN(n767) );
  XNOR2_X1 U811 ( .A(n759), .B(KEYINPUT126), .ZN(n765) );
  NAND2_X1 U812 ( .A1(G224), .A2(G953), .ZN(n760) );
  XNOR2_X1 U813 ( .A(n760), .B(KEYINPUT124), .ZN(n761) );
  XNOR2_X1 U814 ( .A(KEYINPUT61), .B(n761), .ZN(n762) );
  NAND2_X1 U815 ( .A1(n762), .A2(G898), .ZN(n763) );
  XOR2_X1 U816 ( .A(KEYINPUT125), .B(n763), .Z(n764) );
  NAND2_X1 U817 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U818 ( .A(n767), .B(n766), .ZN(G69) );
  XNOR2_X1 U819 ( .A(n768), .B(n769), .ZN(n770) );
  XNOR2_X1 U820 ( .A(n771), .B(n770), .ZN(n774) );
  NAND2_X1 U821 ( .A1(n773), .A2(n370), .ZN(n779) );
  XNOR2_X1 U822 ( .A(G227), .B(n774), .ZN(n775) );
  NAND2_X1 U823 ( .A1(n775), .A2(G900), .ZN(n776) );
  XOR2_X1 U824 ( .A(KEYINPUT127), .B(n776), .Z(n777) );
  NAND2_X1 U825 ( .A1(G953), .A2(n777), .ZN(n778) );
  NAND2_X1 U826 ( .A1(n779), .A2(n778), .ZN(G72) );
  XNOR2_X1 U827 ( .A(G140), .B(n780), .ZN(G42) );
  XOR2_X1 U828 ( .A(KEYINPUT37), .B(KEYINPUT112), .Z(n781) );
  XNOR2_X1 U829 ( .A(n782), .B(n781), .ZN(n783) );
  XNOR2_X1 U830 ( .A(G125), .B(n783), .ZN(G27) );
endmodule

