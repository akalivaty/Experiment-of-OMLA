//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n772,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n850, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959;
  INV_X1    g000(.A(KEYINPUT88), .ZN(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  INV_X1    g002(.A(G36gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT14), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT14), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n206), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT87), .ZN(new_n208));
  AND3_X1   g007(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n208), .B1(new_n205), .B2(new_n207), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AND2_X1   g010(.A1(G43gat), .A2(G50gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(G43gat), .A2(G50gat), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT15), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT85), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(new_n204), .ZN(new_n216));
  NAND2_X1  g015(.A1(KEYINPUT85), .A2(G36gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(G29gat), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT86), .ZN(new_n219));
  INV_X1    g018(.A(G50gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(KEYINPUT86), .A2(G50gat), .ZN(new_n222));
  AOI21_X1  g021(.A(G43gat), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT15), .ZN(new_n224));
  INV_X1    g023(.A(G43gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(new_n220), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n214), .B(new_n218), .C1(new_n223), .C2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n202), .B1(new_n211), .B2(new_n227), .ZN(new_n228));
  NOR3_X1   g027(.A1(new_n206), .A2(G29gat), .A3(G36gat), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT14), .B1(new_n203), .B2(new_n204), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT87), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT86), .B(G50gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(new_n225), .ZN(new_n235));
  INV_X1    g034(.A(new_n226), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n214), .A2(new_n218), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n233), .A2(KEYINPUT88), .A3(new_n237), .A4(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n228), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n229), .A2(new_n230), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n214), .B1(new_n241), .B2(new_n218), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT17), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G15gat), .B(G22gat), .ZN(new_n247));
  INV_X1    g046(.A(G1gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT16), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n247), .A2(G1gat), .ZN(new_n252));
  OAI21_X1  g051(.A(G8gat), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G8gat), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n250), .B(new_n254), .C1(G1gat), .C2(new_n247), .ZN(new_n255));
  AND2_X1   g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n240), .A2(KEYINPUT17), .A3(new_n243), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n246), .A2(KEYINPUT89), .A3(new_n256), .A4(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(G229gat), .A2(G233gat), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT17), .B1(new_n240), .B2(new_n243), .ZN(new_n260));
  AOI211_X1 g059(.A(new_n245), .B(new_n242), .C1(new_n228), .C2(new_n239), .ZN(new_n261));
  INV_X1    g060(.A(new_n256), .ZN(new_n262));
  NOR3_X1   g061(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n256), .B1(new_n240), .B2(new_n243), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT89), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n258), .B(new_n259), .C1(new_n263), .C2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT18), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OR2_X1    g068(.A1(new_n264), .A2(new_n265), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n246), .A2(new_n256), .A3(new_n257), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n272), .A2(KEYINPUT18), .A3(new_n259), .A4(new_n258), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n259), .B(KEYINPUT13), .Z(new_n274));
  AND3_X1   g073(.A1(new_n240), .A2(new_n256), .A3(new_n243), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n274), .B1(new_n275), .B2(new_n264), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT90), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n269), .A2(new_n273), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G113gat), .B(G141gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(G197gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT11), .ZN(new_n281));
  INV_X1    g080(.A(G169gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT12), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n278), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n269), .A2(new_n277), .A3(new_n273), .A4(new_n284), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(KEYINPUT91), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT91), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n278), .A2(new_n289), .A3(new_n285), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G8gat), .B(G36gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n292), .B(KEYINPUT74), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(G64gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(G92gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n297));
  INV_X1    g096(.A(G176gat), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT23), .B1(new_n282), .B2(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  AND2_X1   g101(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n304));
  OAI211_X1 g103(.A(KEYINPUT23), .B(new_n282), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  OR2_X1    g105(.A1(G183gat), .A2(G190gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(G183gat), .A2(G190gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(KEYINPUT24), .A3(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(KEYINPUT24), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n297), .B1(new_n306), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT25), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n314), .B1(new_n300), .B2(KEYINPUT23), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n302), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT66), .B1(new_n316), .B2(new_n312), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT24), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n318), .B1(G183gat), .B2(G190gat), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n310), .B1(new_n319), .B2(new_n307), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT66), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n320), .A2(new_n321), .A3(new_n302), .A4(new_n315), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n313), .A2(new_n317), .A3(new_n322), .ZN(new_n323));
  OR2_X1    g122(.A1(new_n301), .A2(KEYINPUT26), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n301), .A2(KEYINPUT26), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n324), .B(new_n325), .C1(new_n282), .C2(new_n298), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT27), .B(G183gat), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT28), .B1(new_n328), .B2(G190gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT28), .ZN(new_n330));
  INV_X1    g129(.A(G190gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n327), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n326), .A2(new_n329), .A3(new_n332), .A4(new_n308), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n323), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G226gat), .A2(G233gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n335), .B(KEYINPUT72), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT29), .ZN(new_n339));
  AND3_X1   g138(.A1(new_n323), .A2(KEYINPUT73), .A3(new_n333), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT73), .B1(new_n323), .B2(new_n333), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n336), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n338), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G197gat), .B(G204gat), .ZN(new_n345));
  INV_X1    g144(.A(G211gat), .ZN(new_n346));
  INV_X1    g145(.A(G218gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n345), .B1(KEYINPUT22), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G211gat), .B(G218gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT71), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n344), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n351), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n340), .A2(new_n341), .A3(new_n343), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n336), .A2(KEYINPUT29), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n334), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n356), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n296), .B1(new_n355), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT73), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n334), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n323), .A2(KEYINPUT73), .A3(new_n333), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT29), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n337), .B1(new_n367), .B2(new_n336), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n353), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(new_n361), .A3(new_n295), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n363), .A2(KEYINPUT30), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT30), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n369), .A2(new_n372), .A3(new_n361), .A4(new_n295), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G225gat), .A2(G233gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n376), .A2(KEYINPUT5), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT75), .ZN(new_n378));
  XNOR2_X1  g177(.A(G141gat), .B(G148gat), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT2), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n380), .B1(G155gat), .B2(G162gat), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n378), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G155gat), .B(G162gat), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n378), .B(new_n383), .C1(new_n379), .C2(new_n381), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT76), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G127gat), .B(G134gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  XOR2_X1   g190(.A(G113gat), .B(G120gat), .Z(new_n392));
  INV_X1    g191(.A(KEYINPUT67), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT1), .ZN(new_n395));
  XNOR2_X1  g194(.A(G113gat), .B(G120gat), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n395), .B1(new_n396), .B2(KEYINPUT67), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n391), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n392), .A2(new_n390), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT76), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n385), .A2(new_n402), .A3(KEYINPUT3), .A4(new_n386), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n389), .A2(new_n401), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT4), .ZN(new_n406));
  INV_X1    g205(.A(new_n400), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n393), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n396), .A2(KEYINPUT67), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n395), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n407), .B1(new_n410), .B2(new_n391), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n406), .B1(new_n411), .B2(new_n387), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(new_n406), .A3(new_n387), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n412), .B1(KEYINPUT78), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n411), .A2(new_n387), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n415), .A2(KEYINPUT78), .A3(KEYINPUT4), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n377), .B(new_n405), .C1(new_n414), .C2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT5), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n385), .A2(new_n386), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n401), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n415), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n419), .B1(new_n422), .B2(new_n376), .ZN(new_n423));
  NOR3_X1   g222(.A1(new_n401), .A2(new_n420), .A3(KEYINPUT4), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n375), .B1(new_n424), .B2(new_n412), .ZN(new_n425));
  INV_X1    g224(.A(new_n405), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n428));
  XNOR2_X1  g227(.A(G1gat), .B(G29gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(G57gat), .B(G85gat), .ZN(new_n431));
  XOR2_X1   g230(.A(new_n430), .B(new_n431), .Z(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n418), .A2(new_n427), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n433), .B1(new_n418), .B2(new_n427), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n436), .B(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n374), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(G228gat), .A2(G233gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n404), .A2(new_n339), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT81), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n404), .A2(KEYINPUT81), .A3(new_n339), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n353), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n388), .B1(new_n351), .B2(KEYINPUT29), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n420), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n440), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n440), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n441), .A2(new_n351), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT80), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n441), .A2(KEYINPUT80), .A3(new_n351), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n449), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  XOR2_X1   g253(.A(G78gat), .B(G106gat), .Z(new_n455));
  NOR3_X1   g254(.A1(new_n448), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  XOR2_X1   g256(.A(KEYINPUT79), .B(KEYINPUT31), .Z(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(G22gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(G50gat), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n455), .B1(new_n448), .B2(new_n454), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n457), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n460), .ZN(new_n463));
  INV_X1    g262(.A(new_n461), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n463), .B1(new_n464), .B2(new_n456), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n439), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n323), .A2(new_n411), .A3(new_n333), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT69), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n334), .A2(new_n401), .ZN(new_n471));
  NAND2_X1  g270(.A1(G227gat), .A2(G233gat), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT69), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n323), .A2(new_n411), .A3(new_n333), .A4(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n470), .A2(new_n471), .A3(new_n472), .A4(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(KEYINPUT34), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT32), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n470), .A2(new_n471), .A3(new_n474), .ZN(new_n478));
  INV_X1    g277(.A(new_n472), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT33), .B1(new_n478), .B2(new_n479), .ZN(new_n481));
  XNOR2_X1  g280(.A(G15gat), .B(G43gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n482), .B(G71gat), .ZN(new_n483));
  INV_X1    g282(.A(G99gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n480), .A2(new_n481), .A3(new_n486), .ZN(new_n487));
  AOI221_X4 g286(.A(new_n477), .B1(KEYINPUT33), .B2(new_n485), .C1(new_n478), .C2(new_n479), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n476), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n481), .A2(new_n486), .ZN(new_n490));
  INV_X1    g289(.A(new_n480), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n476), .ZN(new_n493));
  INV_X1    g292(.A(new_n488), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n489), .A2(new_n495), .A3(KEYINPUT70), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT36), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT70), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n492), .A2(new_n493), .A3(new_n498), .A4(new_n494), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n489), .A2(new_n495), .A3(KEYINPUT36), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n368), .A2(new_n353), .ZN(new_n503));
  NOR3_X1   g302(.A1(new_n357), .A2(new_n356), .A3(new_n360), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT37), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT38), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT37), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n361), .B(new_n507), .C1(new_n344), .C2(new_n354), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n505), .A2(new_n506), .A3(new_n296), .A4(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n436), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n437), .A2(KEYINPUT83), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT83), .ZN(new_n512));
  AOI211_X1 g311(.A(new_n512), .B(new_n433), .C1(new_n418), .C2(new_n427), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n510), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n437), .A2(KEYINPUT6), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n509), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n508), .A2(new_n296), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n507), .B1(new_n369), .B2(new_n361), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT38), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n370), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n466), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n405), .B1(new_n414), .B2(new_n417), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT39), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n523), .A3(new_n376), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n524), .A2(new_n433), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT84), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n415), .A2(new_n421), .A3(new_n375), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n415), .A2(KEYINPUT4), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT78), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n528), .B1(new_n424), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n426), .B1(new_n530), .B2(new_n416), .ZN(new_n531));
  OAI211_X1 g330(.A(KEYINPUT39), .B(new_n527), .C1(new_n531), .C2(new_n375), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n525), .A2(new_n526), .A3(KEYINPUT40), .A4(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n532), .A2(KEYINPUT40), .A3(new_n433), .A4(new_n524), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT84), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n418), .A2(new_n427), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(new_n432), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n512), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n437), .A2(KEYINPUT83), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n533), .A2(new_n535), .A3(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT82), .B(KEYINPUT40), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n542), .B1(new_n525), .B2(new_n532), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n541), .A2(new_n374), .A3(new_n543), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n468), .B(new_n502), .C1(new_n521), .C2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n466), .A2(new_n495), .A3(new_n489), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT35), .B1(new_n546), .B2(new_n439), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n496), .A2(new_n499), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n514), .A2(new_n515), .B1(new_n371), .B2(new_n373), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT35), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n548), .A2(new_n549), .A3(new_n550), .A4(new_n466), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n291), .B1(new_n545), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(G71gat), .ZN(new_n554));
  INV_X1    g353(.A(G78gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(G71gat), .A2(G78gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT92), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n556), .A2(KEYINPUT92), .A3(new_n557), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(G57gat), .B(G64gat), .Z(new_n563));
  INV_X1    g362(.A(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n557), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(G64gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(G57gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(KEYINPUT93), .B(G57gat), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n569), .B1(new_n570), .B2(new_n568), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n557), .B1(new_n556), .B2(new_n564), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n567), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT94), .B(KEYINPUT21), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n562), .A2(new_n566), .B1(new_n571), .B2(new_n572), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT21), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n578), .A3(new_n256), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n579), .B1(new_n576), .B2(new_n256), .ZN(new_n580));
  XNOR2_X1  g379(.A(G127gat), .B(G155gat), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n580), .A2(new_n581), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g385(.A(G231gat), .B(G233gat), .C1(new_n582), .C2(new_n583), .ZN(new_n587));
  XNOR2_X1  g386(.A(G183gat), .B(G211gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT20), .ZN(new_n589));
  XNOR2_X1  g388(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n586), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n591), .B1(new_n586), .B2(new_n587), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G134gat), .B(G162gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT99), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT98), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT97), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT7), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT7), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT97), .ZN(new_n601));
  AND2_X1   g400(.A1(G85gat), .A2(G92gat), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  OR2_X1    g402(.A1(G85gat), .A2(G92gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(G85gat), .A2(G92gat), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n605), .A2(KEYINPUT97), .A3(new_n600), .ZN(new_n606));
  NAND2_X1  g405(.A1(G99gat), .A2(G106gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT8), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n603), .A2(new_n604), .A3(new_n606), .A4(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n607), .ZN(new_n610));
  NOR2_X1   g409(.A1(G99gat), .A2(G106gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n598), .A2(KEYINPUT7), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n615), .A2(new_n605), .B1(KEYINPUT8), .B2(new_n607), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n616), .A2(new_n612), .A3(new_n604), .A4(new_n603), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n246), .A2(new_n597), .A3(new_n619), .A4(new_n257), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n597), .A2(KEYINPUT17), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n244), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT41), .ZN(new_n624));
  NAND2_X1  g423(.A1(G232gat), .A2(G233gat), .ZN(new_n625));
  OAI22_X1  g424(.A1(new_n623), .A2(new_n619), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n596), .B1(new_n621), .B2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n625), .A2(new_n624), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n244), .A2(new_n622), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n628), .B1(new_n629), .B2(new_n618), .ZN(new_n630));
  INV_X1    g429(.A(new_n596), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(new_n631), .A3(new_n620), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n625), .A2(new_n624), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT96), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(new_n331), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G218gat), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n627), .A2(new_n632), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n636), .B1(new_n627), .B2(new_n632), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n594), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(G230gat), .ZN(new_n643));
  INV_X1    g442(.A(G233gat), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n616), .A2(new_n647), .A3(new_n604), .A4(new_n603), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT101), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n613), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n647), .B1(new_n612), .B2(KEYINPUT101), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n609), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n577), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n573), .ZN(new_n657));
  AOI22_X1  g456(.A1(new_n560), .A2(new_n561), .B1(new_n563), .B2(new_n565), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n614), .B(new_n617), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n654), .B1(new_n653), .B2(new_n659), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n656), .A2(new_n660), .A3(KEYINPUT10), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT10), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n619), .A2(new_n574), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n646), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(G120gat), .B(G148gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(new_n298), .ZN(new_n666));
  INV_X1    g465(.A(G204gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n656), .A2(new_n660), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n664), .B(new_n669), .C1(new_n646), .C2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n653), .A2(new_n659), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT102), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n673), .A2(new_n662), .A3(new_n655), .ZN(new_n674));
  INV_X1    g473(.A(new_n663), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n645), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n670), .A2(new_n646), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n668), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n671), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n642), .A2(KEYINPUT103), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(new_n641), .B2(new_n679), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n553), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n438), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G1gat), .ZN(G1324gat));
  INV_X1    g487(.A(new_n374), .ZN(new_n689));
  OR2_X1    g488(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n690));
  NAND2_X1  g489(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n691));
  AND4_X1   g490(.A1(new_n689), .A2(new_n685), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n254), .B1(new_n685), .B2(new_n689), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT42), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(KEYINPUT42), .B2(new_n692), .ZN(G1325gat));
  AOI21_X1  g494(.A(G15gat), .B1(new_n685), .B2(new_n548), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n500), .A2(G15gat), .A3(new_n501), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT104), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n696), .B1(new_n685), .B2(new_n698), .ZN(G1326gat));
  NAND2_X1  g498(.A1(new_n685), .A2(new_n467), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT43), .B(G22gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1327gat));
  NAND2_X1  g501(.A1(new_n545), .A2(new_n552), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(new_n638), .B2(new_n639), .ZN(new_n705));
  INV_X1    g504(.A(new_n639), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n706), .A2(KEYINPUT108), .A3(new_n637), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n703), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n640), .B1(new_n545), .B2(new_n552), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n291), .A2(new_n594), .A3(new_n679), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(KEYINPUT106), .Z(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(G29gat), .B1(new_n717), .B2(new_n438), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n712), .A2(new_n715), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n719), .A2(new_n203), .A3(new_n686), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT105), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n721), .A2(KEYINPUT45), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(KEYINPUT45), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n718), .B1(new_n722), .B2(new_n723), .ZN(G1328gat));
  OR3_X1    g523(.A1(new_n717), .A2(KEYINPUT109), .A3(new_n374), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n216), .A2(new_n217), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(KEYINPUT109), .B1(new_n717), .B2(new_n374), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n725), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n715), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n730), .A2(new_n727), .A3(new_n374), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT46), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n729), .A2(new_n732), .ZN(G1329gat));
  NAND3_X1  g532(.A1(new_n719), .A2(new_n225), .A3(new_n548), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT110), .ZN(new_n735));
  OAI21_X1  g534(.A(G43gat), .B1(new_n717), .B2(new_n502), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT111), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT47), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n735), .B(new_n736), .C1(new_n738), .C2(KEYINPUT47), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(G1330gat));
  INV_X1    g541(.A(KEYINPUT113), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n719), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n730), .A2(KEYINPUT112), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n745), .A2(new_n467), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n234), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n466), .A2(new_n234), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n714), .A2(new_n716), .A3(new_n749), .ZN(new_n750));
  AOI211_X1 g549(.A(new_n743), .B(KEYINPUT48), .C1(new_n748), .C2(new_n750), .ZN(new_n751));
  OR2_X1    g550(.A1(new_n743), .A2(KEYINPUT48), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n743), .A2(KEYINPUT48), .ZN(new_n753));
  AND4_X1   g552(.A1(new_n752), .A2(new_n748), .A3(new_n753), .A4(new_n750), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n751), .A2(new_n754), .ZN(G1331gat));
  INV_X1    g554(.A(new_n291), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n756), .B1(new_n545), .B2(new_n552), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n641), .A2(new_n680), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n686), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(new_n570), .ZN(G1332gat));
  NOR2_X1   g561(.A1(new_n759), .A2(new_n374), .ZN(new_n763));
  NOR2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  AND2_X1   g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n763), .B2(new_n764), .ZN(G1333gat));
  OAI21_X1  g566(.A(G71gat), .B1(new_n759), .B2(new_n502), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n548), .A2(new_n554), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n759), .B2(new_n769), .ZN(new_n770));
  XOR2_X1   g569(.A(new_n770), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g570(.A1(new_n759), .A2(new_n466), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(new_n555), .ZN(G1335gat));
  NOR2_X1   g572(.A1(new_n756), .A2(new_n594), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n712), .A2(new_n713), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n705), .A2(new_n707), .ZN(new_n776));
  AOI211_X1 g575(.A(new_n776), .B(new_n709), .C1(new_n545), .C2(new_n552), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n679), .B(new_n774), .C1(new_n775), .C2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(G85gat), .B1(new_n778), .B2(new_n438), .ZN(new_n779));
  INV_X1    g578(.A(new_n640), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n703), .A2(new_n780), .A3(new_n774), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT114), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n712), .A2(KEYINPUT51), .A3(new_n774), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n781), .A2(KEYINPUT114), .A3(new_n782), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n438), .A2(new_n680), .A3(G85gat), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n779), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g589(.A(new_n790), .B(KEYINPUT115), .Z(G1336gat));
  OAI21_X1  g590(.A(G92gat), .B1(new_n778), .B2(new_n374), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n374), .A2(G92gat), .A3(new_n680), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n786), .A2(new_n787), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n792), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n783), .A2(KEYINPUT116), .A3(new_n785), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n781), .A2(new_n798), .A3(new_n782), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n797), .A2(new_n793), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n792), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT117), .B1(new_n801), .B2(KEYINPUT52), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n803));
  AOI211_X1 g602(.A(new_n803), .B(new_n795), .C1(new_n792), .C2(new_n800), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n796), .B1(new_n802), .B2(new_n804), .ZN(G1337gat));
  OAI21_X1  g604(.A(G99gat), .B1(new_n778), .B2(new_n502), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n786), .A2(new_n484), .A3(new_n548), .A4(new_n787), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n806), .B1(new_n807), .B2(new_n680), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(KEYINPUT118), .ZN(G1338gat));
  OAI21_X1  g608(.A(G106gat), .B1(new_n778), .B2(new_n466), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n466), .A2(G106gat), .A3(new_n680), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n786), .A2(new_n787), .A3(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n810), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n797), .A2(new_n799), .A3(new_n811), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n814), .B1(new_n816), .B2(new_n813), .ZN(G1339gat));
  INV_X1    g616(.A(new_n594), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n674), .A2(new_n645), .A3(new_n675), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n664), .A2(KEYINPUT54), .A3(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n669), .B1(new_n676), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n820), .A2(new_n822), .A3(KEYINPUT55), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n823), .A2(new_n671), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825));
  INV_X1    g624(.A(new_n820), .ZN(new_n826));
  INV_X1    g625(.A(new_n822), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n288), .A2(new_n824), .A3(new_n290), .A4(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n259), .B1(new_n272), .B2(new_n258), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n275), .A2(new_n264), .A3(new_n274), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n283), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n679), .A2(new_n287), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n708), .B1(new_n829), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n824), .A2(new_n828), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n287), .A2(new_n832), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n835), .A2(new_n776), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n818), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n642), .A2(new_n680), .A3(new_n291), .ZN(new_n839));
  AOI211_X1 g638(.A(new_n438), .B(new_n689), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n840), .A2(new_n466), .A3(new_n548), .ZN(new_n841));
  OAI21_X1  g640(.A(G113gat), .B1(new_n841), .B2(new_n291), .ZN(new_n842));
  INV_X1    g641(.A(new_n546), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n291), .A2(G113gat), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(G1340gat));
  OAI21_X1  g645(.A(G120gat), .B1(new_n841), .B2(new_n680), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n680), .A2(G120gat), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n847), .B1(new_n844), .B2(new_n848), .ZN(G1341gat));
  INV_X1    g648(.A(new_n844), .ZN(new_n850));
  AOI21_X1  g649(.A(G127gat), .B1(new_n850), .B2(new_n594), .ZN(new_n851));
  INV_X1    g650(.A(G127gat), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n841), .A2(new_n852), .A3(new_n818), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n851), .A2(new_n853), .ZN(G1342gat));
  NOR3_X1   g653(.A1(new_n844), .A2(G134gat), .A3(new_n640), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT56), .ZN(new_n856));
  OAI21_X1  g655(.A(G134gat), .B1(new_n841), .B2(new_n640), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1343gat));
  NAND2_X1  g657(.A1(new_n838), .A2(new_n839), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n467), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n502), .A2(new_n686), .A3(new_n374), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n291), .A2(G141gat), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT122), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n861), .B(KEYINPUT119), .ZN(new_n866));
  XOR2_X1   g665(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n867));
  OAI21_X1  g666(.A(new_n867), .B1(new_n826), .B2(new_n827), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n288), .A2(new_n824), .A3(new_n290), .A4(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n780), .B1(new_n869), .B2(new_n833), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n818), .B1(new_n870), .B2(new_n837), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT121), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n873), .B(new_n818), .C1(new_n870), .C2(new_n837), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n839), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(KEYINPUT57), .A3(new_n467), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n860), .A2(new_n877), .ZN(new_n878));
  AOI211_X1 g677(.A(new_n291), .B(new_n866), .C1(new_n876), .C2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(G141gat), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n865), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT58), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT58), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n883), .B(new_n865), .C1(new_n879), .C2(new_n880), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(G1344gat));
  INV_X1    g684(.A(G148gat), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n862), .A2(new_n886), .A3(new_n679), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n866), .B1(new_n876), .B2(new_n878), .ZN(new_n888));
  AOI211_X1 g687(.A(KEYINPUT59), .B(new_n886), .C1(new_n888), .C2(new_n679), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT59), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n466), .A2(KEYINPUT57), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n835), .A2(new_n640), .A3(new_n836), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n818), .B1(new_n870), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n681), .A2(new_n683), .A3(new_n291), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n896), .B1(new_n860), .B2(KEYINPUT57), .ZN(new_n897));
  INV_X1    g696(.A(new_n866), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n897), .A2(new_n679), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n890), .B1(new_n899), .B2(G148gat), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n887), .B1(new_n889), .B2(new_n900), .ZN(G1345gat));
  AOI21_X1  g700(.A(G155gat), .B1(new_n862), .B2(new_n594), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n594), .A2(G155gat), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT123), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n902), .B1(new_n888), .B2(new_n904), .ZN(G1346gat));
  AOI21_X1  g704(.A(G162gat), .B1(new_n862), .B2(new_n780), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n708), .A2(G162gat), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n888), .B2(new_n907), .ZN(G1347gat));
  NOR2_X1   g707(.A1(new_n686), .A2(new_n374), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n548), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(KEYINPUT124), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n859), .A2(new_n466), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n282), .B1(new_n912), .B2(new_n756), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n546), .B1(new_n838), .B2(new_n839), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n909), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n915), .A2(G169gat), .A3(new_n291), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  XOR2_X1   g716(.A(new_n917), .B(KEYINPUT125), .Z(G1348gat));
  INV_X1    g717(.A(new_n915), .ZN(new_n919));
  AOI21_X1  g718(.A(G176gat), .B1(new_n919), .B2(new_n679), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n680), .A2(new_n304), .A3(new_n303), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n912), .B2(new_n921), .ZN(G1349gat));
  NAND2_X1  g721(.A1(new_n912), .A2(new_n594), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(G183gat), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n919), .A2(new_n594), .A3(new_n327), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g726(.A(new_n331), .B1(new_n912), .B2(new_n780), .ZN(new_n928));
  XOR2_X1   g727(.A(new_n928), .B(KEYINPUT61), .Z(new_n929));
  NAND3_X1  g728(.A1(new_n919), .A2(new_n331), .A3(new_n708), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1351gat));
  NAND2_X1  g730(.A1(new_n894), .A2(new_n895), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n891), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n502), .A2(new_n909), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n466), .B1(new_n838), .B2(new_n839), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n933), .B(new_n935), .C1(new_n877), .C2(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(G197gat), .B1(new_n937), .B2(new_n291), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n860), .A2(new_n934), .ZN(new_n939));
  INV_X1    g738(.A(G197gat), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n939), .A2(new_n940), .A3(new_n756), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n938), .A2(new_n941), .ZN(G1352gat));
  NAND3_X1  g741(.A1(new_n939), .A2(new_n667), .A3(new_n679), .ZN(new_n943));
  XOR2_X1   g742(.A(new_n943), .B(KEYINPUT62), .Z(new_n944));
  AND3_X1   g743(.A1(new_n897), .A2(new_n679), .A3(new_n935), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n667), .B2(new_n945), .ZN(G1353gat));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n947), .B1(new_n937), .B2(new_n818), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n897), .A2(KEYINPUT126), .A3(new_n594), .A4(new_n935), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n948), .A2(new_n949), .A3(G211gat), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT63), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n948), .A2(new_n949), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n939), .A2(new_n346), .A3(new_n594), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1354gat));
  NOR3_X1   g755(.A1(new_n937), .A2(new_n347), .A3(new_n640), .ZN(new_n957));
  AOI21_X1  g756(.A(G218gat), .B1(new_n939), .B2(new_n708), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


