//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 1 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n848, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953;
  INV_X1    g000(.A(KEYINPUT64), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT23), .ZN(new_n203));
  NOR3_X1   g002(.A1(new_n203), .A2(G169gat), .A3(G176gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n202), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT23), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n209), .A2(KEYINPUT64), .A3(new_n205), .ZN(new_n210));
  INV_X1    g009(.A(G169gat), .ZN(new_n211));
  INV_X1    g010(.A(G176gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(new_n203), .ZN(new_n214));
  NAND4_X1  g013(.A1(new_n207), .A2(new_n210), .A3(KEYINPUT25), .A4(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216));
  AND2_X1   g015(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n216), .B1(new_n217), .B2(G190gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT24), .ZN(new_n220));
  AND3_X1   g019(.A1(new_n219), .A2(KEYINPUT65), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT65), .B1(new_n219), .B2(new_n220), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n218), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT66), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT66), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n218), .B(new_n225), .C1(new_n221), .C2(new_n222), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n215), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  AND3_X1   g026(.A1(new_n214), .A2(new_n205), .A3(new_n209), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n219), .A2(new_n220), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n218), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT25), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT26), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n205), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT68), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n234), .A3(new_n213), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT68), .B1(new_n236), .B2(new_n208), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n208), .A2(new_n232), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(new_n240), .A3(new_n219), .ZN(new_n241));
  INV_X1    g040(.A(G183gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT27), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT27), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G183gat), .ZN(new_n245));
  INV_X1    g044(.A(G190gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n243), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  AND2_X1   g046(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n248));
  NOR2_X1   g047(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n247), .B(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n241), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n240), .B1(new_n239), .B2(new_n219), .ZN(new_n253));
  OAI22_X1  g052(.A1(new_n227), .A2(new_n231), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT29), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G226gat), .A2(G233gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT75), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n256), .A2(KEYINPUT75), .A3(new_n257), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(new_n257), .B(KEYINPUT73), .Z(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n224), .A2(new_n226), .ZN(new_n265));
  INV_X1    g064(.A(new_n215), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n231), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n239), .A2(new_n219), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT69), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(new_n241), .A3(new_n251), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n264), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G197gat), .B(G204gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT22), .ZN(new_n274));
  INV_X1    g073(.A(G211gat), .ZN(new_n275));
  INV_X1    g074(.A(G218gat), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G211gat), .B(G218gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n279), .A2(new_n273), .A3(new_n277), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n272), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n256), .A2(new_n264), .ZN(new_n286));
  INV_X1    g085(.A(new_n257), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n252), .A2(new_n253), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n287), .B1(new_n288), .B2(new_n267), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT74), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT74), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n254), .A2(new_n291), .A3(new_n287), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n286), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n262), .A2(new_n285), .B1(new_n293), .B2(new_n284), .ZN(new_n294));
  XNOR2_X1  g093(.A(G8gat), .B(G36gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(KEYINPUT76), .ZN(new_n296));
  XNOR2_X1  g095(.A(G64gat), .B(G92gat), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n296), .B(new_n297), .Z(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n294), .A2(KEYINPUT30), .A3(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT78), .B(KEYINPUT30), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n293), .A2(new_n284), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT75), .B1(new_n256), .B2(new_n257), .ZN(new_n303));
  AOI211_X1 g102(.A(new_n259), .B(new_n287), .C1(new_n254), .C2(new_n255), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n285), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n301), .B1(new_n306), .B2(new_n298), .ZN(new_n307));
  NAND2_X1  g106(.A1(G225gat), .A2(G233gat), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT4), .ZN(new_n310));
  OR2_X1    g109(.A1(KEYINPUT81), .A2(G141gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(KEYINPUT81), .A2(G141gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(G148gat), .A3(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G141gat), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT82), .B1(new_n314), .B2(G148gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT82), .ZN(new_n316));
  INV_X1    g115(.A(G148gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(new_n317), .A3(G141gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n313), .A2(new_n315), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT2), .ZN(new_n320));
  INV_X1    g119(.A(G155gat), .ZN(new_n321));
  INV_X1    g120(.A(G162gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n317), .A2(G141gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n314), .A2(G148gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT80), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT2), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n324), .B1(new_n329), .B2(KEYINPUT2), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n328), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT79), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n324), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(KEYINPUT79), .A2(G155gat), .A3(G162gat), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n335), .A2(new_n336), .B1(new_n321), .B2(new_n322), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n319), .A2(new_n325), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT1), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(G113gat), .B2(G120gat), .ZN(new_n340));
  AND2_X1   g139(.A1(G113gat), .A2(G120gat), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT70), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  XOR2_X1   g141(.A(G127gat), .B(G134gat), .Z(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G127gat), .B(G134gat), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n345), .B(KEYINPUT70), .C1(new_n341), .C2(new_n340), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n310), .B1(new_n338), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n309), .B1(new_n348), .B2(KEYINPUT83), .ZN(new_n349));
  INV_X1    g148(.A(new_n312), .ZN(new_n350));
  NOR2_X1   g149(.A1(KEYINPUT81), .A2(G141gat), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n350), .A2(new_n351), .A3(new_n317), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n315), .A2(new_n318), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n325), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n333), .A2(new_n337), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n347), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT4), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT83), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n338), .A2(new_n310), .A3(new_n347), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n315), .A2(new_n318), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n361), .A2(new_n313), .B1(new_n324), .B2(new_n323), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n320), .A2(KEYINPUT80), .B1(G155gat), .B2(G162gat), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n363), .A2(new_n330), .B1(new_n326), .B2(new_n327), .ZN(new_n364));
  INV_X1    g163(.A(new_n336), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT79), .B1(G155gat), .B2(G162gat), .ZN(new_n366));
  OAI22_X1  g165(.A1(new_n365), .A2(new_n366), .B1(G155gat), .B2(G162gat), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT3), .B1(new_n362), .B2(new_n368), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n344), .A2(new_n346), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT3), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n355), .A2(new_n354), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n369), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n349), .A2(new_n360), .A3(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT85), .B(KEYINPUT5), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n355), .A2(new_n354), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n370), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n356), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT84), .B1(new_n378), .B2(new_n309), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n378), .A2(KEYINPUT84), .A3(new_n309), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n374), .B(new_n375), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  XOR2_X1   g180(.A(G1gat), .B(G29gat), .Z(new_n382));
  XNOR2_X1  g181(.A(G57gat), .B(G85gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT86), .B(KEYINPUT0), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n375), .A2(new_n309), .ZN(new_n388));
  AND4_X1   g187(.A1(new_n310), .A2(new_n347), .A3(new_n354), .A4(new_n355), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n373), .B(new_n388), .C1(new_n348), .C2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT87), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n357), .A2(new_n359), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT87), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n392), .A2(new_n393), .A3(new_n373), .A4(new_n388), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n381), .A2(new_n387), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT6), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n387), .B1(new_n381), .B2(new_n395), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI211_X1 g199(.A(new_n397), .B(new_n387), .C1(new_n381), .C2(new_n395), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n300), .B(new_n307), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n347), .B1(new_n288), .B2(new_n267), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n271), .B(new_n370), .C1(new_n231), .C2(new_n227), .ZN(new_n404));
  INV_X1    g203(.A(G227gat), .ZN(new_n405));
  INV_X1    g204(.A(G233gat), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n403), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT32), .ZN(new_n409));
  XOR2_X1   g208(.A(KEYINPUT71), .B(KEYINPUT33), .Z(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G15gat), .B(G43gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(G71gat), .B(G99gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n409), .A2(new_n411), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n410), .B1(new_n414), .B2(KEYINPUT72), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n417), .B1(KEYINPUT72), .B2(new_n414), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n408), .A2(KEYINPUT32), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n407), .B1(new_n403), .B2(new_n404), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT34), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI211_X1 g222(.A(KEYINPUT34), .B(new_n407), .C1(new_n403), .C2(new_n404), .ZN(new_n424));
  OR2_X1    g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n423), .A2(new_n424), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n427), .A2(new_n416), .A3(new_n419), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT88), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n283), .A2(new_n255), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n338), .B1(new_n430), .B2(new_n371), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n283), .B1(new_n372), .B2(new_n255), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n429), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT29), .B1(new_n281), .B2(new_n282), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n376), .B1(new_n434), .B2(KEYINPUT3), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT29), .B1(new_n338), .B2(new_n371), .ZN(new_n436));
  OAI211_X1 g235(.A(KEYINPUT88), .B(new_n435), .C1(new_n436), .C2(new_n283), .ZN(new_n437));
  NAND2_X1  g236(.A1(G228gat), .A2(G233gat), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n433), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n438), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n429), .B(new_n440), .C1(new_n431), .C2(new_n432), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(G22gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n439), .A2(G22gat), .A3(new_n441), .ZN(new_n445));
  XNOR2_X1  g244(.A(G78gat), .B(G106gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(KEYINPUT31), .B(G50gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n446), .B(new_n447), .ZN(new_n448));
  AND4_X1   g247(.A1(KEYINPUT89), .A2(new_n444), .A3(new_n445), .A4(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT89), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n451), .A2(new_n448), .B1(new_n444), .B2(new_n445), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n426), .B(new_n428), .C1(new_n449), .C2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT77), .B1(new_n306), .B2(new_n298), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT77), .ZN(new_n455));
  AOI211_X1 g254(.A(new_n455), .B(new_n299), .C1(new_n302), .C2(new_n305), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n402), .A2(new_n453), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT35), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT91), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT91), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n455), .B1(new_n294), .B2(new_n299), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n306), .A2(KEYINPUT77), .A3(new_n298), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n399), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n465), .A2(new_n397), .A3(new_n396), .ZN(new_n466));
  INV_X1    g265(.A(new_n401), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n464), .A2(new_n468), .A3(new_n300), .A4(new_n307), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n461), .B(KEYINPUT35), .C1(new_n469), .C2(new_n453), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT90), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT35), .B1(new_n466), .B2(new_n467), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n472), .A2(new_n464), .A3(new_n300), .A4(new_n307), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n471), .B1(new_n473), .B2(new_n453), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n300), .A2(new_n307), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n457), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n453), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n476), .A2(KEYINPUT90), .A3(new_n477), .A4(new_n472), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n460), .A2(new_n470), .A3(new_n474), .A4(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n468), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT37), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n294), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n298), .B1(new_n306), .B2(KEYINPUT37), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT38), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n299), .B1(new_n294), .B2(new_n481), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT38), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n481), .B1(new_n293), .B2(new_n283), .ZN(new_n487));
  INV_X1    g286(.A(new_n262), .ZN(new_n488));
  OR2_X1    g287(.A1(new_n272), .A2(new_n283), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n485), .A2(new_n486), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n294), .A2(new_n299), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n480), .A2(new_n484), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n308), .B1(new_n392), .B2(new_n373), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT39), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n386), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT39), .B1(new_n378), .B2(new_n309), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n496), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT40), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n465), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n500), .B1(new_n499), .B2(new_n498), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(new_n457), .B2(new_n475), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n449), .A2(new_n452), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n493), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n469), .A2(new_n503), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n426), .A2(new_n428), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n507), .B(KEYINPUT36), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n505), .A2(new_n506), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n479), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(G190gat), .B(G218gat), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G43gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(G50gat), .ZN(new_n515));
  INV_X1    g314(.A(G50gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(G43gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT14), .ZN(new_n519));
  INV_X1    g318(.A(G29gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n522));
  AOI21_X1  g321(.A(G36gat), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n520), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT92), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT15), .B1(new_n517), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n518), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n527), .ZN(new_n529));
  INV_X1    g328(.A(new_n518), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n529), .B(new_n530), .C1(new_n523), .C2(new_n524), .ZN(new_n531));
  OR3_X1    g330(.A1(new_n523), .A2(KEYINPUT15), .A3(new_n524), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n528), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT93), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n528), .A2(KEYINPUT93), .A3(new_n531), .A4(new_n532), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT17), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(KEYINPUT99), .B(KEYINPUT7), .ZN(new_n539));
  NAND2_X1  g338(.A1(G85gat), .A2(G92gat), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n540), .ZN(new_n542));
  NAND2_X1  g341(.A1(G99gat), .A2(G106gat), .ZN(new_n543));
  INV_X1    g342(.A(G85gat), .ZN(new_n544));
  INV_X1    g343(.A(G92gat), .ZN(new_n545));
  AOI22_X1  g344(.A1(KEYINPUT8), .A2(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n541), .A2(new_n542), .A3(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G99gat), .B(G106gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT100), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n547), .A2(new_n549), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n552), .B1(new_n533), .B2(KEYINPUT17), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n535), .A2(new_n536), .ZN(new_n555));
  AND2_X1   g354(.A1(G232gat), .A2(G233gat), .ZN(new_n556));
  AOI22_X1  g355(.A1(new_n555), .A2(new_n552), .B1(KEYINPUT41), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n513), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n558), .A2(KEYINPUT102), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n554), .A2(new_n513), .A3(new_n557), .ZN(new_n560));
  XOR2_X1   g359(.A(G134gat), .B(G162gat), .Z(new_n561));
  NOR2_X1   g360(.A1(new_n556), .A2(KEYINPUT41), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n558), .A2(KEYINPUT102), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n559), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n563), .B1(new_n560), .B2(new_n558), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT101), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g368(.A(KEYINPUT101), .B(new_n563), .C1(new_n560), .C2(new_n558), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n566), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT9), .ZN(new_n573));
  INV_X1    g372(.A(G71gat), .ZN(new_n574));
  INV_X1    g373(.A(G78gat), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT97), .ZN(new_n577));
  XOR2_X1   g376(.A(G57gat), .B(G64gat), .Z(new_n578));
  INV_X1    g377(.A(KEYINPUT97), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n579), .B(new_n573), .C1(new_n574), .C2(new_n575), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n577), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(G71gat), .B(G78gat), .Z(new_n582));
  AND2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n581), .A2(new_n582), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n585), .A2(KEYINPUT21), .ZN(new_n586));
  AND2_X1   g385(.A1(G231gat), .A2(G233gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(G127gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(G8gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(G15gat), .B(G22gat), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n592), .A2(G1gat), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT94), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n591), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT16), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n592), .B1(new_n596), .B2(G1gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n595), .B(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n599), .B1(KEYINPUT21), .B2(new_n585), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n590), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n588), .B(G127gat), .ZN(new_n602));
  INV_X1    g401(.A(new_n600), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G183gat), .B(G211gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT98), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(new_n321), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n606), .B(new_n608), .ZN(new_n609));
  AND3_X1   g408(.A1(new_n601), .A2(new_n604), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n609), .B1(new_n601), .B2(new_n604), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n572), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(G230gat), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n614), .A2(new_n406), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n547), .A2(new_n549), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n547), .A2(new_n549), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n585), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n581), .B(new_n582), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n550), .A2(new_n619), .A3(new_n551), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT10), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n618), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n552), .A2(KEYINPUT10), .A3(new_n585), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n615), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n618), .A2(new_n620), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n615), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G120gat), .B(G148gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(G176gat), .B(G204gat), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n629), .B(new_n630), .Z(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n628), .A2(new_n632), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n595), .B(new_n598), .Z(new_n637));
  NAND3_X1  g436(.A1(new_n637), .A2(new_n535), .A3(new_n536), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n555), .A2(new_n599), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G229gat), .A2(G233gat), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n641), .B(KEYINPUT95), .Z(new_n642));
  XOR2_X1   g441(.A(new_n642), .B(KEYINPUT13), .Z(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G113gat), .B(G141gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(G197gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT11), .B(G169gat), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n646), .B(new_n647), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT12), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n533), .A2(KEYINPUT17), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n637), .A2(new_n650), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n639), .B(new_n642), .C1(new_n651), .C2(new_n537), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT18), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n644), .B(new_n649), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n652), .A2(new_n653), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT96), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n652), .A2(KEYINPUT96), .A3(new_n653), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n655), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n649), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n644), .B1(new_n652), .B2(new_n653), .ZN(new_n662));
  INV_X1    g461(.A(new_n656), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n613), .A2(new_n636), .A3(new_n666), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n511), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n480), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT103), .B(G1gat), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1324gat));
  INV_X1    g470(.A(new_n668), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT104), .B(KEYINPUT16), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(G8gat), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n672), .A2(new_n476), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n476), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n591), .B1(new_n668), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(KEYINPUT42), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n678), .B1(KEYINPUT42), .B2(new_n675), .ZN(G1325gat));
  OR3_X1    g478(.A1(new_n672), .A2(G15gat), .A3(new_n507), .ZN(new_n680));
  OAI21_X1  g479(.A(G15gat), .B1(new_n672), .B2(new_n509), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(G1326gat));
  NAND2_X1  g481(.A1(new_n668), .A2(new_n503), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT43), .B(G22gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1327gat));
  AOI21_X1  g484(.A(new_n572), .B1(new_n479), .B2(new_n510), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n612), .A2(new_n666), .A3(new_n636), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n689), .A2(new_n520), .A3(new_n480), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT45), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n686), .A2(KEYINPUT44), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693));
  AOI211_X1 g492(.A(new_n693), .B(new_n572), .C1(new_n479), .C2(new_n510), .ZN(new_n694));
  INV_X1    g493(.A(new_n687), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n692), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(G29gat), .B1(new_n697), .B2(new_n468), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n691), .A2(new_n698), .ZN(G1328gat));
  NOR3_X1   g498(.A1(new_n688), .A2(G36gat), .A3(new_n476), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT46), .ZN(new_n701));
  OAI21_X1  g500(.A(G36gat), .B1(new_n697), .B2(new_n476), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(G1329gat));
  XNOR2_X1  g502(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n514), .B1(new_n696), .B2(new_n508), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n688), .A2(G43gat), .A3(new_n507), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n511), .A2(new_n571), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n693), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n686), .A2(KEYINPUT44), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n709), .A2(new_n508), .A3(new_n710), .A4(new_n687), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT106), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n692), .A2(new_n694), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n713), .A2(new_n714), .A3(new_n508), .A4(new_n687), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n712), .A2(new_n715), .A3(G43gat), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT47), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n706), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n707), .B1(new_n716), .B2(new_n718), .ZN(G1330gat));
  NAND2_X1  g518(.A1(new_n689), .A2(KEYINPUT107), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT107), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n504), .B1(new_n688), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(G50gat), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT48), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n504), .A2(new_n516), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n696), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n724), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n727), .ZN(new_n729));
  OAI21_X1  g528(.A(KEYINPUT48), .B1(new_n729), .B2(new_n723), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(G1331gat));
  NAND2_X1  g530(.A1(new_n666), .A2(new_n636), .ZN(new_n732));
  AOI211_X1 g531(.A(new_n613), .B(new_n732), .C1(new_n479), .C2(new_n510), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n480), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g534(.A(new_n476), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT108), .ZN(new_n738));
  NOR2_X1   g537(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(G1333gat));
  NOR2_X1   g539(.A1(new_n509), .A2(new_n574), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n733), .A2(KEYINPUT109), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT109), .B1(new_n733), .B2(new_n741), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n733), .A2(new_n426), .A3(new_n428), .ZN(new_n744));
  OAI22_X1  g543(.A1(new_n742), .A2(new_n743), .B1(G71gat), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g545(.A1(new_n733), .A2(new_n503), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g547(.A1(new_n732), .A2(new_n612), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT110), .Z(new_n750));
  NAND2_X1  g549(.A1(new_n713), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(G85gat), .B1(new_n751), .B2(new_n468), .ZN(new_n752));
  INV_X1    g551(.A(new_n612), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n666), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n686), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n686), .A2(KEYINPUT51), .A3(new_n755), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n760), .A2(new_n544), .A3(new_n480), .A4(new_n636), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n752), .A2(new_n761), .ZN(G1336gat));
  AND4_X1   g561(.A1(KEYINPUT51), .A2(new_n511), .A3(new_n571), .A4(new_n755), .ZN(new_n763));
  XOR2_X1   g562(.A(KEYINPUT111), .B(KEYINPUT51), .Z(new_n764));
  AOI21_X1  g563(.A(new_n764), .B1(new_n686), .B2(new_n755), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n636), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n476), .A2(G92gat), .A3(new_n767), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n709), .A2(new_n676), .A3(new_n710), .A4(new_n750), .ZN(new_n769));
  AOI22_X1  g568(.A1(new_n766), .A2(new_n768), .B1(new_n769), .B2(G92gat), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n760), .A2(new_n768), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n771), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n769), .A2(G92gat), .ZN(new_n774));
  OAI22_X1  g573(.A1(new_n770), .A2(new_n771), .B1(new_n773), .B2(new_n774), .ZN(G1337gat));
  OAI21_X1  g574(.A(G99gat), .B1(new_n751), .B2(new_n509), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n767), .A2(G99gat), .A3(new_n507), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(G1338gat));
  NOR3_X1   g578(.A1(new_n504), .A2(new_n767), .A3(G106gat), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(new_n763), .B2(new_n765), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI211_X1 g582(.A(KEYINPUT112), .B(new_n780), .C1(new_n763), .C2(new_n765), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n709), .A2(new_n503), .A3(new_n710), .A4(new_n750), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G106gat), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n783), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT53), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(KEYINPUT113), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n713), .A2(new_n790), .A3(new_n503), .A4(new_n750), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n789), .A2(new_n791), .A3(G106gat), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT53), .B1(new_n760), .B2(new_n780), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n788), .A2(new_n794), .ZN(G1339gat));
  NAND4_X1  g594(.A1(new_n572), .A2(new_n612), .A3(new_n767), .A4(new_n666), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n658), .A2(new_n659), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n599), .B1(new_n533), .B2(KEYINPUT17), .ZN(new_n799));
  AOI22_X1  g598(.A1(new_n538), .A2(new_n799), .B1(new_n599), .B2(new_n555), .ZN(new_n800));
  OAI22_X1  g599(.A1(new_n800), .A2(new_n642), .B1(new_n640), .B2(new_n643), .ZN(new_n801));
  AOI22_X1  g600(.A1(new_n798), .A2(new_n655), .B1(new_n648), .B2(new_n801), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n622), .A2(new_n623), .A3(new_n615), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n803), .A2(new_n624), .A3(new_n804), .ZN(new_n805));
  XOR2_X1   g604(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  AOI211_X1 g606(.A(new_n615), .B(new_n807), .C1(new_n622), .C2(new_n623), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT115), .B1(new_n808), .B2(new_n631), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n624), .A2(new_n806), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n810), .A2(new_n811), .A3(new_n632), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n805), .B1(new_n809), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n633), .B1(new_n813), .B2(KEYINPUT55), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n809), .A2(new_n812), .ZN(new_n815));
  INV_X1    g614(.A(new_n805), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n571), .A2(new_n802), .A3(new_n814), .A4(new_n819), .ZN(new_n820));
  AOI22_X1  g619(.A1(new_n660), .A2(new_n664), .B1(new_n817), .B2(new_n818), .ZN(new_n821));
  AOI22_X1  g620(.A1(new_n821), .A2(new_n814), .B1(new_n802), .B2(new_n636), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n820), .B1(new_n822), .B2(new_n571), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n797), .B1(new_n823), .B2(new_n753), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n476), .A2(new_n480), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n824), .A2(new_n453), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT116), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n665), .A2(new_n814), .A3(new_n819), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n802), .A2(new_n636), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n571), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n820), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n753), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n796), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n477), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n828), .B1(new_n835), .B2(new_n825), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n827), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(G113gat), .B1(new_n837), .B2(new_n666), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n826), .B(KEYINPUT117), .ZN(new_n839));
  INV_X1    g638(.A(G113gat), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n839), .A2(new_n840), .A3(new_n665), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n838), .A2(new_n841), .ZN(G1340gat));
  OAI21_X1  g641(.A(G120gat), .B1(new_n837), .B2(new_n767), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n767), .A2(G120gat), .ZN(new_n844));
  XOR2_X1   g643(.A(new_n844), .B(KEYINPUT118), .Z(new_n845));
  NAND2_X1  g644(.A1(new_n839), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n843), .A2(new_n846), .ZN(G1341gat));
  NAND3_X1  g646(.A1(new_n826), .A2(new_n589), .A3(new_n612), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n753), .B1(new_n827), .B2(new_n836), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n848), .B1(new_n849), .B2(new_n589), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT119), .ZN(G1342gat));
  OAI21_X1  g650(.A(G134gat), .B1(new_n837), .B2(new_n572), .ZN(new_n852));
  NOR2_X1   g651(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n824), .A2(new_n453), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n476), .A2(new_n571), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n855), .A2(G134gat), .A3(new_n468), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n853), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n857), .B(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n852), .A2(new_n859), .ZN(G1343gat));
  NAND2_X1  g659(.A1(new_n834), .A2(new_n503), .ZN(new_n861));
  XNOR2_X1  g660(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n834), .A2(new_n865), .A3(new_n503), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n825), .A2(new_n508), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n864), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  OAI22_X1  g667(.A1(new_n868), .A2(new_n666), .B1(new_n351), .B2(new_n350), .ZN(new_n869));
  INV_X1    g668(.A(new_n861), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n867), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n314), .A3(new_n665), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT58), .ZN(G1344gat));
  AOI21_X1  g674(.A(KEYINPUT57), .B1(new_n834), .B2(new_n503), .ZN(new_n876));
  AOI211_X1 g675(.A(new_n504), .B(new_n862), .C1(new_n833), .C2(new_n796), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n636), .B(new_n867), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(G148gat), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n864), .A2(new_n636), .A3(new_n866), .A4(new_n867), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n317), .A2(KEYINPUT59), .ZN(new_n881));
  AOI22_X1  g680(.A1(new_n879), .A2(KEYINPUT59), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n871), .A2(G148gat), .A3(new_n767), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT122), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n883), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n880), .A2(new_n881), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n888), .B1(new_n878), .B2(G148gat), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n885), .B(new_n886), .C1(new_n887), .C2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n884), .A2(new_n890), .ZN(G1345gat));
  NAND3_X1  g690(.A1(new_n872), .A2(new_n321), .A3(new_n612), .ZN(new_n892));
  OAI21_X1  g691(.A(G155gat), .B1(new_n868), .B2(new_n753), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT123), .ZN(G1346gat));
  OAI21_X1  g694(.A(G162gat), .B1(new_n868), .B2(new_n572), .ZN(new_n896));
  OR4_X1    g695(.A1(G162gat), .A2(new_n855), .A3(new_n508), .A4(new_n468), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(new_n861), .B2(new_n897), .ZN(G1347gat));
  NOR2_X1   g697(.A1(new_n476), .A2(new_n480), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n854), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n900), .A2(new_n666), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(new_n211), .ZN(G1348gat));
  NOR2_X1   g701(.A1(new_n900), .A2(new_n767), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(new_n212), .ZN(G1349gat));
  NAND3_X1  g703(.A1(new_n854), .A2(new_n612), .A3(new_n899), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n243), .A2(new_n245), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n907), .B1(new_n242), .B2(new_n905), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g708(.A1(new_n854), .A2(new_n571), .A3(new_n899), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n246), .B1(new_n911), .B2(KEYINPUT61), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT61), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n913), .A2(KEYINPUT124), .A3(new_n914), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n910), .A2(G190gat), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n910), .B(new_n912), .C1(new_n911), .C2(KEYINPUT61), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT125), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n915), .A2(KEYINPUT125), .A3(new_n916), .A4(new_n917), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1351gat));
  NAND2_X1  g721(.A1(new_n509), .A2(new_n899), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n861), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(G197gat), .B1(new_n924), .B2(new_n665), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n865), .B1(new_n824), .B2(new_n504), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n834), .A2(new_n503), .A3(new_n863), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n665), .A2(G197gat), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n925), .B1(new_n928), .B2(new_n929), .ZN(G1352gat));
  NOR4_X1   g729(.A1(new_n861), .A2(G204gat), .A3(new_n767), .A4(new_n923), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT62), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n928), .A2(new_n636), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(G204gat), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1353gat));
  INV_X1    g734(.A(KEYINPUT63), .ZN(new_n936));
  INV_X1    g735(.A(new_n923), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n612), .B(new_n937), .C1(new_n876), .C2(new_n877), .ZN(new_n938));
  OAI21_X1  g737(.A(G211gat), .B1(new_n938), .B2(KEYINPUT126), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n940), .B1(new_n928), .B2(new_n612), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n936), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n928), .A2(new_n940), .A3(new_n612), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n938), .A2(KEYINPUT126), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n943), .A2(new_n944), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n924), .A2(new_n275), .A3(new_n612), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1354gat));
  AOI21_X1  g747(.A(G218gat), .B1(new_n924), .B2(new_n571), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT127), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n949), .A2(new_n950), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n572), .A2(new_n276), .ZN(new_n953));
  AOI211_X1 g752(.A(new_n951), .B(new_n952), .C1(new_n928), .C2(new_n953), .ZN(G1355gat));
endmodule


