

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779;

  XNOR2_X1 U374 ( .A(n580), .B(KEYINPUT1), .ZN(n701) );
  NOR2_X1 U375 ( .A1(G237), .A2(G953), .ZN(n508) );
  OR2_X2 U376 ( .A1(n457), .A2(n456), .ZN(n708) );
  XNOR2_X2 U377 ( .A(n371), .B(n370), .ZN(n426) );
  XNOR2_X2 U378 ( .A(n527), .B(n494), .ZN(n554) );
  XNOR2_X2 U379 ( .A(n554), .B(n495), .ZN(n507) );
  AND2_X2 U380 ( .A1(n585), .A2(n569), .ZN(n559) );
  XNOR2_X2 U381 ( .A(n546), .B(n547), .ZN(n585) );
  XNOR2_X1 U382 ( .A(n578), .B(KEYINPUT19), .ZN(n599) );
  INV_X1 U383 ( .A(KEYINPUT64), .ZN(n642) );
  AND2_X1 U384 ( .A1(n749), .A2(n648), .ZN(n750) );
  AND2_X1 U385 ( .A1(n697), .A2(n639), .ZN(n640) );
  AND2_X1 U386 ( .A1(n449), .A2(n447), .ZN(n446) );
  XNOR2_X1 U387 ( .A(n378), .B(n377), .ZN(n685) );
  NOR2_X1 U388 ( .A1(n722), .A2(n571), .ZN(n572) );
  XNOR2_X1 U389 ( .A(n410), .B(KEYINPUT28), .ZN(n568) );
  XNOR2_X1 U390 ( .A(n600), .B(KEYINPUT0), .ZN(n613) );
  INV_X4 U391 ( .A(G953), .ZN(n771) );
  NAND2_X1 U392 ( .A1(n416), .A2(n520), .ZN(n582) );
  XNOR2_X2 U393 ( .A(KEYINPUT20), .B(n488), .ZN(n491) );
  XNOR2_X1 U394 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X1 U395 ( .A1(G237), .A2(G902), .ZN(n514) );
  INV_X1 U396 ( .A(n673), .ZN(n428) );
  NAND2_X1 U397 ( .A1(n643), .A2(n513), .ZN(n458) );
  INV_X1 U398 ( .A(G134), .ZN(n494) );
  XNOR2_X1 U399 ( .A(KEYINPUT4), .B(G131), .ZN(n495) );
  NAND2_X1 U400 ( .A1(n601), .A2(n357), .ZN(n432) );
  NOR2_X1 U401 ( .A1(n387), .A2(n367), .ZN(n431) );
  AND2_X1 U402 ( .A1(n364), .A2(n354), .ZN(n384) );
  NAND2_X1 U403 ( .A1(n603), .A2(n386), .ZN(n385) );
  OR2_X1 U404 ( .A1(n661), .A2(G902), .ZN(n442) );
  NAND2_X2 U405 ( .A1(n398), .A2(n395), .ZN(n705) );
  OR2_X1 U406 ( .A1(n753), .A2(n396), .ZN(n395) );
  AND2_X1 U407 ( .A1(n400), .A2(n399), .ZN(n398) );
  AND2_X1 U408 ( .A1(n575), .A2(n366), .ZN(n407) );
  OR2_X1 U409 ( .A1(n685), .A2(n471), .ZN(n468) );
  NAND2_X1 U410 ( .A1(KEYINPUT80), .A2(KEYINPUT47), .ZN(n471) );
  XNOR2_X1 U411 ( .A(G146), .B(G137), .ZN(n509) );
  AND2_X2 U412 ( .A1(n705), .A2(n706), .ZN(n623) );
  INV_X1 U413 ( .A(KEYINPUT48), .ZN(n463) );
  NAND2_X1 U414 ( .A1(n427), .A2(n630), .ZN(n392) );
  AND2_X1 U415 ( .A1(n429), .A2(n428), .ZN(n427) );
  AND2_X1 U416 ( .A1(n687), .A2(n361), .ZN(n588) );
  NAND2_X1 U417 ( .A1(n458), .A2(n461), .ZN(n457) );
  NAND2_X1 U418 ( .A1(G472), .A2(n460), .ZN(n459) );
  XNOR2_X1 U419 ( .A(n473), .B(n506), .ZN(n522) );
  XNOR2_X1 U420 ( .A(n382), .B(G116), .ZN(n473) );
  XNOR2_X1 U421 ( .A(G113), .B(KEYINPUT3), .ZN(n382) );
  XNOR2_X1 U422 ( .A(G143), .B(G131), .ZN(n537) );
  XNOR2_X1 U423 ( .A(G122), .B(G113), .ZN(n540) );
  XOR2_X1 U424 ( .A(G140), .B(G104), .Z(n541) );
  XNOR2_X1 U425 ( .A(n507), .B(n497), .ZN(n766) );
  XNOR2_X1 U426 ( .A(n424), .B(n423), .ZN(n521) );
  XNOR2_X1 U427 ( .A(G110), .B(G107), .ZN(n423) );
  XNOR2_X1 U428 ( .A(n498), .B(G104), .ZN(n424) );
  INV_X1 U429 ( .A(KEYINPUT72), .ZN(n498) );
  INV_X1 U430 ( .A(G125), .ZN(n485) );
  XOR2_X1 U431 ( .A(KEYINPUT17), .B(KEYINPUT4), .Z(n528) );
  XNOR2_X1 U432 ( .A(n533), .B(KEYINPUT78), .ZN(n534) );
  NOR2_X1 U433 ( .A1(n568), .A2(n580), .ZN(n436) );
  AND2_X1 U434 ( .A1(n435), .A2(n434), .ZN(n433) );
  NAND2_X1 U435 ( .A1(n721), .A2(n367), .ZN(n435) );
  NAND2_X1 U436 ( .A1(n720), .A2(n367), .ZN(n434) );
  NAND2_X1 U437 ( .A1(n446), .A2(n443), .ZN(n394) );
  NAND2_X1 U438 ( .A1(n445), .A2(n444), .ZN(n443) );
  AND2_X1 U439 ( .A1(n717), .A2(n448), .ZN(n444) );
  NAND2_X1 U440 ( .A1(n592), .A2(n718), .ZN(n578) );
  XNOR2_X1 U441 ( .A(n588), .B(KEYINPUT108), .ZN(n376) );
  NOR2_X1 U442 ( .A1(n628), .A2(n732), .ZN(n441) );
  BUF_X1 U443 ( .A(n613), .Z(n628) );
  INV_X1 U444 ( .A(n622), .ZN(n430) );
  XNOR2_X1 U445 ( .A(n389), .B(n368), .ZN(n374) );
  INV_X1 U446 ( .A(KEYINPUT22), .ZN(n602) );
  XNOR2_X1 U447 ( .A(n523), .B(n522), .ZN(n411) );
  XNOR2_X1 U448 ( .A(n521), .B(n421), .ZN(n523) );
  XNOR2_X1 U449 ( .A(n422), .B(G122), .ZN(n421) );
  XNOR2_X1 U450 ( .A(KEYINPUT69), .B(KEYINPUT16), .ZN(n422) );
  XNOR2_X1 U451 ( .A(n467), .B(n465), .ZN(n753) );
  XNOR2_X1 U452 ( .A(n466), .B(n483), .ZN(n465) );
  XNOR2_X1 U453 ( .A(n450), .B(n360), .ZN(n467) );
  INV_X1 U454 ( .A(KEYINPUT70), .ZN(n452) );
  NAND2_X1 U455 ( .A1(n470), .A2(KEYINPUT47), .ZN(n469) );
  INV_X1 U456 ( .A(KEYINPUT46), .ZN(n464) );
  INV_X1 U457 ( .A(n691), .ZN(n380) );
  XNOR2_X1 U458 ( .A(n489), .B(n402), .ZN(n401) );
  XNOR2_X1 U459 ( .A(n490), .B(n359), .ZN(n402) );
  NOR2_X1 U460 ( .A1(n387), .A2(KEYINPUT30), .ZN(n386) );
  NAND2_X1 U461 ( .A1(n513), .A2(G902), .ZN(n461) );
  XOR2_X1 U462 ( .A(KEYINPUT96), .B(KEYINPUT9), .Z(n552) );
  XNOR2_X1 U463 ( .A(G122), .B(KEYINPUT7), .ZN(n551) );
  XOR2_X1 U464 ( .A(G116), .B(G107), .Z(n550) );
  XOR2_X1 U465 ( .A(KEYINPUT94), .B(KEYINPUT12), .Z(n538) );
  XNOR2_X1 U466 ( .A(n480), .B(G137), .ZN(n496) );
  XNOR2_X1 U467 ( .A(KEYINPUT67), .B(G140), .ZN(n480) );
  NAND2_X1 U468 ( .A1(G237), .A2(G234), .ZN(n515) );
  NOR2_X1 U469 ( .A1(n695), .A2(n477), .ZN(n476) );
  INV_X1 U470 ( .A(n651), .ZN(n477) );
  INV_X1 U471 ( .A(KEYINPUT39), .ZN(n448) );
  OR2_X1 U472 ( .A1(n717), .A2(n448), .ZN(n447) );
  INV_X1 U473 ( .A(n401), .ZN(n397) );
  NOR2_X1 U474 ( .A1(n705), .A2(n355), .ZN(n577) );
  NOR2_X1 U475 ( .A1(n613), .A2(n627), .ZN(n629) );
  NAND2_X1 U476 ( .A1(n601), .A2(n706), .ZN(n390) );
  XNOR2_X1 U477 ( .A(n512), .B(n522), .ZN(n472) );
  XNOR2_X1 U478 ( .A(n511), .B(n510), .ZN(n512) );
  INV_X1 U479 ( .A(KEYINPUT23), .ZN(n481) );
  XNOR2_X1 U480 ( .A(n405), .B(n403), .ZN(n450) );
  INV_X1 U481 ( .A(G110), .ZN(n403) );
  XNOR2_X1 U482 ( .A(n496), .B(n484), .ZN(n466) );
  INV_X1 U483 ( .A(KEYINPUT24), .ZN(n484) );
  INV_X1 U484 ( .A(n739), .ZN(n414) );
  NAND2_X1 U485 ( .A1(n433), .A2(n432), .ZN(n733) );
  INV_X1 U486 ( .A(KEYINPUT100), .ZN(n454) );
  NOR2_X1 U487 ( .A1(n388), .A2(n383), .ZN(n416) );
  INV_X1 U488 ( .A(KEYINPUT93), .ZN(n370) );
  NAND2_X1 U489 ( .A1(n372), .A2(n708), .ZN(n371) );
  XNOR2_X1 U490 ( .A(n629), .B(KEYINPUT92), .ZN(n372) );
  XNOR2_X1 U491 ( .A(n356), .B(n543), .ZN(n544) );
  XNOR2_X1 U492 ( .A(n766), .B(n503), .ZN(n661) );
  XNOR2_X1 U493 ( .A(G146), .B(KEYINPUT75), .ZN(n500) );
  XNOR2_X1 U494 ( .A(n411), .B(n531), .ZN(n668) );
  XNOR2_X1 U495 ( .A(n565), .B(n564), .ZN(n779) );
  NAND2_X1 U496 ( .A1(n358), .A2(n433), .ZN(n565) );
  NAND2_X1 U497 ( .A1(n394), .A2(n687), .ZN(n453) );
  AND2_X1 U498 ( .A1(n376), .A2(n375), .ZN(n579) );
  NAND2_X1 U499 ( .A1(n440), .A2(n462), .ZN(n439) );
  XNOR2_X1 U500 ( .A(n441), .B(KEYINPUT34), .ZN(n440) );
  XNOR2_X1 U501 ( .A(n626), .B(n381), .ZN(n691) );
  INV_X1 U502 ( .A(KEYINPUT31), .ZN(n381) );
  NOR2_X1 U503 ( .A1(n628), .A2(n712), .ZN(n626) );
  INV_X1 U504 ( .A(KEYINPUT77), .ZN(n377) );
  NOR2_X1 U505 ( .A1(n568), .A2(n567), .ZN(n378) );
  XNOR2_X1 U506 ( .A(n412), .B(KEYINPUT65), .ZN(n605) );
  NAND2_X1 U507 ( .A1(n374), .A2(n362), .ZN(n412) );
  AND2_X1 U508 ( .A1(n365), .A2(n701), .ZN(n393) );
  XNOR2_X1 U509 ( .A(n753), .B(n752), .ZN(n754) );
  INV_X1 U510 ( .A(KEYINPUT121), .ZN(n474) );
  INV_X1 U511 ( .A(n718), .ZN(n387) );
  OR2_X1 U512 ( .A1(n718), .A2(n478), .ZN(n354) );
  NAND2_X1 U513 ( .A1(n706), .A2(n364), .ZN(n355) );
  XOR2_X1 U514 ( .A(n541), .B(n540), .Z(n356) );
  AND2_X1 U515 ( .A1(n717), .A2(n431), .ZN(n357) );
  XNOR2_X1 U516 ( .A(n708), .B(n576), .ZN(n621) );
  AND2_X1 U517 ( .A1(n432), .A2(n436), .ZN(n358) );
  XOR2_X1 U518 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n359) );
  AND2_X1 U519 ( .A1(n548), .A2(G221), .ZN(n360) );
  AND2_X1 U520 ( .A1(n614), .A2(n577), .ZN(n361) );
  INV_X1 U521 ( .A(n570), .ZN(n470) );
  INV_X1 U522 ( .A(KEYINPUT30), .ZN(n478) );
  AND2_X1 U523 ( .A1(n701), .A2(n604), .ZN(n362) );
  XOR2_X1 U524 ( .A(KEYINPUT11), .B(KEYINPUT95), .Z(n363) );
  AND2_X1 U525 ( .A1(n597), .A2(n519), .ZN(n364) );
  AND2_X1 U526 ( .A1(n621), .A2(n430), .ZN(n365) );
  INV_X1 U527 ( .A(G902), .ZN(n460) );
  AND2_X1 U528 ( .A1(n469), .A2(n574), .ZN(n366) );
  XOR2_X1 U529 ( .A(KEYINPUT106), .B(KEYINPUT41), .Z(n367) );
  XOR2_X1 U530 ( .A(n602), .B(KEYINPUT68), .Z(n368) );
  XNOR2_X1 U531 ( .A(KEYINPUT82), .B(KEYINPUT45), .ZN(n369) );
  INV_X1 U532 ( .A(n426), .ZN(n675) );
  NAND2_X1 U533 ( .A1(n373), .A2(n414), .ZN(n697) );
  NAND2_X1 U534 ( .A1(n373), .A2(n739), .ZN(n743) );
  NAND2_X1 U535 ( .A1(n373), .A2(n771), .ZN(n762) );
  NAND2_X1 U536 ( .A1(n632), .A2(n373), .ZN(n634) );
  XNOR2_X2 U537 ( .A(n379), .B(n369), .ZN(n373) );
  NAND2_X1 U538 ( .A1(n374), .A2(n608), .ZN(n609) );
  AND2_X1 U539 ( .A1(n374), .A2(n393), .ZN(n673) );
  XNOR2_X2 U540 ( .A(n535), .B(n534), .ZN(n592) );
  INV_X1 U541 ( .A(n617), .ZN(n462) );
  NOR2_X1 U542 ( .A1(n615), .A2(n701), .ZN(n616) );
  INV_X1 U543 ( .A(n578), .ZN(n375) );
  NOR2_X1 U544 ( .A1(n408), .A2(n406), .ZN(n420) );
  AND2_X1 U545 ( .A1(n420), .A2(n778), .ZN(n417) );
  XNOR2_X1 U546 ( .A(n392), .B(KEYINPUT83), .ZN(n391) );
  NAND2_X1 U547 ( .A1(n391), .A2(n631), .ZN(n379) );
  NAND2_X1 U548 ( .A1(n426), .A2(n380), .ZN(n425) );
  XNOR2_X1 U549 ( .A(n415), .B(n464), .ZN(n419) );
  XNOR2_X1 U550 ( .A(n539), .B(n363), .ZN(n438) );
  XNOR2_X1 U551 ( .A(n438), .B(n404), .ZN(n545) );
  NAND2_X1 U552 ( .A1(n385), .A2(n384), .ZN(n383) );
  NOR2_X1 U553 ( .A1(n603), .A2(n478), .ZN(n388) );
  XNOR2_X2 U554 ( .A(n708), .B(KEYINPUT99), .ZN(n603) );
  NOR2_X1 U555 ( .A1(n613), .A2(n390), .ZN(n389) );
  NAND2_X1 U556 ( .A1(n394), .A2(n690), .ZN(n651) );
  NAND2_X1 U557 ( .A1(n753), .A2(n401), .ZN(n400) );
  NAND2_X1 U558 ( .A1(n397), .A2(n460), .ZN(n396) );
  NAND2_X1 U559 ( .A1(n401), .A2(G902), .ZN(n399) );
  INV_X1 U560 ( .A(n405), .ZN(n404) );
  XNOR2_X1 U561 ( .A(n766), .B(n405), .ZN(n770) );
  XNOR2_X2 U562 ( .A(n526), .B(KEYINPUT10), .ZN(n405) );
  NAND2_X1 U563 ( .A1(n407), .A2(n468), .ZN(n406) );
  INV_X1 U564 ( .A(n694), .ZN(n408) );
  NAND2_X1 U565 ( .A1(n409), .A2(n624), .ZN(n694) );
  XNOR2_X1 U566 ( .A(n579), .B(KEYINPUT36), .ZN(n409) );
  INV_X1 U567 ( .A(n705), .ZN(n622) );
  NAND2_X1 U568 ( .A1(n577), .A2(n603), .ZN(n410) );
  NAND2_X1 U569 ( .A1(n411), .A2(n758), .ZN(n759) );
  XNOR2_X2 U570 ( .A(n413), .B(n642), .ZN(n751) );
  NAND2_X1 U571 ( .A1(n640), .A2(n641), .ZN(n413) );
  NAND2_X1 U572 ( .A1(n605), .A2(n622), .ZN(n680) );
  XNOR2_X2 U573 ( .A(n507), .B(n472), .ZN(n643) );
  NAND2_X1 U574 ( .A1(n652), .A2(n779), .ZN(n415) );
  NAND2_X1 U575 ( .A1(n437), .A2(n476), .ZN(n475) );
  XNOR2_X1 U576 ( .A(n418), .B(n463), .ZN(n437) );
  NAND2_X1 U577 ( .A1(n419), .A2(n417), .ZN(n418) );
  XNOR2_X1 U578 ( .A(n587), .B(KEYINPUT104), .ZN(n778) );
  NAND2_X1 U579 ( .A1(n425), .A2(n570), .ZN(n429) );
  NAND2_X1 U580 ( .A1(n717), .A2(n718), .ZN(n721) );
  AND2_X1 U581 ( .A1(n437), .A2(n594), .ZN(n637) );
  XNOR2_X2 U582 ( .A(n485), .B(G146), .ZN(n526) );
  XNOR2_X2 U583 ( .A(n559), .B(n558), .ZN(n687) );
  XNOR2_X2 U584 ( .A(n439), .B(KEYINPUT35), .ZN(n775) );
  XNOR2_X2 U585 ( .A(n442), .B(n504), .ZN(n580) );
  NAND2_X1 U586 ( .A1(n582), .A2(KEYINPUT39), .ZN(n449) );
  INV_X1 U587 ( .A(n582), .ZN(n445) );
  XNOR2_X2 U588 ( .A(n487), .B(G902), .ZN(n638) );
  NAND2_X1 U589 ( .A1(n451), .A2(KEYINPUT80), .ZN(n573) );
  XNOR2_X1 U590 ( .A(n572), .B(n452), .ZN(n451) );
  XNOR2_X2 U591 ( .A(n453), .B(n561), .ZN(n652) );
  XNOR2_X1 U592 ( .A(n455), .B(n454), .ZN(n589) );
  NAND2_X1 U593 ( .A1(n588), .A2(n718), .ZN(n455) );
  NOR2_X1 U594 ( .A1(n643), .A2(n459), .ZN(n456) );
  XNOR2_X1 U595 ( .A(n657), .B(n474), .ZN(G63) );
  XNOR2_X2 U596 ( .A(n475), .B(KEYINPUT81), .ZN(n740) );
  XNOR2_X1 U597 ( .A(n747), .B(KEYINPUT59), .ZN(n479) );
  INV_X1 U598 ( .A(KEYINPUT84), .ZN(n610) );
  XNOR2_X1 U599 ( .A(n618), .B(n610), .ZN(n611) );
  XNOR2_X1 U600 ( .A(n482), .B(n481), .ZN(n483) );
  INV_X1 U601 ( .A(n757), .ZN(n648) );
  XNOR2_X1 U602 ( .A(n755), .B(n754), .ZN(n756) );
  XNOR2_X1 U603 ( .A(G128), .B(G119), .ZN(n482) );
  NAND2_X1 U604 ( .A1(n771), .A2(G234), .ZN(n486) );
  XOR2_X1 U605 ( .A(KEYINPUT8), .B(n486), .Z(n548) );
  XOR2_X1 U606 ( .A(KEYINPUT90), .B(KEYINPUT25), .Z(n490) );
  XNOR2_X2 U607 ( .A(KEYINPUT86), .B(KEYINPUT15), .ZN(n487) );
  NAND2_X1 U608 ( .A1(G234), .A2(n638), .ZN(n488) );
  NAND2_X1 U609 ( .A1(n491), .A2(G217), .ZN(n489) );
  NAND2_X1 U610 ( .A1(G221), .A2(n491), .ZN(n493) );
  XNOR2_X1 U611 ( .A(KEYINPUT91), .B(KEYINPUT21), .ZN(n492) );
  XNOR2_X1 U612 ( .A(n493), .B(n492), .ZN(n706) );
  XNOR2_X2 U613 ( .A(G143), .B(G128), .ZN(n527) );
  XNOR2_X1 U614 ( .A(n496), .B(KEYINPUT87), .ZN(n497) );
  NAND2_X1 U615 ( .A1(n771), .A2(G227), .ZN(n499) );
  XNOR2_X1 U616 ( .A(n499), .B(G101), .ZN(n501) );
  XNOR2_X1 U617 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U618 ( .A(n521), .B(n502), .ZN(n503) );
  INV_X1 U619 ( .A(G469), .ZN(n504) );
  INV_X1 U620 ( .A(n580), .ZN(n566) );
  NAND2_X1 U621 ( .A1(n623), .A2(n566), .ZN(n627) );
  INV_X1 U622 ( .A(KEYINPUT102), .ZN(n505) );
  XNOR2_X1 U623 ( .A(n627), .B(n505), .ZN(n520) );
  XOR2_X1 U624 ( .A(G101), .B(G119), .Z(n506) );
  XNOR2_X1 U625 ( .A(n508), .B(KEYINPUT74), .ZN(n542) );
  NAND2_X1 U626 ( .A1(n542), .A2(G210), .ZN(n511) );
  XNOR2_X1 U627 ( .A(n509), .B(KEYINPUT5), .ZN(n510) );
  INV_X1 U628 ( .A(G472), .ZN(n513) );
  XNOR2_X1 U629 ( .A(n514), .B(KEYINPUT71), .ZN(n532) );
  NAND2_X1 U630 ( .A1(n532), .A2(G214), .ZN(n718) );
  XNOR2_X1 U631 ( .A(n515), .B(KEYINPUT14), .ZN(n700) );
  NOR2_X1 U632 ( .A1(G902), .A2(n771), .ZN(n517) );
  NOR2_X1 U633 ( .A1(G953), .A2(G952), .ZN(n516) );
  NOR2_X1 U634 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X1 U635 ( .A1(n700), .A2(n518), .ZN(n597) );
  NAND2_X1 U636 ( .A1(G953), .A2(G900), .ZN(n519) );
  NAND2_X1 U637 ( .A1(G224), .A2(n771), .ZN(n524) );
  XNOR2_X1 U638 ( .A(n524), .B(KEYINPUT18), .ZN(n525) );
  XNOR2_X1 U639 ( .A(n526), .B(n525), .ZN(n530) );
  XNOR2_X1 U640 ( .A(n527), .B(n528), .ZN(n529) );
  XNOR2_X1 U641 ( .A(n530), .B(n529), .ZN(n531) );
  NAND2_X1 U642 ( .A1(n668), .A2(n638), .ZN(n535) );
  AND2_X1 U643 ( .A1(G210), .A2(n532), .ZN(n533) );
  INV_X1 U644 ( .A(KEYINPUT38), .ZN(n536) );
  XNOR2_X1 U645 ( .A(n592), .B(n536), .ZN(n717) );
  XNOR2_X1 U646 ( .A(KEYINPUT13), .B(G475), .ZN(n547) );
  XNOR2_X1 U647 ( .A(n538), .B(n537), .ZN(n539) );
  NAND2_X1 U648 ( .A1(G214), .A2(n542), .ZN(n543) );
  XNOR2_X1 U649 ( .A(n545), .B(n544), .ZN(n747) );
  NOR2_X1 U650 ( .A1(G902), .A2(n747), .ZN(n546) );
  NAND2_X1 U651 ( .A1(G217), .A2(n548), .ZN(n549) );
  XNOR2_X1 U652 ( .A(n550), .B(n549), .ZN(n556) );
  XNOR2_X1 U653 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U654 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U655 ( .A(n556), .B(n555), .ZN(n653) );
  NAND2_X1 U656 ( .A1(n653), .A2(n460), .ZN(n557) );
  XNOR2_X1 U657 ( .A(n557), .B(G478), .ZN(n584) );
  INV_X1 U658 ( .A(n584), .ZN(n569) );
  INV_X1 U659 ( .A(KEYINPUT97), .ZN(n558) );
  INV_X1 U660 ( .A(KEYINPUT105), .ZN(n560) );
  XNOR2_X1 U661 ( .A(n560), .B(KEYINPUT40), .ZN(n561) );
  NOR2_X1 U662 ( .A1(n584), .A2(n585), .ZN(n562) );
  XNOR2_X1 U663 ( .A(n562), .B(KEYINPUT98), .ZN(n601) );
  INV_X1 U664 ( .A(n601), .ZN(n720) );
  INV_X1 U665 ( .A(KEYINPUT107), .ZN(n563) );
  XNOR2_X1 U666 ( .A(n563), .B(KEYINPUT42), .ZN(n564) );
  NAND2_X1 U667 ( .A1(n599), .A2(n566), .ZN(n567) );
  NOR2_X1 U668 ( .A1(n585), .A2(n569), .ZN(n690) );
  NOR2_X1 U669 ( .A1(n687), .A2(n690), .ZN(n722) );
  INV_X1 U670 ( .A(n722), .ZN(n570) );
  XNOR2_X1 U671 ( .A(KEYINPUT66), .B(KEYINPUT47), .ZN(n571) );
  NAND2_X1 U672 ( .A1(n573), .A2(n685), .ZN(n575) );
  OR2_X1 U673 ( .A1(KEYINPUT80), .A2(KEYINPUT47), .ZN(n574) );
  INV_X1 U674 ( .A(KEYINPUT6), .ZN(n576) );
  INV_X1 U675 ( .A(n621), .ZN(n614) );
  INV_X1 U676 ( .A(n701), .ZN(n624) );
  INV_X1 U677 ( .A(n592), .ZN(n581) );
  NOR2_X1 U678 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U679 ( .A(n583), .B(KEYINPUT103), .ZN(n586) );
  NAND2_X1 U680 ( .A1(n585), .A2(n584), .ZN(n617) );
  OR2_X1 U681 ( .A1(n586), .A2(n617), .ZN(n587) );
  AND2_X1 U682 ( .A1(n589), .A2(n701), .ZN(n591) );
  XOR2_X1 U683 ( .A(KEYINPUT101), .B(KEYINPUT43), .Z(n590) );
  XNOR2_X1 U684 ( .A(n591), .B(n590), .ZN(n593) );
  NOR2_X1 U685 ( .A1(n593), .A2(n592), .ZN(n695) );
  INV_X1 U686 ( .A(n695), .ZN(n594) );
  INV_X1 U687 ( .A(KEYINPUT73), .ZN(n595) );
  XNOR2_X1 U688 ( .A(n740), .B(n595), .ZN(n632) );
  NAND2_X1 U689 ( .A1(G898), .A2(G953), .ZN(n596) );
  AND2_X1 U690 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U691 ( .A1(n599), .A2(n598), .ZN(n600) );
  INV_X1 U692 ( .A(n603), .ZN(n604) );
  NAND2_X1 U693 ( .A1(n624), .A2(n621), .ZN(n606) );
  NOR2_X1 U694 ( .A1(n705), .A2(n606), .ZN(n607) );
  XNOR2_X1 U695 ( .A(KEYINPUT76), .B(n607), .ZN(n608) );
  XNOR2_X1 U696 ( .A(n609), .B(KEYINPUT32), .ZN(n777) );
  NAND2_X1 U697 ( .A1(n680), .A2(n777), .ZN(n612) );
  INV_X1 U698 ( .A(KEYINPUT44), .ZN(n618) );
  XNOR2_X1 U699 ( .A(n612), .B(n611), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n623), .A2(n614), .ZN(n615) );
  XNOR2_X1 U701 ( .A(KEYINPUT33), .B(n616), .ZN(n732) );
  NAND2_X1 U702 ( .A1(n618), .A2(n775), .ZN(n619) );
  NAND2_X1 U703 ( .A1(n620), .A2(n619), .ZN(n631) );
  INV_X1 U704 ( .A(n623), .ZN(n702) );
  NOR2_X1 U705 ( .A1(n702), .A2(n708), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n625), .A2(n624), .ZN(n712) );
  NAND2_X1 U707 ( .A1(n775), .A2(KEYINPUT44), .ZN(n630) );
  INV_X1 U708 ( .A(KEYINPUT2), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n634), .A2(n633), .ZN(n641) );
  NAND2_X1 U710 ( .A1(n651), .A2(KEYINPUT2), .ZN(n635) );
  XNOR2_X1 U711 ( .A(n635), .B(KEYINPUT79), .ZN(n636) );
  NAND2_X1 U712 ( .A1(n637), .A2(n636), .ZN(n739) );
  INV_X1 U713 ( .A(n638), .ZN(n639) );
  NAND2_X1 U714 ( .A1(n751), .A2(G472), .ZN(n645) );
  XNOR2_X1 U715 ( .A(n643), .B(KEYINPUT62), .ZN(n644) );
  XNOR2_X1 U716 ( .A(n645), .B(n644), .ZN(n646) );
  INV_X1 U717 ( .A(n646), .ZN(n649) );
  INV_X1 U718 ( .A(G952), .ZN(n647) );
  AND2_X1 U719 ( .A1(n647), .A2(G953), .ZN(n757) );
  NAND2_X1 U720 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U721 ( .A(n650), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U722 ( .A(n651), .B(G134), .ZN(G36) );
  XNOR2_X1 U723 ( .A(n652), .B(G131), .ZN(G33) );
  NAND2_X1 U724 ( .A1(n751), .A2(G478), .ZN(n655) );
  INV_X1 U725 ( .A(n653), .ZN(n654) );
  XNOR2_X1 U726 ( .A(n655), .B(n654), .ZN(n656) );
  NOR2_X2 U727 ( .A1(n656), .A2(n757), .ZN(n657) );
  NAND2_X1 U728 ( .A1(n751), .A2(G469), .ZN(n663) );
  XNOR2_X1 U729 ( .A(KEYINPUT120), .B(KEYINPUT57), .ZN(n659) );
  XNOR2_X1 U730 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n658) );
  XNOR2_X1 U731 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U732 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U733 ( .A(n663), .B(n662), .ZN(n664) );
  NOR2_X1 U734 ( .A1(n664), .A2(n757), .ZN(G54) );
  NAND2_X1 U735 ( .A1(n751), .A2(G210), .ZN(n670) );
  XOR2_X1 U736 ( .A(KEYINPUT118), .B(KEYINPUT54), .Z(n666) );
  XNOR2_X1 U737 ( .A(KEYINPUT55), .B(KEYINPUT85), .ZN(n665) );
  XNOR2_X1 U738 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U739 ( .A(n670), .B(n669), .ZN(n671) );
  NOR2_X2 U740 ( .A1(n671), .A2(n757), .ZN(n672) );
  XNOR2_X1 U741 ( .A(n672), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U742 ( .A(G101), .B(n673), .Z(G3) );
  NAND2_X1 U743 ( .A1(n675), .A2(n687), .ZN(n674) );
  XNOR2_X1 U744 ( .A(n674), .B(G104), .ZN(G6) );
  XOR2_X1 U745 ( .A(KEYINPUT26), .B(KEYINPUT27), .Z(n677) );
  NAND2_X1 U746 ( .A1(n675), .A2(n690), .ZN(n676) );
  XNOR2_X1 U747 ( .A(n677), .B(n676), .ZN(n679) );
  XOR2_X1 U748 ( .A(G107), .B(KEYINPUT109), .Z(n678) );
  XNOR2_X1 U749 ( .A(n679), .B(n678), .ZN(G9) );
  XNOR2_X1 U750 ( .A(n680), .B(G110), .ZN(G12) );
  XOR2_X1 U751 ( .A(KEYINPUT29), .B(KEYINPUT111), .Z(n682) );
  NAND2_X1 U752 ( .A1(n685), .A2(n690), .ZN(n681) );
  XNOR2_X1 U753 ( .A(n682), .B(n681), .ZN(n684) );
  XOR2_X1 U754 ( .A(G128), .B(KEYINPUT110), .Z(n683) );
  XNOR2_X1 U755 ( .A(n684), .B(n683), .ZN(G30) );
  NAND2_X1 U756 ( .A1(n685), .A2(n687), .ZN(n686) );
  XNOR2_X1 U757 ( .A(n686), .B(G146), .ZN(G48) );
  NAND2_X1 U758 ( .A1(n691), .A2(n687), .ZN(n688) );
  XNOR2_X1 U759 ( .A(n688), .B(KEYINPUT112), .ZN(n689) );
  XNOR2_X1 U760 ( .A(G113), .B(n689), .ZN(G15) );
  NAND2_X1 U761 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U762 ( .A(n692), .B(G116), .ZN(G18) );
  XOR2_X1 U763 ( .A(G125), .B(KEYINPUT37), .Z(n693) );
  XNOR2_X1 U764 ( .A(n694), .B(n693), .ZN(G27) );
  XNOR2_X1 U765 ( .A(G140), .B(n695), .ZN(n696) );
  XNOR2_X1 U766 ( .A(n696), .B(KEYINPUT113), .ZN(G42) );
  INV_X1 U767 ( .A(n697), .ZN(n698) );
  NOR2_X1 U768 ( .A1(n698), .A2(n633), .ZN(n699) );
  NOR2_X1 U769 ( .A1(G953), .A2(n699), .ZN(n738) );
  NAND2_X1 U770 ( .A1(G952), .A2(n700), .ZN(n731) );
  NAND2_X1 U771 ( .A1(n702), .A2(n701), .ZN(n704) );
  XNOR2_X1 U772 ( .A(KEYINPUT114), .B(KEYINPUT50), .ZN(n703) );
  XNOR2_X1 U773 ( .A(n704), .B(n703), .ZN(n711) );
  NOR2_X1 U774 ( .A1(n706), .A2(n430), .ZN(n707) );
  XNOR2_X1 U775 ( .A(KEYINPUT49), .B(n707), .ZN(n709) );
  AND2_X1 U776 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U777 ( .A1(n711), .A2(n710), .ZN(n713) );
  NAND2_X1 U778 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U779 ( .A(n714), .B(KEYINPUT115), .Z(n715) );
  XNOR2_X1 U780 ( .A(KEYINPUT51), .B(n715), .ZN(n716) );
  NOR2_X1 U781 ( .A1(n733), .A2(n716), .ZN(n728) );
  NOR2_X1 U782 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U783 ( .A1(n720), .A2(n719), .ZN(n725) );
  NOR2_X1 U784 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U785 ( .A(n723), .B(KEYINPUT116), .ZN(n724) );
  NOR2_X1 U786 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U787 ( .A1(n726), .A2(n732), .ZN(n727) );
  NOR2_X1 U788 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U789 ( .A(n729), .B(KEYINPUT52), .ZN(n730) );
  NOR2_X1 U790 ( .A1(n731), .A2(n730), .ZN(n735) );
  NOR2_X1 U791 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U792 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U793 ( .A(KEYINPUT117), .B(n736), .Z(n737) );
  NAND2_X1 U794 ( .A1(n738), .A2(n737), .ZN(n745) );
  BUF_X1 U795 ( .A(n740), .Z(n741) );
  INV_X1 U796 ( .A(n741), .ZN(n742) );
  NOR2_X1 U797 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U798 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U799 ( .A(KEYINPUT53), .B(n746), .ZN(G75) );
  NAND2_X1 U800 ( .A1(n751), .A2(G475), .ZN(n748) );
  XNOR2_X1 U801 ( .A(n748), .B(n479), .ZN(n749) );
  XNOR2_X1 U802 ( .A(n750), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U803 ( .A1(n751), .A2(G217), .ZN(n755) );
  XOR2_X1 U804 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n752) );
  NOR2_X1 U805 ( .A1(n757), .A2(n756), .ZN(G66) );
  OR2_X1 U806 ( .A1(G898), .A2(n771), .ZN(n758) );
  XNOR2_X1 U807 ( .A(n759), .B(KEYINPUT124), .ZN(n765) );
  NAND2_X1 U808 ( .A1(G953), .A2(G224), .ZN(n760) );
  XNOR2_X1 U809 ( .A(KEYINPUT61), .B(n760), .ZN(n761) );
  NAND2_X1 U810 ( .A1(n761), .A2(G898), .ZN(n763) );
  NAND2_X1 U811 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U812 ( .A(n765), .B(n764), .Z(G69) );
  XOR2_X1 U813 ( .A(G227), .B(n770), .Z(n767) );
  NAND2_X1 U814 ( .A1(n767), .A2(G900), .ZN(n768) );
  NAND2_X1 U815 ( .A1(n768), .A2(G953), .ZN(n769) );
  XOR2_X1 U816 ( .A(KEYINPUT125), .B(n769), .Z(n774) );
  XNOR2_X1 U817 ( .A(n741), .B(n770), .ZN(n772) );
  NAND2_X1 U818 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U819 ( .A1(n774), .A2(n773), .ZN(G72) );
  XOR2_X1 U820 ( .A(n775), .B(G122), .Z(n776) );
  XNOR2_X1 U821 ( .A(KEYINPUT126), .B(n776), .ZN(G24) );
  XNOR2_X1 U822 ( .A(G119), .B(n777), .ZN(G21) );
  XNOR2_X1 U823 ( .A(G143), .B(n778), .ZN(G45) );
  XNOR2_X1 U824 ( .A(G137), .B(n779), .ZN(G39) );
endmodule

