//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 1 1 0 0 0 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  INV_X1    g000(.A(KEYINPUT64), .ZN(new_n187));
  INV_X1    g001(.A(G137), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT64), .A2(G137), .ZN(new_n190));
  AND2_X1   g004(.A1(KEYINPUT11), .A2(G134), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(new_n190), .A3(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT11), .ZN(new_n193));
  INV_X1    g007(.A(G134), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G137), .ZN(new_n195));
  AOI21_X1  g009(.A(G131), .B1(new_n194), .B2(G137), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n192), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT65), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n192), .A2(new_n199), .A3(new_n195), .A4(new_n196), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n192), .B(new_n195), .C1(G134), .C2(new_n188), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G131), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G143), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  AND2_X1   g022(.A1(KEYINPUT0), .A2(G128), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(G143), .B(G146), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT0), .B(G128), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n204), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT1), .B1(new_n207), .B2(G146), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n207), .A2(G146), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n205), .A2(G143), .ZN(new_n218));
  OAI211_X1 g032(.A(G128), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G128), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n206), .B(new_n208), .C1(KEYINPUT1), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n224), .B1(new_n194), .B2(G137), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n188), .A2(KEYINPUT66), .A3(G134), .ZN(new_n226));
  AND2_X1   g040(.A1(KEYINPUT64), .A2(G137), .ZN(new_n227));
  NOR2_X1   g041(.A1(KEYINPUT64), .A2(G137), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n225), .B(new_n226), .C1(new_n229), .C2(G134), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n198), .A2(new_n200), .B1(G131), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n223), .B1(new_n231), .B2(KEYINPUT67), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(G131), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n201), .A2(KEYINPUT67), .A3(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n215), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT72), .ZN(new_n236));
  INV_X1    g050(.A(G119), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G116), .ZN(new_n238));
  INV_X1    g052(.A(G116), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G119), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n238), .A2(new_n240), .A3(KEYINPUT68), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT2), .B(G113), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  OR2_X1    g060(.A1(new_n241), .A2(new_n245), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n235), .A2(new_n236), .A3(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT71), .B(KEYINPUT28), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n235), .A2(new_n248), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT11), .B1(new_n188), .B2(G134), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n252), .B1(new_n229), .B2(new_n191), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n199), .B1(new_n253), .B2(new_n196), .ZN(new_n254));
  INV_X1    g068(.A(new_n200), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n223), .B(new_n233), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n248), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n198), .A2(new_n200), .B1(G131), .B2(new_n202), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n213), .A2(KEYINPUT69), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n210), .B(new_n260), .C1(new_n211), .C2(new_n212), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n256), .B(new_n257), .C1(new_n258), .C2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT72), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n249), .B(new_n250), .C1(new_n251), .C2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT28), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n263), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n266), .B1(new_n263), .B2(new_n267), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G237), .ZN(new_n271));
  INV_X1    g085(.A(G953), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(G210), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n273), .B(KEYINPUT27), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(G101), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n274), .B(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n265), .A2(new_n270), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT29), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT30), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n279), .B(new_n215), .C1(new_n232), .C2(new_n234), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n256), .B1(new_n258), .B2(new_n262), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT30), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n248), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n263), .ZN(new_n285));
  INV_X1    g099(.A(new_n276), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n277), .A2(new_n278), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n263), .A2(KEYINPUT76), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n204), .A2(new_n261), .A3(new_n259), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT76), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n291), .A2(new_n292), .A3(new_n257), .A4(new_n256), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n281), .A2(new_n248), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n290), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n270), .B1(new_n296), .B2(new_n267), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n276), .A2(KEYINPUT29), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n289), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G472), .B1(new_n288), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT31), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT70), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n263), .A2(new_n302), .A3(new_n276), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n302), .B1(new_n263), .B2(new_n276), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n257), .B1(new_n280), .B2(new_n282), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n301), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n263), .A2(new_n276), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT70), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n263), .A2(new_n302), .A3(new_n276), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n284), .A2(new_n311), .A3(KEYINPUT31), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n249), .A2(new_n250), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n264), .B1(new_n248), .B2(new_n235), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n270), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AOI22_X1  g129(.A1(new_n307), .A2(new_n312), .B1(new_n315), .B2(new_n286), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(G472), .A2(G902), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(KEYINPUT32), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n300), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n321));
  INV_X1    g135(.A(new_n318), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n321), .B1(new_n316), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT32), .ZN(new_n324));
  NOR3_X1   g138(.A1(new_n305), .A2(new_n306), .A3(new_n301), .ZN(new_n325));
  AOI21_X1  g139(.A(KEYINPUT31), .B1(new_n284), .B2(new_n311), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n276), .B1(new_n265), .B2(new_n270), .ZN(new_n328));
  OAI211_X1 g142(.A(KEYINPUT74), .B(new_n318), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n323), .A2(new_n324), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n323), .A2(new_n329), .A3(KEYINPUT75), .A4(new_n324), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n320), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(G214), .B1(G237), .B2(G902), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT94), .ZN(new_n337));
  INV_X1    g151(.A(G122), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n337), .B1(G116), .B2(new_n338), .ZN(new_n339));
  NOR3_X1   g153(.A1(new_n239), .A2(KEYINPUT94), .A3(G122), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G107), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n239), .A2(G122), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n344), .B(KEYINPUT14), .ZN(new_n346));
  OAI21_X1  g160(.A(G107), .B1(new_n346), .B2(new_n341), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n207), .A2(G128), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n220), .A2(G143), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n350), .B(G134), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n345), .A2(new_n347), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT95), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT95), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n345), .A2(new_n347), .A3(new_n354), .A4(new_n351), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n342), .A2(new_n344), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G107), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n345), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT13), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n194), .B1(new_n349), .B2(new_n360), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n361), .A2(new_n350), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n350), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n359), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT9), .B(G234), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(G217), .A3(new_n272), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n356), .A2(new_n364), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n368), .B1(new_n356), .B2(new_n364), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n289), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G478), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(KEYINPUT15), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n356), .A2(new_n364), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n367), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n356), .A2(new_n364), .A3(new_n368), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n373), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n289), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n374), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(G113), .B(G122), .ZN(new_n383));
  INV_X1    g197(.A(G104), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n383), .B(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n271), .A2(new_n272), .A3(G214), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n207), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n271), .A2(new_n272), .A3(G143), .A4(G214), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G131), .ZN(new_n390));
  INV_X1    g204(.A(G131), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n387), .A2(new_n391), .A3(new_n388), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(G125), .B(G140), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT16), .ZN(new_n395));
  INV_X1    g209(.A(G125), .ZN(new_n396));
  OR2_X1    g210(.A1(new_n396), .A2(G140), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n395), .B(G146), .C1(KEYINPUT16), .C2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT19), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n394), .B(new_n399), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n393), .B(new_n398), .C1(G146), .C2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n394), .A2(new_n205), .ZN(new_n402));
  INV_X1    g216(.A(new_n394), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G146), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT92), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n387), .A2(new_n405), .A3(new_n388), .ZN(new_n406));
  NAND2_X1  g220(.A1(KEYINPUT18), .A2(G131), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  AOI22_X1  g222(.A1(new_n402), .A2(new_n404), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  OR2_X1    g223(.A1(new_n406), .A2(new_n408), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n385), .B1(new_n401), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n395), .B1(KEYINPUT16), .B2(new_n397), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n205), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n389), .A2(KEYINPUT17), .A3(G131), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n414), .A2(new_n415), .A3(new_n398), .ZN(new_n416));
  OR2_X1    g230(.A1(new_n393), .A2(KEYINPUT17), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n416), .A2(new_n417), .B1(new_n410), .B2(new_n409), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n412), .B1(new_n418), .B2(new_n385), .ZN(new_n419));
  NOR2_X1   g233(.A1(G475), .A2(G902), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n420), .B(KEYINPUT93), .ZN(new_n421));
  OAI21_X1  g235(.A(KEYINPUT20), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n416), .A2(new_n417), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(new_n385), .A3(new_n411), .ZN(new_n424));
  INV_X1    g238(.A(new_n412), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT20), .ZN(new_n427));
  INV_X1    g241(.A(new_n421), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n424), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n418), .A2(new_n385), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n289), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n422), .A2(new_n429), .B1(new_n432), .B2(G475), .ZN(new_n433));
  INV_X1    g247(.A(G952), .ZN(new_n434));
  AOI211_X1 g248(.A(G953), .B(new_n434), .C1(G234), .C2(G237), .ZN(new_n435));
  AOI211_X1 g249(.A(new_n289), .B(new_n272), .C1(G234), .C2(G237), .ZN(new_n436));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(G898), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n382), .A2(new_n433), .A3(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(G210), .B1(G237), .B2(G902), .ZN(new_n441));
  XOR2_X1   g255(.A(new_n441), .B(KEYINPUT91), .Z(new_n442));
  NAND2_X1  g256(.A1(new_n272), .A2(G224), .ZN(new_n443));
  XOR2_X1   g257(.A(new_n443), .B(KEYINPUT89), .Z(new_n444));
  NAND2_X1  g258(.A1(new_n213), .A2(G125), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT86), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n445), .B(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT87), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n445), .B(KEYINPUT86), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT87), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n222), .A2(new_n396), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT88), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n453), .B(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n444), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n453), .B(KEYINPUT88), .ZN(new_n457));
  INV_X1    g271(.A(new_n444), .ZN(new_n458));
  AOI211_X1 g272(.A(new_n457), .B(new_n458), .C1(new_n448), .C2(new_n451), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(G110), .B(G122), .ZN(new_n461));
  OAI21_X1  g275(.A(KEYINPUT3), .B1(new_n384), .B2(G107), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT3), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(new_n343), .A3(G104), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n384), .A2(G107), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(G101), .ZN(new_n467));
  INV_X1    g281(.A(G101), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n462), .A2(new_n464), .A3(new_n468), .A4(new_n465), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(KEYINPUT4), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT4), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n466), .A2(new_n471), .A3(G101), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n248), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT84), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n384), .A2(G107), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n343), .A2(G104), .ZN(new_n477));
  OAI21_X1  g291(.A(G101), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n469), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT5), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n481), .B1(new_n243), .B2(new_n244), .ZN(new_n482));
  OAI21_X1  g296(.A(G113), .B1(new_n238), .B2(KEYINPUT5), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n480), .B(new_n247), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n248), .A2(KEYINPUT84), .A3(new_n470), .A4(new_n472), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n475), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT85), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n461), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n475), .A2(KEYINPUT85), .A3(new_n484), .A4(new_n485), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n475), .A2(new_n484), .A3(new_n485), .A4(new_n461), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT6), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n488), .A2(KEYINPUT6), .A3(new_n489), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n460), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n455), .A2(new_n449), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n443), .A2(KEYINPUT7), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n247), .B(new_n479), .C1(new_n482), .C2(new_n483), .ZN(new_n498));
  XOR2_X1   g312(.A(new_n461), .B(KEYINPUT8), .Z(new_n499));
  NOR2_X1   g313(.A1(new_n241), .A2(new_n481), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n247), .B1(new_n500), .B2(new_n483), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n499), .B1(new_n501), .B2(new_n480), .ZN(new_n502));
  AOI22_X1  g316(.A1(new_n496), .A2(new_n497), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n452), .A2(new_n455), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT7), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT90), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n505), .B1(new_n443), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n507), .B1(new_n506), .B2(new_n443), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n503), .B(new_n491), .C1(new_n504), .C2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n289), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n442), .B1(new_n495), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n494), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n488), .A2(new_n489), .B1(KEYINPUT6), .B2(new_n491), .ZN(new_n513));
  OAI22_X1  g327(.A1(new_n512), .A2(new_n513), .B1(new_n459), .B2(new_n456), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n514), .A2(new_n289), .A3(new_n441), .A4(new_n509), .ZN(new_n515));
  AOI211_X1 g329(.A(new_n336), .B(new_n440), .C1(new_n511), .C2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(G221), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n517), .B1(new_n366), .B2(new_n289), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT12), .ZN(new_n519));
  OR2_X1    g333(.A1(new_n519), .A2(KEYINPUT80), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(KEYINPUT80), .ZN(new_n521));
  AND4_X1   g335(.A1(new_n221), .A2(new_n219), .A3(new_n469), .A4(new_n478), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n221), .A2(new_n219), .B1(new_n469), .B2(new_n478), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n520), .B(new_n521), .C1(new_n524), .C2(new_n258), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n222), .A2(new_n479), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n219), .A2(new_n469), .A3(new_n478), .A4(new_n221), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n204), .A2(KEYINPUT80), .A3(new_n519), .A4(new_n528), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT10), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n527), .B(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT79), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n259), .A2(new_n261), .A3(new_n472), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n534), .B1(new_n535), .B2(new_n470), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n259), .A2(new_n261), .A3(new_n472), .ZN(new_n537));
  INV_X1    g351(.A(new_n470), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT79), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n258), .B(new_n533), .C1(new_n536), .C2(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(G110), .B(G140), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n272), .A2(G227), .ZN(new_n542));
  XOR2_X1   g356(.A(new_n541), .B(new_n542), .Z(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n530), .A2(new_n540), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT82), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n535), .A2(new_n534), .A3(new_n470), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT79), .B1(new_n537), .B2(new_n538), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n532), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n550), .A2(new_n258), .ZN(new_n551));
  AOI211_X1 g365(.A(new_n204), .B(new_n532), .C1(new_n548), .C2(new_n549), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n543), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n530), .A2(new_n540), .A3(KEYINPUT82), .A4(new_n544), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n547), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  XOR2_X1   g369(.A(KEYINPUT81), .B(G469), .Z(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n289), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT83), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n555), .A2(KEYINPUT83), .A3(new_n289), .A4(new_n556), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OR2_X1    g375(.A1(new_n550), .A2(new_n258), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n543), .B1(new_n550), .B2(new_n258), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n530), .A2(new_n540), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n543), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(G469), .B1(new_n567), .B2(G902), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n518), .B1(new_n561), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n516), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT23), .B1(new_n220), .B2(G119), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT77), .B1(new_n237), .B2(G128), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n571), .B(new_n572), .Z(new_n573));
  XNOR2_X1  g387(.A(G119), .B(G128), .ZN(new_n574));
  XOR2_X1   g388(.A(KEYINPUT24), .B(G110), .Z(new_n575));
  OAI22_X1  g389(.A1(new_n573), .A2(G110), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(new_n398), .A3(new_n402), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n414), .A2(new_n398), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n575), .A2(new_n574), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n573), .A2(G110), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT22), .B(G137), .ZN(new_n583));
  INV_X1    g397(.A(G234), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n517), .A2(new_n584), .A3(G953), .ZN(new_n585));
  XOR2_X1   g399(.A(new_n583), .B(new_n585), .Z(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n577), .A2(new_n581), .A3(new_n586), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n588), .A2(new_n289), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT78), .ZN(new_n591));
  AOI21_X1  g405(.A(KEYINPUT25), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(G217), .B1(new_n584), .B2(G902), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n590), .A2(new_n591), .A3(KEYINPUT25), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n588), .A2(new_n589), .ZN(new_n597));
  AOI21_X1  g411(.A(G902), .B1(new_n584), .B2(G217), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n334), .A2(new_n570), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(new_n468), .ZN(G3));
  INV_X1    g416(.A(new_n569), .ZN(new_n603));
  OAI21_X1  g417(.A(G472), .B1(new_n316), .B2(G902), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n323), .A2(new_n604), .A3(new_n329), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n603), .A2(new_n600), .A3(new_n605), .ZN(new_n606));
  MUX2_X1   g420(.A(new_n289), .B(new_n371), .S(new_n372), .Z(new_n607));
  NAND2_X1  g421(.A1(new_n378), .A2(KEYINPUT33), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT33), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n376), .A2(new_n609), .A3(new_n377), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n608), .A2(G478), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n612), .A2(new_n433), .A3(new_n438), .ZN(new_n613));
  INV_X1    g427(.A(new_n441), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n614), .B1(new_n495), .B2(new_n510), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n336), .B1(new_n615), .B2(new_n515), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n606), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT34), .B(G104), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT98), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n617), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G6));
  NAND3_X1  g436(.A1(new_n422), .A2(new_n429), .A3(KEYINPUT99), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT99), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n624), .B(KEYINPUT20), .C1(new_n419), .C2(new_n421), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n432), .A2(G475), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n623), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  AND4_X1   g442(.A1(new_n381), .A2(new_n616), .A3(new_n439), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n606), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT35), .B(G107), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  NOR2_X1   g446(.A1(new_n587), .A2(KEYINPUT36), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n582), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n598), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n596), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n637), .A2(new_n440), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n511), .A2(new_n515), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n638), .A2(new_n335), .A3(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n603), .A2(new_n640), .A3(new_n605), .ZN(new_n641));
  XNOR2_X1  g455(.A(KEYINPUT37), .B(G110), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G12));
  NAND2_X1  g457(.A1(new_n332), .A2(new_n333), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n300), .A2(new_n319), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(G900), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n435), .B1(new_n436), .B2(new_n647), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n382), .A2(new_n627), .A3(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n569), .A2(new_n616), .A3(new_n636), .A4(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n646), .A2(KEYINPUT100), .A3(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n653), .B1(new_n334), .B2(new_n650), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G128), .ZN(G30));
  XOR2_X1   g470(.A(new_n648), .B(KEYINPUT39), .Z(new_n657));
  NAND2_X1  g471(.A1(new_n569), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(KEYINPUT40), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT38), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n511), .A2(new_n515), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n660), .B1(new_n511), .B2(new_n515), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n382), .A2(new_n433), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n637), .A2(new_n335), .A3(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n659), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n319), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n284), .A2(new_n311), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n668), .B1(new_n296), .B2(new_n276), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n289), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n667), .B1(G472), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n644), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n658), .A2(KEYINPUT40), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n666), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT101), .B(G143), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G45));
  NOR3_X1   g490(.A1(new_n612), .A2(new_n433), .A3(new_n648), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n569), .A2(new_n616), .A3(new_n636), .A4(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n334), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(new_n205), .ZN(G48));
  AOI21_X1  g494(.A(new_n600), .B1(new_n644), .B2(new_n645), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n555), .A2(new_n289), .ZN(new_n682));
  AOI22_X1  g496(.A1(new_n559), .A2(new_n560), .B1(G469), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n518), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n683), .A2(new_n616), .A3(new_n684), .A4(new_n613), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(KEYINPUT102), .B1(new_n681), .B2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT102), .ZN(new_n688));
  NOR4_X1   g502(.A1(new_n334), .A2(new_n688), .A3(new_n600), .A4(new_n685), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT41), .B(G113), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G15));
  NAND2_X1  g506(.A1(new_n682), .A2(G469), .ZN(new_n693));
  AND3_X1   g507(.A1(new_n561), .A2(new_n684), .A3(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n681), .A2(new_n629), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  AND3_X1   g510(.A1(new_n694), .A2(new_n616), .A3(new_n638), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n646), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G119), .ZN(G21));
  NAND2_X1  g513(.A1(new_n683), .A2(new_n684), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n297), .A2(new_n286), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n701), .B(new_n318), .C1(new_n702), .C2(new_n327), .ZN(new_n703));
  AOI22_X1  g517(.A1(new_n307), .A2(new_n312), .B1(new_n297), .B2(new_n286), .ZN(new_n704));
  OAI21_X1  g518(.A(KEYINPUT103), .B1(new_n704), .B2(new_n322), .ZN(new_n705));
  INV_X1    g519(.A(new_n600), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n703), .A2(new_n705), .A3(new_n604), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n616), .A2(new_n664), .ZN(new_n708));
  NOR4_X1   g522(.A1(new_n700), .A2(new_n707), .A3(new_n708), .A4(new_n438), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n338), .ZN(G24));
  NAND4_X1  g524(.A1(new_n683), .A2(new_n616), .A3(new_n684), .A4(new_n677), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n703), .A2(new_n705), .A3(new_n604), .A4(new_n636), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n396), .ZN(G27));
  AOI21_X1  g528(.A(G902), .B1(new_n564), .B2(new_n566), .ZN(new_n715));
  INV_X1    g529(.A(G469), .ZN(new_n716));
  OAI21_X1  g530(.A(KEYINPUT104), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n716), .A2(KEYINPUT104), .A3(G902), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n567), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n561), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n722), .A3(new_n684), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n559), .A2(new_n560), .B1(new_n717), .B2(new_n719), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT105), .B1(new_n724), .B2(new_n518), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n511), .A2(new_n515), .A3(new_n335), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n723), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n677), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(KEYINPUT42), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n728), .A2(new_n646), .A3(new_n706), .A4(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n324), .B1(new_n316), .B2(new_n322), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n645), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n706), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n723), .A2(new_n725), .A3(new_n677), .A4(new_n727), .ZN(new_n735));
  OAI21_X1  g549(.A(KEYINPUT42), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G131), .ZN(G33));
  NAND3_X1  g552(.A1(new_n681), .A2(new_n649), .A3(new_n728), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G134), .ZN(G36));
  NAND2_X1  g554(.A1(G469), .A2(G902), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n564), .A2(new_n566), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(G469), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n742), .A2(new_n743), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n741), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT46), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n567), .A2(KEYINPUT45), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(G469), .A3(new_n744), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(KEYINPUT46), .A3(new_n741), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n749), .A2(new_n561), .A3(new_n752), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n753), .A2(new_n684), .A3(new_n657), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n607), .A2(new_n433), .A3(new_n611), .ZN(new_n755));
  XOR2_X1   g569(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n607), .A2(new_n433), .A3(new_n611), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n605), .A2(new_n762), .A3(KEYINPUT44), .A4(new_n636), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT44), .ZN(new_n764));
  INV_X1    g578(.A(new_n605), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n762), .A2(new_n636), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n754), .A2(new_n727), .A3(new_n763), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G137), .ZN(G39));
  NOR3_X1   g583(.A1(new_n729), .A2(new_n706), .A3(new_n726), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n753), .A2(KEYINPUT47), .A3(new_n684), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT47), .B1(new_n753), .B2(new_n684), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n334), .B(new_n770), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(KEYINPUT107), .B(G140), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(G42));
  INV_X1    g589(.A(new_n672), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n600), .A2(new_n755), .A3(new_n518), .A4(new_n336), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n663), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n683), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n778), .B1(KEYINPUT49), .B2(new_n779), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n776), .B(new_n780), .C1(KEYINPUT49), .C2(new_n779), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n782));
  AOI211_X1 g596(.A(new_n336), .B(new_n438), .C1(new_n511), .C2(new_n515), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n765), .A2(new_n569), .A3(new_n706), .A4(new_n783), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n784), .A2(new_n433), .A3(new_n612), .ZN(new_n785));
  OAI21_X1  g599(.A(KEYINPUT108), .B1(new_n601), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n433), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n784), .A2(new_n382), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n641), .ZN(new_n789));
  INV_X1    g603(.A(new_n570), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n646), .A2(new_n706), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n612), .A2(new_n433), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n606), .A2(new_n792), .A3(new_n783), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT108), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n791), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n786), .A2(new_n789), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n709), .B1(new_n646), .B2(new_n697), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n797), .B(new_n695), .C1(new_n687), .C2(new_n689), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  AND4_X1   g613(.A1(new_n677), .A2(new_n723), .A3(new_n725), .A4(new_n727), .ZN(new_n800));
  AND4_X1   g614(.A1(new_n604), .A2(new_n703), .A3(new_n705), .A4(new_n636), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT109), .ZN(new_n802));
  INV_X1    g616(.A(new_n648), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n374), .A2(new_n380), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n802), .B1(new_n628), .B2(new_n805), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n627), .A2(new_n804), .A3(KEYINPUT109), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n726), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n808), .A2(new_n569), .A3(new_n636), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n800), .A2(new_n801), .B1(new_n646), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n810), .A2(new_n736), .A3(new_n739), .A4(new_n731), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n796), .A2(new_n799), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n678), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n713), .B1(new_n646), .B2(new_n814), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n708), .A2(new_n636), .A3(new_n648), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n672), .A2(new_n684), .A3(new_n721), .A4(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT100), .B1(new_n646), .B2(new_n651), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n334), .A2(new_n653), .A3(new_n650), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n815), .B(new_n817), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n801), .A2(new_n694), .A3(new_n616), .A4(new_n677), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n823), .B1(new_n334), .B2(new_n678), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n824), .B1(new_n652), .B2(new_n654), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT52), .B1(new_n825), .B2(new_n817), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n782), .B1(new_n813), .B2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n820), .A2(new_n821), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n825), .A2(KEYINPUT52), .A3(new_n817), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n798), .A2(new_n811), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n832), .A2(new_n833), .A3(KEYINPUT53), .A4(new_n796), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n828), .A2(new_n829), .A3(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n700), .A2(new_n726), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(new_n435), .A3(new_n762), .ZN(new_n837));
  AOI211_X1 g651(.A(new_n734), .B(new_n837), .C1(KEYINPUT120), .C2(KEYINPUT48), .ZN(new_n838));
  NOR2_X1   g652(.A1(KEYINPUT120), .A2(KEYINPUT48), .ZN(new_n839));
  XOR2_X1   g653(.A(new_n838), .B(new_n839), .Z(new_n840));
  NAND2_X1  g654(.A1(new_n762), .A2(new_n435), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n707), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n842), .A2(new_n616), .A3(new_n694), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(G952), .A3(new_n272), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n836), .A2(new_n706), .A3(new_n435), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n845), .A2(new_n672), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n844), .B1(new_n846), .B2(new_n792), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT119), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n840), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT51), .ZN(new_n850));
  OR3_X1    g664(.A1(new_n837), .A2(KEYINPUT116), .A3(new_n712), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT116), .B1(new_n837), .B2(new_n712), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n787), .B1(new_n607), .B2(new_n611), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n851), .A2(new_n852), .B1(new_n846), .B2(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n663), .A2(new_n694), .A3(new_n336), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n855), .A2(new_n856), .A3(new_n842), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n841), .A2(new_n707), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n663), .A2(new_n694), .A3(new_n336), .ZN(new_n859));
  OAI21_X1  g673(.A(KEYINPUT114), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT50), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n857), .A2(new_n860), .A3(KEYINPUT115), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n855), .A2(new_n842), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n862), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT50), .B1(new_n863), .B2(KEYINPUT114), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT115), .B1(new_n865), .B2(new_n857), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n854), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n771), .A2(new_n772), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n683), .A2(new_n518), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT118), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n842), .A2(new_n727), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n874), .B(KEYINPUT112), .Z(new_n875));
  NAND2_X1  g689(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n850), .B1(new_n869), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n871), .B(KEYINPUT113), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT51), .B1(new_n870), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n880), .B1(KEYINPUT117), .B2(new_n850), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n867), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n849), .B1(new_n877), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n834), .A2(KEYINPUT111), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n786), .A2(new_n789), .A3(new_n795), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n885), .A2(new_n798), .A3(new_n811), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT111), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n886), .A2(new_n887), .A3(KEYINPUT53), .A4(new_n832), .ZN(new_n888));
  AOI211_X1 g702(.A(KEYINPUT110), .B(KEYINPUT53), .C1(new_n886), .C2(new_n832), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT110), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n832), .A2(new_n796), .A3(new_n833), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n890), .B1(new_n891), .B2(new_n782), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n884), .B(new_n888), .C1(new_n889), .C2(new_n892), .ZN(new_n893));
  AOI211_X1 g707(.A(new_n835), .B(new_n883), .C1(new_n893), .C2(KEYINPUT54), .ZN(new_n894));
  NOR2_X1   g708(.A1(G952), .A2(G953), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n781), .B1(new_n894), .B2(new_n895), .ZN(G75));
  NOR2_X1   g710(.A1(new_n272), .A2(G952), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n289), .B1(new_n828), .B2(new_n834), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT56), .B1(new_n899), .B2(G210), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n512), .A2(new_n513), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n460), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n514), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT55), .Z(new_n904));
  OAI21_X1  g718(.A(new_n898), .B1(new_n900), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT56), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n899), .B2(new_n442), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n908), .A2(KEYINPUT121), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(KEYINPUT121), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n905), .B1(new_n909), .B2(new_n910), .ZN(G51));
  XOR2_X1   g725(.A(new_n741), .B(KEYINPUT57), .Z(new_n912));
  AOI21_X1  g726(.A(new_n829), .B1(new_n828), .B2(new_n834), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n912), .B1(new_n835), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n555), .ZN(new_n915));
  INV_X1    g729(.A(new_n899), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n916), .A2(new_n751), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n897), .B1(new_n915), .B2(new_n917), .ZN(G54));
  NAND2_X1  g732(.A1(KEYINPUT58), .A2(G475), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n916), .A2(new_n419), .A3(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n919), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n426), .B1(new_n899), .B2(new_n921), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n920), .A2(new_n897), .A3(new_n922), .ZN(G60));
  NAND2_X1  g737(.A1(new_n608), .A2(new_n610), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n372), .A2(new_n289), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT59), .Z(new_n926));
  OAI211_X1 g740(.A(new_n924), .B(new_n926), .C1(new_n835), .C2(new_n913), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n898), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n828), .A2(KEYINPUT110), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT53), .B1(new_n886), .B2(new_n832), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n890), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n884), .A2(new_n888), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n829), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n926), .B1(new_n934), .B2(new_n835), .ZN(new_n935));
  INV_X1    g749(.A(new_n924), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n928), .B1(new_n935), .B2(new_n936), .ZN(G63));
  NAND2_X1  g751(.A1(new_n828), .A2(new_n834), .ZN(new_n938));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT60), .Z(new_n940));
  NAND2_X1  g754(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n597), .B(KEYINPUT122), .Z(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n834), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n634), .B(new_n940), .C1(new_n944), .C2(new_n930), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n943), .A2(new_n898), .A3(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n943), .A2(KEYINPUT61), .A3(new_n898), .A4(new_n945), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(G66));
  INV_X1    g764(.A(G224), .ZN(new_n951));
  OAI21_X1  g765(.A(G953), .B1(new_n437), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n885), .A2(new_n798), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n952), .B1(new_n953), .B2(G953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n901), .B1(G898), .B2(new_n272), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(G69));
  INV_X1    g770(.A(new_n708), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n754), .A2(new_n706), .A3(new_n957), .A4(new_n733), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n773), .A2(new_n768), .A3(new_n958), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n959), .A2(new_n737), .A3(new_n739), .A4(new_n825), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(KEYINPUT125), .ZN(new_n961));
  AND4_X1   g775(.A1(new_n739), .A2(new_n773), .A3(new_n768), .A4(new_n958), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT125), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n962), .A2(new_n963), .A3(new_n737), .A4(new_n825), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n961), .A2(new_n272), .A3(new_n964), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n283), .B(new_n400), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n966), .B1(G900), .B2(G953), .ZN(new_n967));
  AOI21_X1  g781(.A(KEYINPUT124), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n272), .B1(G227), .B2(G900), .ZN(new_n969));
  OR3_X1    g783(.A1(new_n968), .A2(KEYINPUT126), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n825), .A2(new_n674), .ZN(new_n971));
  OR3_X1    g785(.A1(new_n971), .A2(KEYINPUT123), .A3(KEYINPUT62), .ZN(new_n972));
  OAI21_X1  g786(.A(KEYINPUT123), .B1(new_n971), .B2(KEYINPUT62), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n787), .A2(new_n382), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n727), .B1(new_n792), .B2(new_n975), .ZN(new_n976));
  NOR4_X1   g790(.A1(new_n334), .A2(new_n600), .A3(new_n658), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n773), .A2(new_n768), .ZN(new_n978));
  AOI211_X1 g792(.A(new_n977), .B(new_n978), .C1(new_n971), .C2(KEYINPUT62), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n974), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n272), .ZN(new_n981));
  AOI22_X1  g795(.A1(new_n981), .A2(new_n966), .B1(new_n965), .B2(new_n967), .ZN(new_n982));
  OAI21_X1  g796(.A(KEYINPUT126), .B1(new_n968), .B2(new_n969), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n970), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n982), .B1(new_n970), .B2(new_n983), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(G72));
  NAND3_X1  g800(.A1(new_n974), .A2(new_n953), .A3(new_n979), .ZN(new_n987));
  NAND2_X1  g801(.A1(G472), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT63), .Z(new_n989));
  NAND2_X1  g803(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n990), .A2(new_n276), .A3(new_n285), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n285), .A2(new_n276), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n961), .A2(new_n953), .A3(new_n964), .ZN(new_n993));
  INV_X1    g807(.A(new_n989), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n991), .A2(new_n898), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n994), .B1(new_n287), .B2(new_n668), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n893), .A2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT127), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n893), .A2(KEYINPUT127), .A3(new_n997), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n996), .B1(new_n1000), .B2(new_n1001), .ZN(G57));
endmodule


