//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n444, new_n445, new_n446, new_n451, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n562, new_n564, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n609, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1129;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  INV_X1    g017(.A(G2072), .ZN(new_n443));
  INV_X1    g018(.A(G2078), .ZN(new_n444));
  NOR2_X1   g019(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g020(.A1(new_n445), .A2(G2084), .A3(G2090), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g022(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g023(.A(G452), .Z(G391));
  AND2_X1   g024(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g027(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g029(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n455));
  XNOR2_X1  g030(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n455), .B(new_n456), .ZN(new_n457));
  NOR4_X1   g032(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g036(.A(G261), .ZN(G325));
  NAND2_X1  g037(.A1(new_n457), .A2(G2106), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT68), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n464), .B1(G567), .B2(new_n459), .ZN(G319));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n468), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT69), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n469), .A2(new_n481), .A3(G125), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n473), .B1(new_n483), .B2(G2105), .ZN(G160));
  NAND2_X1  g059(.A1(new_n469), .A2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n477), .A2(G2105), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n488), .A2(KEYINPUT70), .A3(G136), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n490));
  INV_X1    g065(.A(G136), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n471), .B2(new_n491), .ZN(new_n492));
  OR2_X1    g067(.A1(G100), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n487), .A2(new_n489), .A3(new_n492), .A4(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  NAND4_X1  g071(.A1(new_n474), .A2(new_n476), .A3(G138), .A4(new_n470), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(G126), .A2(G2105), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n470), .A2(G138), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(new_n498), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(new_n469), .ZN(new_n503));
  OR2_X1    g078(.A1(G102), .A2(G2105), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n504), .B(G2104), .C1(G114), .C2(new_n470), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n499), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT72), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n499), .A2(new_n503), .A3(new_n508), .A4(new_n505), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(G164));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT73), .A2(KEYINPUT5), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  AND3_X1   g097(.A1(new_n512), .A2(new_n514), .A3(G543), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n522), .A2(G88), .B1(G50), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n525), .A2(new_n511), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n524), .A2(new_n526), .ZN(G166));
  AND2_X1   g102(.A1(new_n522), .A2(G89), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n523), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n528), .A2(new_n533), .ZN(G168));
  NAND2_X1  g109(.A1(new_n523), .A2(G52), .ZN(new_n535));
  XNOR2_X1  g110(.A(KEYINPUT74), .B(G90), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n521), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n511), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n537), .A2(new_n539), .ZN(G171));
  NAND2_X1  g115(.A1(new_n523), .A2(G43), .ZN(new_n541));
  INV_X1    g116(.A(G81), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OAI221_X1 g118(.A(new_n541), .B1(new_n521), .B2(new_n542), .C1(new_n543), .C2(new_n511), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(G188));
  NAND2_X1  g127(.A1(new_n522), .A2(G91), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT76), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n520), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(new_n511), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n523), .A2(G53), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT9), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n554), .A2(new_n556), .A3(new_n558), .ZN(G299));
  INV_X1    g134(.A(G171), .ZN(G301));
  INV_X1    g135(.A(G168), .ZN(G286));
  INV_X1    g136(.A(KEYINPUT77), .ZN(new_n562));
  XNOR2_X1  g137(.A(G166), .B(new_n562), .ZN(G303));
  OAI21_X1  g138(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n564));
  INV_X1    g139(.A(G87), .ZN(new_n565));
  INV_X1    g140(.A(G49), .ZN(new_n566));
  INV_X1    g141(.A(new_n523), .ZN(new_n567));
  OAI221_X1 g142(.A(new_n564), .B1(new_n521), .B2(new_n565), .C1(new_n566), .C2(new_n567), .ZN(G288));
  NAND2_X1  g143(.A1(new_n523), .A2(G48), .ZN(new_n569));
  INV_X1    g144(.A(G86), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n521), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n520), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n511), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G305));
  NAND2_X1  g150(.A1(new_n523), .A2(G47), .ZN(new_n576));
  INV_X1    g151(.A(G85), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n521), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(new_n511), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G290));
  INV_X1    g157(.A(G868), .ZN(new_n583));
  OAI21_X1  g158(.A(KEYINPUT78), .B1(G171), .B2(new_n583), .ZN(new_n584));
  OR3_X1    g159(.A1(G171), .A2(KEYINPUT78), .A3(new_n583), .ZN(new_n585));
  INV_X1    g160(.A(G92), .ZN(new_n586));
  OAI21_X1  g161(.A(KEYINPUT79), .B1(new_n521), .B2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT79), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n515), .A2(new_n520), .A3(new_n588), .A4(G92), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n520), .A2(G66), .ZN(new_n593));
  INV_X1    g168(.A(G79), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n594), .B2(new_n517), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(G54), .B2(new_n523), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n587), .A2(KEYINPUT10), .A3(new_n589), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n592), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT80), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n592), .A2(KEYINPUT80), .A3(new_n596), .A4(new_n597), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n584), .B(new_n585), .C1(new_n603), .C2(G868), .ZN(G284));
  OAI211_X1 g179(.A(new_n584), .B(new_n585), .C1(new_n603), .C2(G868), .ZN(G321));
  NAND2_X1  g180(.A1(G299), .A2(new_n583), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n583), .B2(G168), .ZN(G297));
  OAI21_X1  g182(.A(new_n606), .B1(new_n583), .B2(G168), .ZN(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n603), .B1(new_n609), .B2(G860), .ZN(G148));
  NOR2_X1   g185(.A1(new_n546), .A2(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n603), .A2(new_n609), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(G868), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT81), .Z(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n469), .A2(new_n467), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2100), .ZN(new_n619));
  INV_X1    g194(.A(G135), .ZN(new_n620));
  OR3_X1    g195(.A1(new_n471), .A2(KEYINPUT82), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(KEYINPUT82), .B1(new_n471), .B2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n486), .A2(G123), .ZN(new_n623));
  OR2_X1    g198(.A1(G99), .A2(G2105), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n624), .B(G2104), .C1(G111), .C2(new_n470), .ZN(new_n625));
  NAND4_X1  g200(.A1(new_n621), .A2(new_n622), .A3(new_n623), .A4(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(G2096), .Z(new_n627));
  NAND2_X1  g202(.A1(new_n619), .A2(new_n627), .ZN(G156));
  XNOR2_X1  g203(.A(G2427), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT15), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2435), .Z(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(KEYINPUT14), .ZN(new_n633));
  XOR2_X1   g208(.A(G2443), .B(G2446), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(G1341), .B(G1348), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n635), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(G14), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n640), .A2(new_n641), .ZN(G401));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2067), .B(G2678), .Z(new_n645));
  NOR2_X1   g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n646), .B1(KEYINPUT83), .B2(KEYINPUT17), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n644), .A2(new_n645), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n647), .B(new_n648), .C1(KEYINPUT83), .C2(KEYINPUT17), .ZN(new_n649));
  INV_X1    g224(.A(KEYINPUT18), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g226(.A1(G2072), .A2(G2078), .ZN(new_n652));
  OAI22_X1  g227(.A1(new_n646), .A2(new_n650), .B1(new_n445), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n651), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2096), .B(G2100), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n654), .B(new_n655), .Z(G227));
  XOR2_X1   g231(.A(G1956), .B(G2474), .Z(new_n657));
  XOR2_X1   g232(.A(G1961), .B(G1966), .Z(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT85), .Z(new_n662));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n660), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT20), .Z(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(new_n659), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT84), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n665), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1991), .B(G1996), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G1981), .ZN(new_n674));
  INV_X1    g249(.A(G1986), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n672), .B(new_n676), .Z(G229));
  INV_X1    g252(.A(G16), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G6), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(new_n574), .B2(new_n678), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT32), .ZN(new_n681));
  INV_X1    g256(.A(G1981), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(G16), .A2(G22), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(G166), .B2(G16), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n685), .A2(G1971), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(G1971), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n678), .A2(G23), .ZN(new_n688));
  INV_X1    g263(.A(G288), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n688), .B1(new_n689), .B2(new_n678), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT33), .B(G1976), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT87), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n690), .B(new_n692), .ZN(new_n693));
  NAND4_X1  g268(.A1(new_n683), .A2(new_n686), .A3(new_n687), .A4(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT34), .Z(new_n695));
  NAND2_X1  g270(.A1(new_n678), .A2(G24), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(new_n581), .B2(new_n678), .ZN(new_n697));
  MUX2_X1   g272(.A(new_n696), .B(new_n697), .S(KEYINPUT86), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(new_n675), .ZN(new_n699));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G25), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n486), .A2(G119), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n488), .A2(G131), .ZN(new_n703));
  OR2_X1    g278(.A1(G95), .A2(G2105), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n704), .B(G2104), .C1(G107), .C2(new_n470), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n701), .B1(new_n707), .B2(new_n700), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT35), .B(G1991), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n695), .A2(new_n699), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT36), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n712), .A2(KEYINPUT88), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n711), .B(new_n713), .Z(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT31), .B(G11), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(G299), .A2(G16), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n678), .A2(KEYINPUT23), .A3(G20), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT23), .ZN(new_n719));
  INV_X1    g294(.A(G20), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(G16), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n717), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G1956), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  NOR2_X1   g300(.A1(G29), .A2(G35), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G162), .B2(G29), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT99), .B(KEYINPUT29), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G2090), .ZN(new_n731));
  OAI22_X1  g306(.A1(new_n724), .A2(new_n725), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n732), .A2(KEYINPUT100), .ZN(new_n733));
  OR2_X1    g308(.A1(G29), .A2(G33), .ZN(new_n734));
  NAND2_X1  g309(.A1(G115), .A2(G2104), .ZN(new_n735));
  INV_X1    g310(.A(G127), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n477), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G2105), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT93), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n488), .A2(G139), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT92), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT91), .B(KEYINPUT25), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n467), .A2(G103), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n740), .A2(new_n743), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT94), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n734), .B1(new_n748), .B2(new_n700), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G2072), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n443), .B(new_n734), .C1(new_n748), .C2(new_n700), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(G160), .A2(G29), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT24), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n700), .B1(new_n754), .B2(G34), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT95), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n754), .A2(G34), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n755), .A2(new_n756), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n753), .A2(G2084), .A3(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(G29), .A2(G32), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n486), .A2(G129), .B1(new_n488), .B2(G141), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n467), .A2(G105), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT96), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT26), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n762), .B1(new_n769), .B2(G29), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT27), .B(G1996), .Z(new_n771));
  OR2_X1    g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n752), .A2(new_n761), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(KEYINPUT97), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT97), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n752), .A2(new_n775), .A3(new_n761), .A4(new_n772), .ZN(new_n776));
  AOI211_X1 g351(.A(new_n716), .B(new_n733), .C1(new_n774), .C2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n700), .A2(G27), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G164), .B2(new_n700), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(new_n444), .ZN(new_n780));
  OAI21_X1  g355(.A(KEYINPUT98), .B1(G5), .B2(G16), .ZN(new_n781));
  OR3_X1    g356(.A1(KEYINPUT98), .A2(G5), .A3(G16), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n781), .B(new_n782), .C1(G301), .C2(new_n678), .ZN(new_n783));
  INV_X1    g358(.A(G1961), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n780), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n603), .A2(new_n678), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G4), .B2(new_n678), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT89), .B(G1348), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n777), .A2(new_n786), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n626), .A2(new_n700), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n732), .A2(KEYINPUT100), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT30), .B(G28), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n770), .A2(new_n771), .B1(new_n700), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n678), .A2(G19), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n546), .B2(new_n678), .ZN(new_n799));
  OAI221_X1 g374(.A(new_n797), .B1(G1341), .B2(new_n799), .C1(new_n729), .C2(G2090), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n753), .A2(new_n760), .ZN(new_n802));
  INV_X1    g377(.A(G2084), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n799), .A2(G1341), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT28), .ZN(new_n806));
  INV_X1    g381(.A(G26), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(G29), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n807), .A2(G29), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n486), .A2(G128), .B1(new_n488), .B2(G140), .ZN(new_n810));
  OAI21_X1  g385(.A(G2104), .B1(new_n470), .B2(G116), .ZN(new_n811));
  NOR2_X1   g386(.A1(G104), .A2(G2105), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT90), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n810), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n809), .B1(new_n814), .B2(G29), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n808), .B1(new_n815), .B2(new_n806), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(G2067), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(G2067), .ZN(new_n818));
  AND3_X1   g393(.A1(new_n805), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n801), .A2(new_n804), .A3(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(G168), .A2(G16), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G16), .B2(G21), .ZN(new_n823));
  INV_X1    g398(.A(G1966), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n825), .B(new_n826), .C1(new_n783), .C2(new_n784), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n794), .A2(new_n795), .A3(new_n821), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(KEYINPUT101), .ZN(new_n830));
  NOR4_X1   g405(.A1(new_n792), .A2(new_n820), .A3(new_n827), .A4(new_n793), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT101), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n831), .A2(new_n832), .A3(new_n795), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n714), .B1(new_n830), .B2(new_n833), .ZN(G311));
  INV_X1    g409(.A(new_n714), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n829), .A2(KEYINPUT101), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n832), .B1(new_n831), .B2(new_n795), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(G150));
  NAND2_X1  g413(.A1(new_n523), .A2(G55), .ZN(new_n839));
  INV_X1    g414(.A(G93), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n521), .B2(new_n840), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n842), .A2(new_n511), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(G860), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT37), .Z(new_n847));
  NOR2_X1   g422(.A1(new_n602), .A2(new_n609), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n546), .A2(new_n845), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n844), .A2(new_n544), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n848), .B(new_n851), .ZN(new_n852));
  XOR2_X1   g427(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n847), .B1(new_n854), .B2(G860), .ZN(G145));
  XNOR2_X1  g430(.A(new_n814), .B(new_n506), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n769), .ZN(new_n857));
  INV_X1    g432(.A(new_n748), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT103), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n747), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n861), .B1(new_n862), .B2(new_n857), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n488), .A2(G142), .ZN(new_n864));
  OAI21_X1  g439(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n470), .A2(G118), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(G130), .B2(new_n486), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(new_n617), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n706), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n863), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n863), .A2(new_n870), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(KEYINPUT104), .A3(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(G160), .B(KEYINPUT102), .Z(new_n874));
  XNOR2_X1  g449(.A(new_n626), .B(new_n495), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n873), .B(new_n876), .C1(KEYINPUT104), .C2(new_n872), .ZN(new_n877));
  INV_X1    g452(.A(G37), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n871), .A2(new_n872), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n877), .B(new_n878), .C1(new_n879), .C2(new_n876), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g456(.A1(new_n845), .A2(new_n583), .ZN(new_n882));
  XOR2_X1   g457(.A(G299), .B(new_n598), .Z(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(KEYINPUT41), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n612), .B(new_n851), .ZN(new_n885));
  MUX2_X1   g460(.A(new_n883), .B(new_n884), .S(new_n885), .Z(new_n886));
  XNOR2_X1  g461(.A(G166), .B(G288), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n574), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(G290), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT42), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n886), .B(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n882), .B1(new_n891), .B2(new_n583), .ZN(G295));
  OAI21_X1  g467(.A(new_n882), .B1(new_n891), .B2(new_n583), .ZN(G331));
  INV_X1    g468(.A(new_n851), .ZN(new_n894));
  XNOR2_X1  g469(.A(G168), .B(G171), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n884), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n897), .B(KEYINPUT105), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n896), .A2(new_n883), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n902), .A3(new_n889), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n889), .B1(new_n899), .B2(new_n902), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n904), .A2(new_n905), .A3(G37), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(KEYINPUT43), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n900), .A2(new_n896), .ZN(new_n908));
  AOI22_X1  g483(.A1(new_n908), .A2(new_n884), .B1(new_n897), .B2(new_n901), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n878), .B(new_n903), .C1(new_n909), .C2(new_n889), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n907), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n906), .A2(KEYINPUT43), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n910), .B(KEYINPUT106), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n915), .B1(new_n916), .B2(KEYINPUT43), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n914), .B1(new_n917), .B2(new_n913), .ZN(G397));
  INV_X1    g493(.A(new_n769), .ZN(new_n919));
  XNOR2_X1  g494(.A(KEYINPUT107), .B(G40), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(G160), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G1384), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n506), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT45), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n919), .A2(G1996), .A3(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT110), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n814), .B(G2067), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n927), .ZN(new_n931));
  OR3_X1    g506(.A1(new_n922), .A2(new_n926), .A3(G1996), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT109), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n929), .B(new_n931), .C1(new_n919), .C2(new_n933), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n707), .A2(new_n709), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n707), .A2(new_n709), .ZN(new_n936));
  AOI211_X1 g511(.A(new_n922), .B(new_n926), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n927), .A2(G1986), .A3(G290), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n927), .A2(new_n675), .A3(new_n581), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XOR2_X1   g515(.A(new_n940), .B(KEYINPUT108), .Z(new_n941));
  NOR3_X1   g516(.A1(new_n934), .A2(new_n937), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(G8), .ZN(new_n943));
  AOI211_X1 g518(.A(new_n920), .B(new_n473), .C1(G2105), .C2(new_n483), .ZN(new_n944));
  INV_X1    g519(.A(new_n924), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G1976), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n946), .B1(new_n947), .B2(G288), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n948), .A2(KEYINPUT52), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n949), .B1(G1976), .B2(new_n689), .ZN(new_n950));
  XNOR2_X1  g525(.A(KEYINPUT113), .B(G1981), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n574), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n952), .B1(new_n682), .B2(new_n574), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT49), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n946), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n948), .A2(KEYINPUT52), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n956), .A2(KEYINPUT112), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(KEYINPUT112), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n950), .B(new_n955), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT111), .ZN(new_n961));
  NAND2_X1  g536(.A1(G303), .A2(G8), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT55), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n963), .ZN(new_n965));
  NAND4_X1  g540(.A1(G303), .A2(KEYINPUT111), .A3(KEYINPUT55), .A4(G8), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n507), .A2(new_n923), .A3(new_n509), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n925), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n506), .A2(KEYINPUT45), .A3(new_n923), .ZN(new_n970));
  AND2_X1   g545(.A1(G160), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(new_n971), .A3(new_n921), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n973), .A2(G1971), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n922), .B1(KEYINPUT50), .B2(new_n968), .ZN(new_n976));
  OR2_X1    g551(.A1(new_n924), .A2(KEYINPUT50), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(new_n731), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n943), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n967), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n924), .A2(KEYINPUT50), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n944), .B(new_n981), .C1(new_n968), .C2(KEYINPUT50), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(G2090), .ZN(new_n983));
  OAI21_X1  g558(.A(G8), .B1(new_n974), .B2(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n984), .A2(new_n964), .A3(new_n965), .A4(new_n966), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n960), .A2(new_n980), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n923), .A4(new_n509), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(KEYINPUT114), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n926), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n944), .B1(new_n988), .B2(KEYINPUT114), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n824), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT115), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n976), .A2(new_n803), .A3(new_n977), .ZN(new_n995));
  OAI211_X1 g570(.A(KEYINPUT115), .B(new_n824), .C1(new_n990), .C2(new_n991), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n994), .A2(G168), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n997), .A2(KEYINPUT123), .A3(G8), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT123), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT122), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n997), .A2(new_n1002), .A3(G8), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1000), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(new_n1001), .A3(KEYINPUT51), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1006), .A2(G8), .A3(G286), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT62), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(new_n972), .B2(G2078), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT124), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n990), .A2(new_n991), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1010), .A2(G2078), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT124), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1016), .B(new_n1010), .C1(new_n972), .C2(G2078), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n976), .A2(new_n977), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n784), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1012), .A2(new_n1015), .A3(new_n1017), .A4(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(G171), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1003), .A2(new_n1001), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1023), .A2(new_n999), .A3(new_n998), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT62), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1024), .A2(new_n1025), .A3(new_n1007), .A4(new_n1005), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1009), .A2(new_n1022), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n1028));
  NAND2_X1  g603(.A1(G299), .A2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n554), .A2(KEYINPUT57), .A3(new_n556), .A4(new_n558), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g606(.A(KEYINPUT56), .B(G2072), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1032), .B(KEYINPUT117), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n973), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n982), .A2(new_n723), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1031), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1031), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G1348), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1018), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G2067), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n945), .A2(G160), .A3(new_n1043), .A4(new_n921), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1044), .B(KEYINPUT118), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n602), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1036), .B1(new_n1040), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1042), .A2(KEYINPUT60), .A3(new_n1045), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT120), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n603), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n602), .A2(KEYINPUT120), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1048), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n602), .A2(KEYINPUT120), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1053), .A2(new_n1042), .A3(KEYINPUT60), .A4(new_n1045), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT60), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1052), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT121), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1052), .A2(KEYINPUT121), .A3(new_n1054), .A4(new_n1057), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1039), .A2(new_n1036), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT61), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OR3_X1    g640(.A1(new_n972), .A2(KEYINPUT119), .A3(G1996), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT119), .B1(new_n972), .B2(G1996), .ZN(new_n1067));
  XOR2_X1   g642(.A(KEYINPUT58), .B(G1341), .Z(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n922), .B2(new_n924), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1066), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n546), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1039), .A2(KEYINPUT61), .A3(new_n1036), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1070), .A2(KEYINPUT59), .A3(new_n546), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1065), .A2(new_n1073), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1047), .B1(new_n1062), .B2(new_n1076), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1011), .A2(KEYINPUT124), .B1(new_n784), .B2(new_n1018), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n971), .A2(G40), .A3(new_n1014), .A4(new_n926), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1078), .A2(G301), .A3(new_n1017), .A4(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1021), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT125), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT125), .ZN(new_n1084));
  AOI211_X1 g659(.A(new_n1084), .B(KEYINPUT54), .C1(new_n1021), .C2(new_n1080), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1024), .A2(new_n1007), .A3(new_n1005), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1078), .A2(new_n1017), .A3(new_n1079), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1082), .B1(new_n1088), .B2(G171), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(G171), .B2(new_n1020), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1077), .A2(new_n1086), .A3(new_n1087), .A4(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n987), .B1(new_n1027), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n955), .A2(new_n947), .A3(new_n689), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n952), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(new_n946), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1006), .A2(G8), .A3(G168), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT63), .B1(new_n986), .B2(new_n1096), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n967), .A2(KEYINPUT116), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1096), .B1(new_n1098), .B2(new_n979), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n979), .B1(new_n967), .B2(KEYINPUT116), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1100), .A2(new_n960), .A3(KEYINPUT63), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  OAI221_X1 g677(.A(new_n1095), .B1(new_n980), .B2(new_n959), .C1(new_n1097), .C2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n942), .B1(new_n1092), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT126), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT126), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1106), .B(new_n942), .C1(new_n1092), .C2(new_n1103), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n927), .B1(new_n930), .B2(new_n919), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n933), .A2(KEYINPUT46), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n933), .A2(KEYINPUT46), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1112), .B(KEYINPUT47), .ZN(new_n1113));
  OAI22_X1  g688(.A1(new_n934), .A2(new_n936), .B1(G2067), .B2(new_n814), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n927), .ZN(new_n1115));
  XOR2_X1   g690(.A(new_n939), .B(KEYINPUT48), .Z(new_n1116));
  OR3_X1    g691(.A1(new_n934), .A2(new_n937), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1113), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  XOR2_X1   g693(.A(new_n1118), .B(KEYINPUT127), .Z(new_n1119));
  NAND2_X1  g694(.A1(new_n1108), .A2(new_n1119), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g695(.A(G401), .ZN(new_n1122));
  INV_X1    g696(.A(G227), .ZN(new_n1123));
  NAND3_X1  g697(.A1(new_n880), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  AND3_X1   g698(.A1(new_n907), .A2(new_n912), .A3(G319), .ZN(new_n1125));
  INV_X1    g699(.A(G229), .ZN(new_n1126));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g701(.A1(new_n1124), .A2(new_n1127), .ZN(G308));
  AND2_X1   g702(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1129));
  NAND4_X1  g703(.A1(new_n1129), .A2(new_n1122), .A3(new_n1123), .A4(new_n880), .ZN(G225));
endmodule


