//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934;
  XOR2_X1   g000(.A(G113gat), .B(G141gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT11), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT97), .ZN(new_n204));
  XNOR2_X1  g003(.A(G169gat), .B(G197gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209));
  XOR2_X1   g008(.A(G43gat), .B(G50gat), .Z(new_n210));
  OR3_X1    g009(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT98), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n211), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n215), .B1(new_n214), .B2(new_n211), .ZN(new_n216));
  INV_X1    g015(.A(G29gat), .ZN(new_n217));
  INV_X1    g016(.A(G36gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  AOI211_X1 g019(.A(new_n209), .B(new_n210), .C1(new_n216), .C2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT99), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n210), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n223), .B(new_n209), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n211), .B1(new_n213), .B2(KEYINPUT100), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(KEYINPUT100), .B2(new_n211), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n226), .A3(new_n220), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT101), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n224), .A2(KEYINPUT101), .A3(new_n226), .A4(new_n220), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n221), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT16), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n232), .A2(G1gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(G15gat), .B(G22gat), .ZN(new_n234));
  MUX2_X1   g033(.A(G1gat), .B(new_n233), .S(new_n234), .Z(new_n235));
  XNOR2_X1  g034(.A(new_n235), .B(G8gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(new_n231), .B(KEYINPUT17), .Z(new_n238));
  AOI21_X1  g037(.A(new_n237), .B1(new_n238), .B2(new_n236), .ZN(new_n239));
  NAND2_X1  g038(.A1(G229gat), .A2(G233gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(KEYINPUT18), .A3(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n231), .B(new_n236), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n240), .B(KEYINPUT13), .Z(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT18), .B1(new_n239), .B2(new_n240), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n208), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n239), .A2(new_n240), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT18), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n250), .A2(new_n241), .A3(new_n244), .A4(new_n207), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n255));
  NAND2_X1  g054(.A1(G183gat), .A2(G190gat), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT24), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(G183gat), .A2(G190gat), .ZN(new_n260));
  NOR3_X1   g059(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G169gat), .ZN(new_n262));
  INV_X1    g061(.A(G176gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT23), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT23), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n265), .B1(G169gat), .B2(G176gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(G169gat), .A2(G176gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n264), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n255), .B1(new_n261), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT65), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n256), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT66), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT66), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT24), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n271), .A2(new_n272), .A3(new_n273), .A4(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT67), .ZN(new_n277));
  INV_X1    g076(.A(new_n256), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n260), .B1(new_n278), .B2(KEYINPUT24), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n276), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT25), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n268), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n277), .B1(new_n276), .B2(new_n279), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n254), .B(new_n269), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n276), .A2(new_n279), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT67), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(new_n280), .A3(new_n282), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n254), .B1(new_n289), .B2(new_n269), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT27), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(G183gat), .ZN(new_n292));
  INV_X1    g091(.A(G183gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n293), .A2(KEYINPUT27), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT70), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G190gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n293), .A2(KEYINPUT27), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n291), .A2(G183gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT70), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n295), .A2(new_n296), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT28), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT28), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT69), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT27), .B(G183gat), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n304), .B1(new_n305), .B2(new_n296), .ZN(new_n306));
  AND4_X1   g105(.A1(new_n304), .A2(new_n297), .A3(new_n298), .A4(new_n296), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n303), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT71), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n302), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT72), .ZN(new_n311));
  OR2_X1    g110(.A1(new_n311), .A2(KEYINPUT26), .ZN(new_n312));
  INV_X1    g111(.A(new_n267), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n311), .B1(new_n313), .B2(KEYINPUT26), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n278), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n310), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n309), .B1(new_n302), .B2(new_n308), .ZN(new_n317));
  OAI22_X1  g116(.A1(new_n286), .A2(new_n290), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT74), .ZN(new_n319));
  INV_X1    g118(.A(G120gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(KEYINPUT74), .A2(G120gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(G113gat), .A3(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n320), .A2(G113gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT75), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT75), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n323), .A2(new_n328), .A3(new_n325), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(G127gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(G134gat), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT1), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G134gat), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n334), .B1(G127gat), .B2(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(KEYINPUT73), .B(G134gat), .Z(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(G127gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(new_n332), .ZN(new_n339));
  INV_X1    g138(.A(G113gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n340), .A2(G120gat), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n333), .B1(new_n324), .B2(new_n341), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n330), .A2(new_n336), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n318), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(G227gat), .ZN(new_n345));
  INV_X1    g144(.A(G233gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n317), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(new_n310), .A3(new_n315), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n269), .B1(new_n283), .B2(new_n284), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT68), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n285), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n323), .A2(new_n328), .A3(new_n325), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n328), .B1(new_n323), .B2(new_n325), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n336), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n342), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n349), .A2(new_n352), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n344), .A2(new_n347), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT33), .ZN(new_n360));
  XOR2_X1   g159(.A(G15gat), .B(G43gat), .Z(new_n361));
  XNOR2_X1  g160(.A(G71gat), .B(G99gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n359), .B(KEYINPUT32), .C1(new_n360), .C2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n364), .B1(new_n359), .B2(KEYINPUT32), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n359), .A2(new_n360), .ZN(new_n367));
  AND3_X1   g166(.A1(new_n366), .A2(KEYINPUT76), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT76), .B1(new_n366), .B2(new_n367), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n365), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n344), .A2(new_n358), .ZN(new_n371));
  INV_X1    g170(.A(new_n347), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  XOR2_X1   g172(.A(KEYINPUT77), .B(KEYINPUT34), .Z(new_n374));
  XOR2_X1   g173(.A(new_n373), .B(new_n374), .Z(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n370), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n375), .B(new_n365), .C1(new_n369), .C2(new_n368), .ZN(new_n378));
  INV_X1    g177(.A(G22gat), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT3), .ZN(new_n380));
  XOR2_X1   g179(.A(G197gat), .B(G204gat), .Z(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT78), .B(G211gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G218gat), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT22), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n381), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n385), .A2(KEYINPUT79), .ZN(new_n386));
  XNOR2_X1  g185(.A(G211gat), .B(G218gat), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(new_n385), .B2(KEYINPUT79), .ZN(new_n388));
  OR2_X1    g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n388), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n380), .B1(new_n391), .B2(KEYINPUT29), .ZN(new_n392));
  INV_X1    g191(.A(G155gat), .ZN(new_n393));
  INV_X1    g192(.A(G162gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(G155gat), .A2(G162gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT82), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n395), .A2(KEYINPUT82), .A3(new_n396), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  XOR2_X1   g200(.A(G141gat), .B(G148gat), .Z(new_n402));
  NAND2_X1  g201(.A1(new_n396), .A2(KEYINPUT2), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT83), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n396), .A2(KEYINPUT83), .A3(KEYINPUT2), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n402), .A2(new_n407), .A3(new_n397), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n392), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT29), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n402), .A2(new_n397), .A3(new_n407), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n413), .A2(new_n408), .B1(new_n401), .B2(new_n404), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n380), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n389), .A2(new_n390), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(G228gat), .A2(G233gat), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n419), .B1(new_n416), .B2(KEYINPUT88), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n411), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n420), .B1(new_n411), .B2(new_n417), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n379), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n385), .A2(KEYINPUT79), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n388), .B(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT3), .B1(new_n425), .B2(new_n412), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n417), .B1(new_n426), .B2(new_n414), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n427), .B(new_n419), .C1(KEYINPUT88), .C2(new_n416), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n417), .A3(new_n420), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(G22gat), .A3(new_n429), .ZN(new_n430));
  XOR2_X1   g229(.A(G78gat), .B(G106gat), .Z(new_n431));
  XNOR2_X1  g230(.A(KEYINPUT31), .B(G50gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT89), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n423), .A2(new_n430), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n435), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n428), .A2(G22gat), .A3(new_n429), .A4(new_n437), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n379), .B(new_n433), .C1(new_n421), .C2(new_n422), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n377), .A2(new_n378), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT95), .ZN(new_n442));
  AND2_X1   g241(.A1(G226gat), .A2(G233gat), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n349), .A2(new_n352), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n350), .B1(new_n316), .B2(new_n317), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n443), .A2(KEYINPUT29), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n391), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n350), .B(new_n443), .C1(new_n316), .C2(new_n317), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n310), .A2(new_n315), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n451), .A2(new_n348), .B1(new_n351), .B2(new_n285), .ZN(new_n452));
  INV_X1    g251(.A(new_n446), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n391), .B(new_n450), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(G8gat), .B(G36gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(G64gat), .B(G92gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n455), .B(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n449), .A2(KEYINPUT30), .A3(new_n454), .A4(new_n458), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n452), .A2(new_n443), .B1(new_n446), .B2(new_n445), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n454), .B1(new_n460), .B2(new_n391), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n457), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n463), .B(KEYINPUT80), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n414), .A2(new_n356), .A3(new_n355), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT4), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT86), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n357), .A2(KEYINPUT4), .A3(new_n410), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT85), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT85), .B1(new_n465), .B2(KEYINPUT4), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT86), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n465), .A2(new_n472), .A3(KEYINPUT4), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n467), .A2(new_n470), .A3(new_n471), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n410), .A2(KEYINPUT3), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n415), .A2(new_n475), .A3(new_n357), .ZN(new_n476));
  NAND2_X1  g275(.A1(G225gat), .A2(G233gat), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n478), .A2(KEYINPUT5), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n474), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT4), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n481), .B1(new_n343), .B2(new_n414), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n477), .B(new_n476), .C1(new_n482), .C2(new_n468), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT5), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n357), .A2(new_n410), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n465), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n484), .B1(new_n486), .B2(new_n478), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n483), .A2(KEYINPUT84), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT84), .B1(new_n483), .B2(new_n487), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n480), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G1gat), .B(G29gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(KEYINPUT0), .ZN(new_n492));
  XNOR2_X1  g291(.A(G57gat), .B(G85gat), .ZN(new_n493));
  XOR2_X1   g292(.A(new_n492), .B(new_n493), .Z(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(KEYINPUT87), .B(KEYINPUT6), .Z(new_n497));
  OAI211_X1 g296(.A(new_n480), .B(new_n494), .C1(new_n488), .C2(new_n489), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n497), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n490), .A2(new_n495), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  OR3_X1    g301(.A1(new_n461), .A2(KEYINPUT81), .A3(new_n457), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT30), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT81), .B1(new_n461), .B2(new_n457), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n464), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT95), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n377), .A2(new_n440), .A3(new_n378), .A4(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n442), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n377), .A2(KEYINPUT94), .A3(new_n378), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT94), .B1(new_n377), .B2(new_n378), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT35), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n506), .A2(new_n463), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT92), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT92), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n490), .A2(new_n518), .A3(new_n495), .A4(new_n500), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n499), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  AND4_X1   g319(.A1(new_n515), .A2(new_n516), .A3(new_n440), .A4(new_n520), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n511), .A2(KEYINPUT35), .B1(new_n514), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n377), .A2(new_n378), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT36), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n377), .A2(new_n525), .A3(new_n378), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT38), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n458), .B1(new_n461), .B2(KEYINPUT37), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT93), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT37), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n454), .B(new_n532), .C1(new_n460), .C2(new_n391), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n534), .B1(new_n529), .B2(new_n530), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n528), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n425), .B(new_n450), .C1(new_n452), .C2(new_n453), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n537), .B(KEYINPUT37), .C1(new_n460), .C2(new_n425), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n458), .A2(KEYINPUT38), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n533), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT91), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT91), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n533), .A2(new_n538), .A3(new_n542), .A4(new_n539), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n541), .A2(new_n505), .A3(new_n503), .A4(new_n543), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n536), .A2(new_n520), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT40), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n477), .B1(new_n474), .B2(new_n476), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT90), .B(KEYINPUT39), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT39), .B1(new_n486), .B2(new_n478), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n494), .B1(new_n547), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n546), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  OR2_X1    g353(.A1(new_n547), .A2(new_n552), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n555), .A2(KEYINPUT40), .A3(new_n494), .A4(new_n550), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n554), .A2(new_n556), .A3(new_n496), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n516), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n440), .B1(new_n545), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n440), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n508), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n527), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n522), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT96), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT96), .B1(new_n522), .B2(new_n562), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n253), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G134gat), .B(G162gat), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n568), .B(new_n569), .Z(new_n570));
  NAND3_X1  g369(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(G99gat), .A2(G106gat), .ZN(new_n572));
  INV_X1    g371(.A(G85gat), .ZN(new_n573));
  INV_X1    g372(.A(G92gat), .ZN(new_n574));
  AOI22_X1  g373(.A1(KEYINPUT8), .A2(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT105), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G85gat), .A2(G92gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT7), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G99gat), .B(G106gat), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n580), .B(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT106), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n571), .B1(new_n584), .B2(new_n231), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT107), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n238), .A2(new_n584), .ZN(new_n587));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT108), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n570), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT109), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n589), .B1(new_n586), .B2(new_n587), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n594), .B1(new_n596), .B2(new_n590), .ZN(new_n597));
  INV_X1    g396(.A(new_n590), .ZN(new_n598));
  NOR3_X1   g397(.A1(new_n598), .A2(KEYINPUT109), .A3(new_n595), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n593), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(KEYINPUT109), .B1(new_n598), .B2(new_n595), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n596), .A2(new_n594), .A3(new_n590), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n601), .A2(new_n602), .A3(new_n592), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G183gat), .B(G211gat), .Z(new_n606));
  XNOR2_X1  g405(.A(G127gat), .B(G155gat), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n607), .B(KEYINPUT20), .Z(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT103), .ZN(new_n610));
  XOR2_X1   g409(.A(G57gat), .B(G64gat), .Z(new_n611));
  AND2_X1   g410(.A1(G71gat), .A2(G78gat), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n611), .B1(KEYINPUT9), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT102), .ZN(new_n614));
  XNOR2_X1  g413(.A(G71gat), .B(G78gat), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n616), .B1(new_n614), .B2(new_n615), .ZN(new_n617));
  INV_X1    g416(.A(new_n615), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT21), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n610), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n620), .A2(new_n610), .A3(new_n621), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n623), .A2(G231gat), .A3(G233gat), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G231gat), .A2(G233gat), .ZN(new_n626));
  INV_X1    g425(.A(new_n624), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n626), .B1(new_n627), .B2(new_n622), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT104), .B(KEYINPUT19), .Z(new_n629));
  NAND3_X1  g428(.A1(new_n625), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n629), .B1(new_n625), .B2(new_n628), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n609), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n625), .A2(new_n628), .ZN(new_n634));
  INV_X1    g433(.A(new_n629), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n636), .A2(new_n608), .A3(new_n630), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n236), .B1(new_n620), .B2(new_n621), .ZN(new_n638));
  AND3_X1   g437(.A1(new_n633), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n638), .B1(new_n633), .B2(new_n637), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n606), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n633), .A2(new_n637), .ZN(new_n642));
  INV_X1    g441(.A(new_n638), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n633), .A2(new_n637), .A3(new_n638), .ZN(new_n645));
  INV_X1    g444(.A(new_n606), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n583), .B(new_n620), .ZN(new_n649));
  NAND2_X1  g448(.A1(G230gat), .A2(G233gat), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n652), .B(KEYINPUT110), .Z(new_n653));
  OR2_X1    g452(.A1(new_n649), .A2(KEYINPUT10), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n617), .A2(KEYINPUT10), .A3(new_n619), .ZN(new_n655));
  OR2_X1    g454(.A1(new_n584), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(new_n650), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G120gat), .B(G148gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(G176gat), .B(G204gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n662), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n653), .A2(new_n664), .A3(new_n658), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n605), .A2(new_n648), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n567), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(new_n502), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n669), .B(G1gat), .Z(G1324gat));
  INV_X1    g469(.A(new_n516), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n567), .A2(new_n671), .A3(new_n667), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(G8gat), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(KEYINPUT42), .ZN(new_n674));
  NOR2_X1   g473(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n675));
  AND2_X1   g474(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n672), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  MUX2_X1   g476(.A(new_n674), .B(KEYINPUT42), .S(new_n677), .Z(G1325gat));
  INV_X1    g477(.A(new_n527), .ZN(new_n679));
  OAI21_X1  g478(.A(G15gat), .B1(new_n668), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n514), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n681), .A2(G15gat), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n680), .B1(new_n668), .B2(new_n682), .ZN(G1326gat));
  XNOR2_X1  g482(.A(KEYINPUT43), .B(G22gat), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT112), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n565), .A2(new_n566), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n687), .A2(new_n252), .A3(new_n560), .A4(new_n667), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT111), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT111), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n567), .A2(new_n690), .A3(new_n560), .A4(new_n667), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n686), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n689), .A2(new_n686), .A3(new_n691), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n685), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n694), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n696), .A2(new_n692), .A3(new_n684), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n695), .A2(new_n697), .ZN(G1327gat));
  NAND2_X1  g497(.A1(new_n687), .A2(new_n252), .ZN(new_n699));
  INV_X1    g498(.A(new_n666), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n605), .A2(new_n648), .A3(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n502), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n702), .A2(new_n217), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT45), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n605), .A2(KEYINPUT44), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n687), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n559), .A2(new_n561), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n679), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n511), .A2(KEYINPUT35), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n514), .A2(new_n521), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(KEYINPUT44), .B1(new_n713), .B2(new_n605), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n641), .A2(new_n647), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n253), .A2(new_n716), .A3(new_n666), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n708), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(G29gat), .B1(new_n718), .B2(new_n502), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n705), .A2(new_n719), .ZN(G1328gat));
  NAND3_X1  g519(.A1(new_n702), .A2(new_n218), .A3(new_n671), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT46), .Z(new_n722));
  OAI21_X1  g521(.A(G36gat), .B1(new_n718), .B2(new_n516), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(G1329gat));
  NOR3_X1   g523(.A1(new_n699), .A2(new_n681), .A3(new_n701), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n527), .A2(G43gat), .ZN(new_n726));
  OAI22_X1  g525(.A1(new_n725), .A2(G43gat), .B1(new_n718), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g527(.A1(new_n699), .A2(new_n440), .A3(new_n701), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n560), .A2(G50gat), .ZN(new_n730));
  OAI22_X1  g529(.A1(new_n729), .A2(G50gat), .B1(new_n718), .B2(new_n730), .ZN(new_n731));
  XOR2_X1   g530(.A(KEYINPUT113), .B(KEYINPUT48), .Z(new_n732));
  XOR2_X1   g531(.A(new_n731), .B(new_n732), .Z(G1331gat));
  AOI211_X1 g532(.A(new_n252), .B(new_n648), .C1(new_n603), .C2(new_n600), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n713), .A2(new_n666), .A3(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n703), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(G57gat), .ZN(G1332gat));
  INV_X1    g537(.A(KEYINPUT49), .ZN(new_n739));
  INV_X1    g538(.A(G64gat), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n736), .B(new_n671), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n740), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1333gat));
  OAI21_X1  g542(.A(G71gat), .B1(new_n735), .B2(new_n679), .ZN(new_n744));
  OR2_X1    g543(.A1(new_n681), .A2(G71gat), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n735), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g546(.A1(new_n736), .A2(new_n560), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(G78gat), .ZN(G1335gat));
  INV_X1    g548(.A(KEYINPUT114), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n648), .A2(new_n253), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(KEYINPUT114), .B1(new_n716), .B2(new_n252), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n713), .A2(KEYINPUT51), .A3(new_n605), .A4(new_n753), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n605), .B(new_n753), .C1(new_n522), .C2(new_n562), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT51), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n700), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(G85gat), .B1(new_n758), .B2(new_n703), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n706), .B1(new_n565), .B2(new_n566), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n753), .A2(new_n666), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n760), .A2(new_n714), .A3(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n502), .A2(new_n573), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n759), .B1(new_n762), .B2(new_n763), .ZN(G1336gat));
  AOI21_X1  g563(.A(G92gat), .B1(new_n758), .B2(new_n671), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n516), .A2(new_n574), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NOR4_X1   g566(.A1(new_n760), .A2(new_n714), .A3(new_n761), .A4(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(KEYINPUT115), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n755), .A2(new_n756), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n756), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n671), .B(new_n666), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n574), .ZN(new_n773));
  INV_X1    g572(.A(new_n761), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n708), .A2(new_n715), .A3(new_n774), .A4(new_n766), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT116), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  OAI211_X1 g575(.A(KEYINPUT52), .B(new_n769), .C1(new_n776), .C2(KEYINPUT115), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT115), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n765), .A2(new_n768), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n778), .B(new_n779), .C1(new_n780), .C2(KEYINPUT116), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n777), .A2(new_n781), .ZN(G1337gat));
  AOI21_X1  g581(.A(G99gat), .B1(new_n758), .B2(new_n514), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n527), .A2(G99gat), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n762), .B2(new_n784), .ZN(G1338gat));
  INV_X1    g584(.A(G106gat), .ZN(new_n786));
  INV_X1    g585(.A(new_n758), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n787), .B2(new_n440), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n762), .A2(G106gat), .A3(new_n560), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT117), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n790), .A2(KEYINPUT53), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(KEYINPUT53), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n792), .B(new_n793), .ZN(G1339gat));
  NOR2_X1   g593(.A1(new_n671), .A2(new_n502), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n654), .A2(new_n656), .A3(new_n651), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n658), .A2(KEYINPUT54), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n651), .B1(new_n654), .B2(new_n656), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n664), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n797), .A2(KEYINPUT55), .A3(new_n800), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n804), .A2(new_n665), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n252), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n239), .A2(new_n240), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n242), .A2(new_n243), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n206), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n666), .A2(new_n251), .A3(new_n809), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n601), .A2(new_n602), .A3(new_n592), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n592), .B1(new_n601), .B2(new_n602), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n806), .B(new_n810), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n805), .A2(new_n251), .A3(new_n809), .A4(new_n803), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n600), .A2(new_n814), .A3(new_n603), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n813), .A2(new_n648), .A3(new_n815), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n604), .A2(new_n253), .A3(new_n716), .A4(new_n700), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT118), .B1(new_n818), .B2(new_n440), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n820));
  AOI211_X1 g619(.A(new_n820), .B(new_n560), .C1(new_n816), .C2(new_n817), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n514), .B(new_n795), .C1(new_n819), .C2(new_n821), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n822), .A2(new_n340), .A3(new_n253), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n442), .A2(new_n510), .ZN(new_n824));
  INV_X1    g623(.A(new_n795), .ZN(new_n825));
  AOI211_X1 g624(.A(new_n824), .B(new_n825), .C1(new_n816), .C2(new_n817), .ZN(new_n826));
  AOI21_X1  g625(.A(G113gat), .B1(new_n826), .B2(new_n252), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n823), .A2(new_n827), .ZN(G1340gat));
  OAI21_X1  g627(.A(G120gat), .B1(new_n822), .B2(new_n700), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n826), .A2(new_n321), .A3(new_n322), .A4(new_n666), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(G1341gat));
  OAI21_X1  g630(.A(G127gat), .B1(new_n822), .B2(new_n648), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n826), .A2(new_n331), .A3(new_n716), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(G1342gat));
  AOI21_X1  g633(.A(new_n502), .B1(new_n816), .B2(new_n817), .ZN(new_n835));
  INV_X1    g634(.A(new_n824), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n604), .A2(new_n671), .ZN(new_n837));
  AND4_X1   g636(.A1(new_n337), .A2(new_n835), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n839), .A2(KEYINPUT56), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(KEYINPUT119), .ZN(new_n841));
  OAI21_X1  g640(.A(G134gat), .B1(new_n822), .B2(new_n604), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n839), .A2(KEYINPUT56), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(G1343gat));
  NOR2_X1   g643(.A1(new_n825), .A2(new_n527), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n560), .A2(KEYINPUT57), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT120), .ZN(new_n847));
  AOI22_X1  g646(.A1(new_n816), .A2(new_n847), .B1(new_n734), .B2(new_n700), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n813), .A2(KEYINPUT120), .A3(new_n648), .A4(new_n815), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n846), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n440), .B1(new_n816), .B2(new_n817), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n851), .A2(KEYINPUT57), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n252), .B(new_n845), .C1(new_n850), .C2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(G141gat), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n527), .A2(new_n440), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n253), .A2(G141gat), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n818), .A2(new_n795), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n854), .A2(new_n855), .A3(new_n858), .ZN(new_n859));
  XOR2_X1   g658(.A(new_n858), .B(KEYINPUT121), .Z(new_n860));
  NAND2_X1  g659(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT122), .B1(new_n861), .B2(KEYINPUT58), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT122), .ZN(new_n863));
  AOI211_X1 g662(.A(new_n863), .B(new_n855), .C1(new_n854), .C2(new_n860), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n859), .B1(new_n862), .B2(new_n864), .ZN(G1344gat));
  AND2_X1   g664(.A1(new_n835), .A2(new_n856), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n700), .A2(new_n671), .A3(G148gat), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n851), .B(KEYINPUT57), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n870), .A2(new_n666), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n845), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n869), .B1(new_n872), .B2(G148gat), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n869), .A2(G148gat), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n850), .A2(new_n852), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n875), .A2(new_n527), .A3(new_n825), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n874), .B1(new_n876), .B2(new_n666), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n868), .B1(new_n873), .B2(new_n877), .ZN(G1345gat));
  NOR2_X1   g677(.A1(new_n648), .A2(new_n393), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n818), .A2(new_n716), .A3(new_n795), .A4(new_n856), .ZN(new_n880));
  AOI22_X1  g679(.A1(new_n876), .A2(new_n879), .B1(new_n393), .B2(new_n880), .ZN(G1346gat));
  NAND3_X1  g680(.A1(new_n866), .A2(new_n394), .A3(new_n837), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT123), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n876), .A2(new_n605), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n883), .B1(new_n884), .B2(new_n394), .ZN(G1347gat));
  NOR2_X1   g684(.A1(new_n516), .A2(new_n703), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n514), .B(new_n886), .C1(new_n819), .C2(new_n821), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n887), .A2(new_n262), .A3(new_n253), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n836), .A2(new_n671), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT124), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n890), .A2(new_n502), .A3(new_n818), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(G169gat), .B1(new_n892), .B2(new_n252), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n888), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT125), .ZN(G1348gat));
  OAI21_X1  g694(.A(G176gat), .B1(new_n887), .B2(new_n700), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n892), .A2(new_n263), .A3(new_n666), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1349gat));
  NOR2_X1   g697(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n899));
  OAI21_X1  g698(.A(G183gat), .B1(new_n887), .B2(new_n648), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n892), .A2(new_n295), .A3(new_n300), .A4(new_n716), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AND2_X1   g701(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n902), .B(new_n903), .ZN(G1350gat));
  OAI21_X1  g703(.A(G190gat), .B1(new_n887), .B2(new_n604), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n905), .A2(KEYINPUT61), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT61), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n907), .B(G190gat), .C1(new_n887), .C2(new_n604), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n605), .A2(new_n296), .ZN(new_n910));
  OAI22_X1  g709(.A1(new_n906), .A2(new_n909), .B1(new_n891), .B2(new_n910), .ZN(G1351gat));
  NOR3_X1   g710(.A1(new_n527), .A2(new_n703), .A3(new_n516), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n851), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(G197gat), .B1(new_n914), .B2(new_n252), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n870), .A2(new_n912), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n252), .A2(G197gat), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(G1352gat));
  OR3_X1    g718(.A1(new_n913), .A2(G204gat), .A3(new_n700), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(KEYINPUT62), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT127), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n921), .B(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n871), .A2(new_n912), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G204gat), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n920), .A2(KEYINPUT62), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n923), .A2(new_n925), .A3(new_n926), .ZN(G1353gat));
  OR3_X1    g726(.A1(new_n913), .A2(new_n382), .A3(new_n648), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n870), .A2(new_n716), .A3(new_n912), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n929), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT63), .B1(new_n929), .B2(G211gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(G1354gat));
  OAI21_X1  g731(.A(G218gat), .B1(new_n916), .B2(new_n604), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n604), .A2(G218gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n933), .B1(new_n913), .B2(new_n934), .ZN(G1355gat));
endmodule


