//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n562, new_n563, new_n564,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n632, new_n633, new_n634, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1184,
    new_n1185;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n461), .A2(new_n463), .A3(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT67), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n466));
  NAND4_X1  g041(.A1(new_n461), .A2(new_n463), .A3(new_n466), .A4(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n475), .B1(new_n462), .B2(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n460), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n476), .A2(new_n477), .A3(new_n471), .A4(new_n463), .ZN(new_n478));
  INV_X1    g053(.A(G137), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n474), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n470), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  XOR2_X1   g058(.A(new_n478), .B(KEYINPUT69), .Z(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n476), .A2(new_n477), .A3(G2105), .A4(new_n463), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT70), .Z(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT71), .B1(G100), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NOR3_X1   g065(.A1(KEYINPUT71), .A2(G100), .A3(G2105), .ZN(new_n491));
  OAI221_X1 g066(.A(G2104), .B1(G112), .B2(new_n471), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n485), .A2(new_n488), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n476), .A2(new_n477), .A3(new_n496), .A4(new_n463), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n461), .A2(new_n463), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n495), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n497), .A2(KEYINPUT4), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G126), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n471), .A2(G114), .ZN(new_n502));
  OAI21_X1  g077(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n503));
  OAI22_X1  g078(.A1(new_n486), .A2(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n500), .A2(new_n504), .ZN(G164));
  OR2_X1    g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  AND2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n515), .A2(new_n516), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n511), .A2(new_n523), .ZN(G166));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  INV_X1    g101(.A(G89), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n527), .B2(new_n521), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT72), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n526), .B(KEYINPUT72), .C1(new_n527), .C2(new_n521), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n518), .A2(new_n517), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n510), .ZN(new_n533));
  INV_X1    g108(.A(G543), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n534), .B1(new_n512), .B2(new_n513), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n533), .A2(G63), .B1(G51), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n530), .A2(new_n531), .A3(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT73), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n530), .A2(KEYINPUT73), .A3(new_n531), .A4(new_n536), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(G168));
  AOI22_X1  g116(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n510), .ZN(new_n543));
  INV_X1    g118(.A(G52), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n515), .A2(new_n544), .B1(new_n521), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(G171));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n532), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G651), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(KEYINPUT74), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n506), .A2(new_n507), .B1(new_n512), .B2(new_n513), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n553), .A2(G81), .B1(new_n535), .B2(G43), .ZN(new_n554));
  AND2_X1   g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n551), .A2(KEYINPUT74), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT75), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(new_n564));
  XOR2_X1   g139(.A(new_n564), .B(KEYINPUT76), .Z(G188));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n515), .B2(new_n569), .ZN(new_n570));
  OAI211_X1 g145(.A(new_n535), .B(G53), .C1(new_n566), .C2(new_n567), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n570), .A2(new_n571), .B1(G91), .B2(new_n553), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n508), .A2(KEYINPUT78), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n532), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n574), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  AND2_X1   g153(.A1(G78), .A2(G543), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT79), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n582));
  OAI211_X1 g157(.A(new_n582), .B(G651), .C1(new_n578), .C2(new_n579), .ZN(new_n583));
  AOI211_X1 g158(.A(KEYINPUT80), .B(new_n573), .C1(new_n581), .C2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT80), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n581), .A2(new_n583), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n585), .B1(new_n586), .B2(new_n572), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(G299));
  INV_X1    g163(.A(G171), .ZN(G301));
  INV_X1    g164(.A(G168), .ZN(G286));
  INV_X1    g165(.A(G166), .ZN(G303));
  AOI22_X1  g166(.A1(new_n553), .A2(G87), .B1(new_n535), .B2(G49), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(KEYINPUT81), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT81), .ZN(new_n595));
  OAI211_X1 g170(.A(new_n595), .B(G651), .C1(new_n508), .C2(G74), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n592), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT82), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n598), .ZN(new_n600));
  AND2_X1   g175(.A1(new_n599), .A2(new_n600), .ZN(G288));
  OAI211_X1 g176(.A(G48), .B(G543), .C1(new_n519), .C2(new_n520), .ZN(new_n602));
  INV_X1    g177(.A(G86), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n521), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(G61), .B1(new_n518), .B2(new_n517), .ZN(new_n605));
  NAND2_X1  g180(.A1(G73), .A2(G543), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n510), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G305));
  AOI22_X1  g184(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n610), .A2(new_n510), .ZN(new_n611));
  INV_X1    g186(.A(G47), .ZN(new_n612));
  INV_X1    g187(.A(G85), .ZN(new_n613));
  OAI22_X1  g188(.A1(new_n515), .A2(new_n612), .B1(new_n521), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(G290));
  NAND2_X1  g191(.A1(G301), .A2(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n553), .A2(G92), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT10), .Z(new_n619));
  INV_X1    g194(.A(G66), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(new_n575), .B2(new_n577), .ZN(new_n621));
  NAND2_X1  g196(.A1(G79), .A2(G543), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT84), .Z(new_n623));
  OAI21_X1  g198(.A(G651), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(G54), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT83), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n625), .B1(new_n515), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(new_n626), .B2(new_n515), .ZN(new_n628));
  AND3_X1   g203(.A1(new_n619), .A2(new_n624), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n617), .B1(new_n629), .B2(G868), .ZN(G284));
  OAI21_X1  g205(.A(new_n617), .B1(new_n629), .B2(G868), .ZN(G321));
  NAND2_X1  g206(.A1(G286), .A2(G868), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT85), .ZN(new_n633));
  INV_X1    g208(.A(G299), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n633), .B1(G868), .B2(new_n634), .ZN(G297));
  OAI21_X1  g210(.A(new_n633), .B1(G868), .B2(new_n634), .ZN(G280));
  INV_X1    g211(.A(G559), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n629), .B1(new_n637), .B2(G860), .ZN(G148));
  INV_X1    g213(.A(G868), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n557), .A2(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(new_n629), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n641), .A2(G559), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n640), .B1(new_n642), .B2(new_n639), .ZN(G323));
  XNOR2_X1  g218(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g219(.A1(new_n487), .A2(G123), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n484), .A2(G135), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n471), .A2(G111), .ZN(new_n647));
  OAI21_X1  g222(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n645), .B(new_n646), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT89), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(G2096), .Z(new_n651));
  NAND2_X1  g226(.A1(new_n498), .A2(new_n473), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT87), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(KEYINPUT88), .B(G2100), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT13), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n655), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n651), .A2(new_n658), .ZN(G156));
  XOR2_X1   g234(.A(KEYINPUT15), .B(G2435), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2438), .ZN(new_n661));
  XOR2_X1   g236(.A(G2427), .B(G2430), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT90), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n663), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n664), .A2(KEYINPUT14), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2443), .B(G2446), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G1341), .B(G1348), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2451), .B(G2454), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT16), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT91), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n671), .A2(new_n674), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n675), .A2(G14), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT92), .Z(G401));
  INV_X1    g253(.A(KEYINPUT18), .ZN(new_n679));
  XOR2_X1   g254(.A(G2084), .B(G2090), .Z(new_n680));
  XNOR2_X1  g255(.A(G2067), .B(G2678), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(KEYINPUT17), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n680), .A2(new_n681), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n679), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G2100), .ZN(new_n686));
  XOR2_X1   g261(.A(G2072), .B(G2078), .Z(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(new_n682), .B2(KEYINPUT18), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G2096), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n686), .B(new_n689), .ZN(G227));
  XOR2_X1   g265(.A(G1971), .B(G1976), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT19), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1956), .B(G2474), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1961), .B(G1966), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  NOR3_X1   g271(.A1(new_n692), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n692), .A2(new_n695), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT20), .Z(new_n699));
  AOI211_X1 g274(.A(new_n697), .B(new_n699), .C1(new_n692), .C2(new_n696), .ZN(new_n700));
  INV_X1    g275(.A(G1981), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT93), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1991), .B(G1996), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n702), .B(new_n706), .Z(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT94), .B(G1986), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n702), .B(new_n706), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(new_n708), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n712), .ZN(G229));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(KEYINPUT95), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(KEYINPUT95), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n718), .A2(G19), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n558), .B2(new_n718), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(G1341), .Z(new_n721));
  NAND2_X1  g296(.A1(new_n714), .A2(G5), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G171), .B2(new_n714), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n723), .A2(G1961), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(G1961), .ZN(new_n725));
  INV_X1    g300(.A(G28), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n726), .A2(KEYINPUT30), .ZN(new_n727));
  AOI21_X1  g302(.A(G29), .B1(new_n726), .B2(KEYINPUT30), .ZN(new_n728));
  OR2_X1    g303(.A1(KEYINPUT31), .A2(G11), .ZN(new_n729));
  NAND2_X1  g304(.A1(KEYINPUT31), .A2(G11), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n727), .A2(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n725), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G2084), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT24), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n734), .A2(G34), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(G34), .ZN(new_n736));
  AOI21_X1  g311(.A(G29), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n482), .B2(G29), .ZN(new_n738));
  AOI211_X1 g313(.A(new_n724), .B(new_n732), .C1(new_n733), .C2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(G4), .A2(G16), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n629), .B2(G16), .ZN(new_n741));
  INV_X1    g316(.A(G1348), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n484), .A2(G139), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT25), .ZN(new_n745));
  NAND2_X1  g320(.A1(G103), .A2(G2104), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(G2105), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n471), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n498), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n744), .B(new_n749), .C1(new_n471), .C2(new_n750), .ZN(new_n751));
  MUX2_X1   g326(.A(G33), .B(new_n751), .S(G29), .Z(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G2072), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n721), .A2(new_n739), .A3(new_n743), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT27), .B(G1996), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT101), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n484), .A2(G141), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n487), .A2(G129), .ZN(new_n758));
  NAND3_X1  g333(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT99), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n760), .A2(KEYINPUT26), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(KEYINPUT26), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n761), .A2(new_n762), .B1(G105), .B2(new_n473), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n757), .A2(new_n758), .A3(new_n763), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT100), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G29), .ZN(new_n766));
  OR2_X1    g341(.A1(G29), .A2(G32), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n756), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(G27), .A2(G29), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G164), .B2(G29), .ZN(new_n770));
  INV_X1    g345(.A(G2078), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G29), .ZN(new_n773));
  OAI221_X1 g348(.A(new_n772), .B1(new_n733), .B2(new_n738), .C1(new_n650), .C2(new_n773), .ZN(new_n774));
  NOR3_X1   g349(.A1(new_n754), .A2(new_n768), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n717), .A2(G20), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT23), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n634), .B2(new_n714), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT102), .B(G1956), .Z(new_n779));
  NOR2_X1   g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n773), .A2(G35), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G162), .B2(new_n773), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT29), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n783), .A2(G2090), .ZN(new_n784));
  AND3_X1   g359(.A1(new_n766), .A2(new_n756), .A3(new_n767), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n780), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n752), .A2(G2072), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT98), .ZN(new_n788));
  NOR2_X1   g363(.A1(G16), .A2(G21), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G168), .B2(G16), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G1966), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n487), .A2(G128), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n484), .A2(G140), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n471), .A2(G116), .ZN(new_n794));
  OAI21_X1  g369(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n792), .B(new_n793), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n796), .A2(G29), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n773), .A2(G26), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT28), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G2067), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n788), .A2(new_n791), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n778), .A2(new_n779), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n783), .A2(G2090), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n775), .A2(new_n786), .A3(new_n802), .A4(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT103), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR4_X1   g384(.A1(new_n805), .A2(new_n754), .A3(new_n768), .A4(new_n774), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n810), .A2(KEYINPUT103), .A3(new_n786), .A4(new_n802), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT97), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n717), .A2(G22), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT96), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G303), .B2(new_n718), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G1971), .ZN(new_n818));
  MUX2_X1   g393(.A(G23), .B(new_n597), .S(G16), .Z(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT33), .B(G1976), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(G6), .A2(G16), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(new_n608), .B2(G16), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT32), .B(G1981), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n818), .A2(new_n821), .A3(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT34), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n487), .A2(G119), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n484), .A2(G131), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n471), .A2(G107), .ZN(new_n831));
  OAI21_X1  g406(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n829), .B(new_n830), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  MUX2_X1   g408(.A(G25), .B(new_n833), .S(G29), .Z(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT35), .B(G1991), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n718), .A2(G24), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(new_n615), .B2(new_n718), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(G1986), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n813), .B1(new_n828), .B2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n828), .A2(new_n840), .A3(new_n813), .ZN(new_n843));
  AOI21_X1  g418(.A(KEYINPUT36), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n843), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT36), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n845), .A2(new_n846), .A3(new_n841), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT104), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n812), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n849), .B1(new_n812), .B2(new_n848), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(G311));
  NAND2_X1  g427(.A1(new_n812), .A2(new_n848), .ZN(G150));
  AOI22_X1  g428(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n854), .A2(new_n510), .ZN(new_n855));
  INV_X1    g430(.A(G55), .ZN(new_n856));
  INV_X1    g431(.A(G93), .ZN(new_n857));
  OAI22_X1  g432(.A1(new_n515), .A2(new_n856), .B1(new_n521), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT105), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n858), .A2(new_n859), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n855), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(G860), .ZN(new_n863));
  XOR2_X1   g438(.A(KEYINPUT109), .B(KEYINPUT37), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT107), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n629), .A2(G559), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT106), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT38), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n557), .A2(new_n862), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n858), .B(new_n859), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n871), .A2(new_n555), .A3(new_n556), .A4(new_n855), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n869), .B(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n866), .B1(new_n874), .B2(KEYINPUT39), .ZN(new_n875));
  INV_X1    g450(.A(new_n873), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n869), .B(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n877), .A2(KEYINPUT107), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(G860), .B1(new_n874), .B2(KEYINPUT39), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n880), .A2(KEYINPUT108), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(KEYINPUT108), .B1(new_n880), .B2(new_n881), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n865), .B1(new_n882), .B2(new_n883), .ZN(G145));
  MUX2_X1   g459(.A(new_n765), .B(new_n764), .S(new_n751), .Z(new_n885));
  NOR2_X1   g460(.A1(new_n502), .A2(new_n503), .ZN(new_n886));
  AND4_X1   g461(.A1(G2105), .A2(new_n476), .A3(new_n463), .A4(new_n477), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n886), .B1(new_n887), .B2(G126), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n498), .A2(new_n499), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n796), .B(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n885), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n885), .A2(new_n894), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n833), .B(new_n655), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n484), .A2(G142), .ZN(new_n898));
  OR2_X1    g473(.A1(G106), .A2(G2105), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n899), .B(G2104), .C1(G118), .C2(new_n471), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n901), .B1(G130), .B2(new_n487), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n897), .B(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n895), .A2(new_n896), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT110), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n895), .A2(new_n896), .ZN(new_n906));
  INV_X1    g481(.A(new_n903), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT110), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n895), .A2(new_n896), .A3(new_n909), .A4(new_n903), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n650), .B(G160), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(new_n493), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n905), .A2(new_n908), .A3(new_n910), .A4(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(G37), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n908), .A2(new_n904), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n913), .B(new_n914), .C1(new_n915), .C2(new_n912), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g492(.A1(new_n586), .A2(new_n572), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT80), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n573), .B1(new_n581), .B2(new_n583), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n585), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(new_n921), .A3(new_n629), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n641), .B1(new_n584), .B2(new_n587), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT41), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n642), .B(new_n876), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT41), .B1(new_n922), .B2(new_n923), .ZN(new_n926));
  OR3_X1    g501(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n925), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n922), .A2(new_n923), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  XOR2_X1   g505(.A(new_n615), .B(new_n597), .Z(new_n931));
  OR2_X1    g506(.A1(new_n931), .A2(KEYINPUT111), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(KEYINPUT111), .ZN(new_n933));
  XNOR2_X1  g508(.A(G166), .B(new_n608), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n933), .A2(new_n934), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT42), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n930), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n639), .B1(new_n930), .B2(new_n938), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n939), .A2(new_n940), .A3(KEYINPUT112), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT112), .B1(new_n862), .B2(new_n639), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(G295));
  AOI21_X1  g519(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(G331));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT113), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n539), .A2(new_n540), .A3(G301), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(G301), .B1(new_n539), .B2(new_n540), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n873), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(G168), .A2(G171), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n952), .A2(new_n870), .A3(new_n872), .A4(new_n948), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n947), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n948), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT113), .B1(new_n955), .B2(new_n873), .ZN(new_n956));
  OAI22_X1  g531(.A1(new_n924), .A2(new_n926), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n937), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n929), .A2(new_n951), .A3(new_n953), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n960), .A2(new_n914), .ZN(new_n961));
  INV_X1    g536(.A(new_n954), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT115), .ZN(new_n963));
  INV_X1    g538(.A(new_n956), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n962), .A2(new_n963), .A3(new_n929), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n951), .A2(new_n953), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(new_n924), .B2(new_n926), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n954), .A2(new_n956), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n963), .B1(new_n969), .B2(new_n929), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n937), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n961), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT116), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n961), .A2(new_n971), .A3(KEYINPUT116), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n946), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n957), .A2(new_n959), .ZN(new_n977));
  OR2_X1    g552(.A1(new_n977), .A2(KEYINPUT114), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(KEYINPUT114), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(new_n937), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT43), .B1(new_n980), .B2(new_n961), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT44), .B1(new_n976), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n946), .B1(new_n980), .B2(new_n961), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n982), .A2(new_n986), .ZN(G397));
  INV_X1    g562(.A(G1384), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n988), .B1(new_n500), .B2(new_n504), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n470), .A2(new_n481), .A3(G40), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1996), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n765), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G2067), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n796), .B(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n764), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n995), .B(new_n997), .C1(new_n994), .C2(new_n998), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n999), .A2(new_n835), .A3(new_n833), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n796), .A2(G2067), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n993), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n993), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n1003), .A2(G1986), .A3(G290), .ZN(new_n1004));
  XOR2_X1   g579(.A(new_n1004), .B(KEYINPUT48), .Z(new_n1005));
  XNOR2_X1  g580(.A(new_n833), .B(new_n835), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n999), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1005), .B1(new_n1007), .B2(new_n1003), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1003), .B1(new_n997), .B2(new_n998), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n993), .A2(new_n994), .ZN(new_n1010));
  XOR2_X1   g585(.A(new_n1010), .B(KEYINPUT46), .Z(new_n1011));
  NOR2_X1   g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g587(.A(new_n1012), .B(KEYINPUT47), .Z(new_n1013));
  AND3_X1   g588(.A1(new_n1002), .A2(new_n1008), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT119), .B1(new_n608), .B2(new_n701), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT119), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1016), .B(G1981), .C1(new_n604), .C2(new_n607), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n605), .A2(new_n606), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(G651), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n553), .A2(G86), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1020), .A2(new_n1021), .A3(new_n701), .A4(new_n602), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT118), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT118), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n608), .A2(new_n1024), .A3(new_n701), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1018), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT49), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G8), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n464), .A2(KEYINPUT67), .B1(G113), .B2(G2104), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n471), .B1(new_n1031), .B2(new_n467), .ZN(new_n1032));
  INV_X1    g607(.A(G40), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n1032), .A2(new_n1033), .A3(new_n480), .ZN(new_n1034));
  INV_X1    g609(.A(new_n989), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1030), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1018), .A2(new_n1026), .A3(KEYINPUT49), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1029), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G1976), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n599), .A2(new_n1039), .A3(new_n600), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n1041));
  OR2_X1    g616(.A1(new_n597), .A2(new_n1039), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1040), .A2(new_n1036), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1036), .A2(new_n1042), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT52), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1038), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(G166), .A2(new_n1030), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1047), .B(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n989), .A2(KEYINPUT50), .ZN(new_n1050));
  INV_X1    g625(.A(G2090), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT50), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1052), .B(new_n988), .C1(new_n500), .C2(new_n504), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1050), .A2(new_n1034), .A3(new_n1051), .A4(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n1055));
  OAI211_X1 g630(.A(KEYINPUT45), .B(new_n988), .C1(new_n500), .C2(new_n504), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n991), .A2(new_n1034), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1971), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1054), .A2(new_n1055), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n992), .B1(KEYINPUT50), .B2(new_n989), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1060), .A2(KEYINPUT117), .A3(new_n1051), .A4(new_n1053), .ZN(new_n1061));
  AOI211_X1 g636(.A(new_n1030), .B(new_n1049), .C1(new_n1059), .C2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1046), .A2(new_n1062), .ZN(new_n1063));
  AOI211_X1 g638(.A(G1976), .B(G288), .C1(new_n1029), .C2(new_n1037), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1026), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1036), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(G286), .A2(G8), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT122), .ZN(new_n1069));
  INV_X1    g644(.A(G1966), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1057), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1050), .A2(new_n1034), .A3(new_n733), .A4(new_n1053), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1069), .B1(new_n1057), .B2(new_n1070), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT125), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n991), .A2(new_n1034), .A3(new_n1056), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT122), .B1(new_n1076), .B2(G1966), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT125), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1077), .A2(new_n1078), .A3(new_n1072), .A4(new_n1071), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1068), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1075), .A2(G168), .A3(new_n1079), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT51), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1082), .A2(new_n1030), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(G8), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1085), .A2(new_n1082), .A3(new_n1068), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1080), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1038), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1062), .A2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n991), .A2(new_n1034), .A3(new_n771), .A4(new_n1056), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1050), .A2(new_n1034), .A3(new_n1053), .ZN(new_n1092));
  INV_X1    g667(.A(G1961), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1090), .A2(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1094), .B1(new_n1091), .B2(new_n1090), .ZN(new_n1095));
  XNOR2_X1  g670(.A(G171), .B(KEYINPUT54), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT126), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1076), .A2(new_n1098), .A3(KEYINPUT53), .A4(new_n771), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1096), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1090), .A2(KEYINPUT126), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1094), .A2(new_n1099), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1097), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1052), .B1(new_n892), .B2(new_n988), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1104), .B1(new_n1105), .B2(new_n992), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1050), .A2(new_n1034), .A3(KEYINPUT120), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1106), .A2(new_n1051), .A3(new_n1053), .A4(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1108), .A2(KEYINPUT121), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT121), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n1110), .A2(new_n1111), .A3(new_n1030), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1049), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1089), .B(new_n1103), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1087), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT61), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1106), .A2(new_n1053), .A3(new_n1107), .ZN(new_n1117));
  INV_X1    g692(.A(G1956), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n920), .B(KEYINPUT57), .ZN(new_n1120));
  XNOR2_X1  g695(.A(KEYINPUT56), .B(G2072), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1076), .A2(new_n1121), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1119), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1120), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1116), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1120), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1119), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(KEYINPUT61), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT60), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1092), .A2(new_n742), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1034), .A2(new_n1035), .A3(new_n996), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n629), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n641), .A2(new_n1133), .A3(new_n1132), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1131), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT59), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n991), .A2(new_n1034), .A3(new_n994), .A4(new_n1056), .ZN(new_n1139));
  XOR2_X1   g714(.A(KEYINPUT58), .B(G1341), .Z(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(new_n992), .B2(new_n989), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1138), .B1(new_n1142), .B2(new_n558), .ZN(new_n1143));
  AOI211_X1 g718(.A(KEYINPUT59), .B(new_n557), .C1(new_n1139), .C2(new_n1141), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n629), .A2(new_n1131), .ZN(new_n1145));
  OAI22_X1  g720(.A1(new_n1143), .A2(new_n1144), .B1(new_n1134), .B2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1137), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1125), .A2(new_n1130), .A3(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1123), .A2(new_n1135), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1149), .A2(new_n1124), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1067), .B1(new_n1115), .B2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g727(.A(G8), .B(G168), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT63), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1062), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT123), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1061), .A2(new_n1157), .A3(new_n1109), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(G8), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(new_n1049), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1156), .B1(new_n1160), .B2(new_n1046), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1113), .B1(new_n1158), .B2(G8), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1162), .A2(new_n1088), .A3(KEYINPUT123), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1155), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1089), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1154), .B1(new_n1167), .B2(new_n1153), .ZN(new_n1168));
  OAI211_X1 g743(.A(KEYINPUT124), .B(new_n1155), .C1(new_n1161), .C2(new_n1163), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1166), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  AND3_X1   g745(.A1(new_n1152), .A2(KEYINPUT127), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(KEYINPUT127), .B1(new_n1152), .B2(new_n1170), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n1173));
  AND2_X1   g748(.A1(new_n1087), .A2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1087), .A2(new_n1173), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1094), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(G171), .ZN(new_n1177));
  NOR4_X1   g752(.A1(new_n1174), .A2(new_n1175), .A3(new_n1167), .A4(new_n1177), .ZN(new_n1178));
  NOR3_X1   g753(.A1(new_n1171), .A2(new_n1172), .A3(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n615), .B(G1986), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1003), .B1(new_n1007), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1014), .B1(new_n1179), .B2(new_n1181), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g757(.A1(G227), .A2(new_n458), .ZN(new_n1184));
  AND4_X1   g758(.A1(new_n677), .A2(new_n710), .A3(new_n712), .A4(new_n1184), .ZN(new_n1185));
  OAI211_X1 g759(.A(new_n916), .B(new_n1185), .C1(new_n984), .C2(new_n985), .ZN(G225));
  INV_X1    g760(.A(G225), .ZN(G308));
endmodule


