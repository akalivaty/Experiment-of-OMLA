//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1 1 0 1 0 1 1 0 0 0 0 0 0 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1338, new_n1339, new_n1340, new_n1341;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT0), .Z(new_n208));
  AOI22_X1  g0008(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT65), .Z(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n213));
  NAND3_X1  g0013(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n205), .B1(new_n210), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT1), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(KEYINPUT64), .ZN(new_n218));
  INV_X1    g0018(.A(KEYINPUT64), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n219), .A2(G1), .A3(G13), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  AOI211_X1 g0025(.A(new_n208), .B(new_n216), .C1(new_n223), .C2(new_n225), .ZN(G361));
  XOR2_X1   g0026(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n227));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G226), .B(G232), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n232), .B(new_n233), .Z(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n231), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT67), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  INV_X1    g0044(.A(KEYINPUT14), .ZN(new_n245));
  INV_X1    g0045(.A(G41), .ZN(new_n246));
  INV_X1    g0046(.A(G45), .ZN(new_n247));
  AOI21_X1  g0047(.A(G1), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G274), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g0051(.A(KEYINPUT68), .B1(G33), .B2(G41), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(new_n217), .ZN(new_n253));
  NAND3_X1  g0053(.A1(KEYINPUT68), .A2(G33), .A3(G41), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n249), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n251), .B1(new_n257), .B2(G238), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n221), .B1(G33), .B2(G41), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n264));
  AND3_X1   g0064(.A1(new_n262), .A2(new_n264), .A3(KEYINPUT69), .ZN(new_n265));
  AOI21_X1  g0065(.A(KEYINPUT69), .B1(new_n262), .B2(new_n264), .ZN(new_n266));
  OAI211_X1 g0066(.A(G226), .B(new_n260), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G97), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g0069(.A(G232), .B(G1698), .C1(new_n265), .C2(new_n266), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT74), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT69), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n261), .A2(G33), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n262), .A2(new_n264), .A3(KEYINPUT69), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n278), .A2(KEYINPUT74), .A3(G232), .A4(G1698), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n269), .B1(new_n272), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n259), .B1(new_n280), .B2(KEYINPUT75), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n272), .A2(new_n279), .ZN(new_n282));
  INV_X1    g0082(.A(new_n269), .ZN(new_n283));
  AND3_X1   g0083(.A1(new_n282), .A2(KEYINPUT75), .A3(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n258), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT13), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT13), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n287), .B(new_n258), .C1(new_n281), .C2(new_n284), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n245), .B1(new_n289), .B2(G169), .ZN(new_n290));
  INV_X1    g0090(.A(G169), .ZN(new_n291));
  AOI211_X1 g0091(.A(KEYINPUT14), .B(new_n291), .C1(new_n286), .C2(new_n288), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT78), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT77), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n286), .A2(new_n295), .A3(new_n288), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n282), .A2(new_n283), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT75), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n280), .A2(KEYINPUT75), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(new_n300), .A3(new_n259), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n301), .A2(KEYINPUT77), .A3(new_n287), .A4(new_n258), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n294), .B1(new_n303), .B2(G179), .ZN(new_n304));
  INV_X1    g0104(.A(G179), .ZN(new_n305));
  AOI211_X1 g0105(.A(KEYINPUT78), .B(new_n305), .C1(new_n296), .C2(new_n302), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n293), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n263), .A2(G20), .ZN(new_n308));
  INV_X1    g0108(.A(G68), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n308), .A2(G77), .B1(G20), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G50), .ZN(new_n311));
  NOR2_X1   g0111(.A1(G20), .A2(G33), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n310), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n205), .A2(new_n263), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n315), .B1(new_n218), .B2(new_n220), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  XOR2_X1   g0118(.A(new_n318), .B(KEYINPUT11), .Z(new_n319));
  INV_X1    g0119(.A(G13), .ZN(new_n320));
  NOR3_X1   g0120(.A1(new_n320), .A2(new_n222), .A3(G1), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n309), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT12), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n316), .B1(G1), .B2(new_n222), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n323), .B1(new_n309), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n319), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n307), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G200), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n286), .B2(new_n288), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n330), .B(KEYINPUT76), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n327), .B1(new_n303), .B2(G190), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n251), .ZN(new_n334));
  INV_X1    g0134(.A(G244), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n334), .B1(new_n256), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n278), .A2(G232), .A3(new_n260), .ZN(new_n337));
  INV_X1    g0137(.A(G107), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n278), .A2(G1698), .ZN(new_n339));
  INV_X1    g0139(.A(G238), .ZN(new_n340));
  OAI221_X1 g0140(.A(new_n337), .B1(new_n338), .B2(new_n278), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n336), .B1(new_n341), .B2(new_n259), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G190), .ZN(new_n343));
  XNOR2_X1  g0143(.A(KEYINPUT8), .B(G58), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n344), .A2(new_n313), .B1(new_n222), .B2(new_n202), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT71), .ZN(new_n346));
  XOR2_X1   g0146(.A(KEYINPUT15), .B(G87), .Z(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n308), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n345), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n346), .B2(new_n348), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n317), .ZN(new_n351));
  INV_X1    g0151(.A(new_n321), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(G77), .ZN(new_n353));
  INV_X1    g0153(.A(new_n324), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n353), .B1(new_n354), .B2(G77), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n343), .B(new_n357), .C1(new_n329), .C2(new_n342), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n342), .A2(new_n305), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n356), .B1(new_n342), .B2(G169), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(KEYINPUT72), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  OR2_X1    g0164(.A1(new_n361), .A2(new_n362), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT72), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n365), .A2(new_n366), .A3(new_n358), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g0168(.A(G58), .B(G68), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n369), .A2(G20), .B1(G159), .B2(new_n312), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n276), .A2(new_n222), .A3(new_n277), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT7), .ZN(new_n372));
  XNOR2_X1  g0172(.A(KEYINPUT79), .B(G33), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n264), .B1(new_n373), .B2(KEYINPUT3), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n372), .A2(G20), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n371), .A2(new_n372), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n370), .B1(new_n376), .B2(new_n309), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT16), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n274), .B1(new_n373), .B2(KEYINPUT3), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT7), .B1(new_n380), .B2(G20), .ZN(new_n381));
  AND2_X1   g0181(.A1(KEYINPUT79), .A2(G33), .ZN(new_n382));
  NOR2_X1   g0182(.A1(KEYINPUT79), .A2(G33), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT3), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n262), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n385), .A2(new_n372), .A3(new_n222), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n381), .A2(G68), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n387), .A2(KEYINPUT16), .A3(new_n370), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n379), .A2(new_n317), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(KEYINPUT70), .A2(G58), .ZN(new_n390));
  XNOR2_X1  g0190(.A(new_n390), .B(KEYINPUT8), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n352), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n354), .B2(new_n392), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n251), .B1(new_n257), .B2(G232), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n259), .ZN(new_n397));
  INV_X1    g0197(.A(G226), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(G1698), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n380), .B(new_n399), .C1(G223), .C2(G1698), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G33), .A2(G87), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n397), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(G169), .B1(new_n396), .B2(new_n402), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n400), .A2(new_n401), .ZN(new_n404));
  OAI211_X1 g0204(.A(G179), .B(new_n395), .C1(new_n404), .C2(new_n397), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n389), .A2(new_n394), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT18), .ZN(new_n407));
  OAI211_X1 g0207(.A(G190), .B(new_n395), .C1(new_n404), .C2(new_n397), .ZN(new_n408));
  OAI21_X1  g0208(.A(G200), .B1(new_n396), .B2(new_n402), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n389), .A2(new_n394), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n410), .B(KEYINPUT17), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n352), .A2(G50), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(new_n354), .B2(G50), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n391), .A2(new_n308), .ZN(new_n414));
  INV_X1    g0214(.A(G150), .ZN(new_n415));
  OAI22_X1  g0215(.A1(new_n415), .A2(new_n313), .B1(new_n201), .B2(new_n222), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n317), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n334), .B1(new_n256), .B2(new_n398), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n278), .A2(G222), .A3(new_n260), .ZN(new_n420));
  INV_X1    g0220(.A(G223), .ZN(new_n421));
  OAI221_X1 g0221(.A(new_n420), .B1(new_n202), .B2(new_n278), .C1(new_n339), .C2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n419), .B1(new_n422), .B2(new_n259), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n418), .B1(new_n423), .B2(G169), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n305), .B2(new_n423), .ZN(new_n425));
  INV_X1    g0225(.A(new_n423), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(G200), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT73), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n418), .A2(new_n428), .A3(KEYINPUT9), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n428), .A2(KEYINPUT9), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(KEYINPUT9), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n413), .A2(new_n430), .A3(new_n417), .A4(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n423), .A2(G190), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n427), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT10), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT10), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n427), .A2(new_n437), .A3(new_n433), .A4(new_n434), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n425), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n368), .A2(new_n407), .A3(new_n411), .A4(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n328), .A2(new_n333), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G1), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n321), .B1(new_n443), .B2(G33), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n316), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G107), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n321), .A2(new_n338), .ZN(new_n448));
  XOR2_X1   g0248(.A(new_n448), .B(KEYINPUT25), .Z(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT88), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n380), .A2(new_n452), .A3(new_n222), .A4(G87), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n384), .A2(new_n222), .A3(G87), .A4(new_n262), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT88), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(new_n455), .A3(KEYINPUT22), .ZN(new_n456));
  XOR2_X1   g0256(.A(KEYINPUT89), .B(KEYINPUT22), .Z(new_n457));
  NAND4_X1  g0257(.A1(new_n278), .A2(new_n222), .A3(G87), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n338), .A2(G20), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT23), .ZN(new_n461));
  OR2_X1    g0261(.A1(new_n460), .A2(KEYINPUT23), .ZN(new_n462));
  INV_X1    g0262(.A(new_n373), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G116), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n461), .B(new_n462), .C1(new_n464), .C2(G20), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT24), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n465), .B1(new_n456), .B2(new_n458), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n317), .B1(new_n470), .B2(KEYINPUT24), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n451), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n443), .A2(G45), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n246), .A2(KEYINPUT5), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT5), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G41), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n474), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  OR2_X1    g0278(.A1(new_n478), .A2(new_n250), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n255), .A2(new_n478), .ZN(new_n480));
  INV_X1    g0280(.A(G264), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n380), .A2(KEYINPUT90), .A3(G250), .A4(new_n260), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT90), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n260), .A2(G250), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n484), .B1(new_n385), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n380), .A2(G257), .A3(G1698), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n463), .A2(G294), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n483), .A2(new_n486), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  AOI211_X1 g0289(.A(G179), .B(new_n482), .C1(new_n489), .C2(new_n259), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n482), .B1(new_n489), .B2(new_n259), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n490), .B1(new_n291), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n472), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n265), .A2(new_n266), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G303), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT85), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n380), .A2(new_n497), .A3(G257), .A4(new_n260), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n384), .A2(G257), .A3(new_n260), .A4(new_n262), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT85), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n380), .A2(G264), .A3(G1698), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n496), .A2(new_n498), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n480), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n502), .A2(new_n259), .B1(G270), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n479), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G33), .A2(G283), .ZN(new_n507));
  INV_X1    g0307(.A(G97), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n507), .B(new_n222), .C1(G33), .C2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n222), .B2(G116), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(new_n316), .ZN(new_n511));
  OAI21_X1  g0311(.A(KEYINPUT86), .B1(new_n511), .B2(KEYINPUT20), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT86), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT20), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n513), .B(new_n514), .C1(new_n510), .C2(new_n316), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n511), .A2(KEYINPUT20), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n512), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n352), .A2(G116), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n518), .B1(new_n446), .B2(G116), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n506), .A2(G179), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n291), .B1(new_n517), .B2(new_n519), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n505), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT21), .B1(new_n523), .B2(KEYINPUT87), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT87), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT21), .ZN(new_n526));
  AOI211_X1 g0326(.A(new_n525), .B(new_n526), .C1(new_n505), .C2(new_n522), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n494), .B(new_n521), .C1(new_n524), .C2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n508), .A2(new_n338), .A3(KEYINPUT6), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT6), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G97), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n338), .A2(KEYINPUT80), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT80), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G107), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n529), .A2(new_n531), .A3(new_n532), .A4(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n529), .A2(new_n531), .B1(new_n532), .B2(new_n534), .ZN(new_n537));
  OAI21_X1  g0337(.A(G20), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT81), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n312), .A2(G77), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n529), .A2(new_n531), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n532), .A2(new_n534), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n222), .B1(new_n544), .B2(new_n535), .ZN(new_n545));
  INV_X1    g0345(.A(new_n540), .ZN(new_n546));
  OAI21_X1  g0346(.A(KEYINPUT81), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n541), .B(new_n547), .C1(new_n338), .C2(new_n376), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n317), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n352), .A2(G97), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n550), .B1(new_n446), .B2(G97), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT83), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n551), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n555), .B1(new_n548), .B2(new_n317), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(KEYINPUT83), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(G257), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n479), .B1(new_n480), .B2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n384), .A2(G244), .A3(new_n260), .A4(new_n262), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT4), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n562), .A2(new_n335), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n260), .B(new_n564), .C1(new_n265), .C2(new_n266), .ZN(new_n565));
  OAI211_X1 g0365(.A(G250), .B(G1698), .C1(new_n265), .C2(new_n266), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n563), .A2(new_n565), .A3(new_n566), .A4(new_n507), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n560), .B1(new_n567), .B2(new_n259), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G179), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n291), .B2(new_n568), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n558), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n473), .A2(G250), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n255), .A2(new_n573), .B1(G274), .B2(new_n474), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n340), .A2(G1698), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n384), .A2(new_n262), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT84), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n384), .A2(G244), .A3(G1698), .A4(new_n262), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT84), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n384), .A2(new_n580), .A3(new_n262), .A4(new_n576), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n578), .A2(new_n464), .A3(new_n579), .A4(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n575), .B1(new_n582), .B2(new_n259), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n305), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n380), .A2(new_n222), .A3(G68), .ZN(new_n585));
  AOI21_X1  g0385(.A(KEYINPUT19), .B1(new_n308), .B2(G97), .ZN(new_n586));
  INV_X1    g0386(.A(G87), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(new_n508), .A3(new_n338), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT19), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n222), .B1(new_n268), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n586), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n316), .B1(new_n585), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n352), .A2(new_n347), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n446), .A2(new_n347), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n584), .B(new_n596), .C1(G169), .C2(new_n583), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n582), .A2(new_n259), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n598), .A2(G190), .A3(new_n574), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n445), .A2(new_n587), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n592), .A2(new_n600), .A3(new_n593), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n599), .B(new_n601), .C1(new_n329), .C2(new_n583), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n471), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n470), .A2(KEYINPUT24), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n450), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(G190), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n492), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n491), .A2(new_n329), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n603), .B1(new_n606), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n520), .B1(new_n505), .B2(G200), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(new_n607), .B2(new_n505), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT82), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n568), .A2(G190), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n549), .A2(new_n615), .A3(new_n551), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n568), .A2(new_n329), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n614), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n617), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n619), .A2(KEYINPUT82), .A3(new_n556), .A4(new_n615), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n571), .A2(new_n611), .A3(new_n613), .A4(new_n621), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n442), .A2(new_n528), .A3(new_n622), .ZN(G372));
  AOI21_X1  g0423(.A(new_n363), .B1(new_n307), .B2(new_n327), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n333), .A2(new_n411), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n407), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n436), .A2(new_n438), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n425), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n597), .A2(new_n570), .A3(new_n552), .A4(new_n602), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n597), .B1(new_n629), .B2(KEYINPUT26), .ZN(new_n630));
  INV_X1    g0430(.A(new_n570), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n554), .B2(new_n557), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n597), .A2(new_n602), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n630), .B1(new_n634), .B2(KEYINPUT26), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n528), .A2(new_n571), .A3(new_n621), .A4(new_n611), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n628), .B1(new_n442), .B2(new_n638), .ZN(G369));
  OAI21_X1  g0439(.A(new_n521), .B1(new_n524), .B2(new_n527), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n320), .A2(G20), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n443), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(G213), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(G343), .ZN(new_n647));
  XOR2_X1   g0447(.A(new_n647), .B(KEYINPUT91), .Z(new_n648));
  AND2_X1   g0448(.A1(new_n648), .A2(new_n520), .ZN(new_n649));
  XNOR2_X1  g0449(.A(new_n640), .B(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n650), .A2(new_n613), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G330), .ZN(new_n652));
  INV_X1    g0452(.A(new_n648), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n606), .A2(new_n653), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n472), .A2(new_n608), .A3(new_n609), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n494), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n494), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n653), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n652), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n640), .A2(new_n653), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n658), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n660), .A2(new_n664), .ZN(G399));
  INV_X1    g0465(.A(new_n206), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(G41), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n588), .A2(G116), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G1), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n224), .B2(new_n668), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT28), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n637), .A2(new_n653), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT29), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT26), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n558), .A2(new_n633), .A3(new_n676), .A4(new_n570), .ZN(new_n677));
  INV_X1    g0477(.A(new_n597), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n678), .B1(new_n629), .B2(KEYINPUT26), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT93), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n677), .A2(new_n679), .A3(KEYINPUT93), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(new_n636), .A3(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n684), .A2(KEYINPUT29), .A3(new_n653), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n675), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n504), .A2(new_n491), .A3(new_n583), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT30), .ZN(new_n688));
  OR3_X1    g0488(.A1(new_n687), .A2(new_n688), .A3(new_n569), .ZN(new_n689));
  NOR3_X1   g0489(.A1(new_n491), .A2(new_n583), .A3(G179), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n567), .A2(new_n259), .ZN(new_n691));
  OAI211_X1 g0491(.A(new_n690), .B(new_n505), .C1(new_n691), .C2(new_n560), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n688), .B1(new_n687), .B2(new_n569), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n689), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n694), .A2(KEYINPUT31), .A3(new_n648), .ZN(new_n695));
  AOI21_X1  g0495(.A(KEYINPUT31), .B1(new_n694), .B2(new_n648), .ZN(new_n696));
  OAI21_X1  g0496(.A(KEYINPUT92), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n694), .A2(new_n648), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT31), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT92), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n694), .A2(KEYINPUT31), .A3(new_n648), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n697), .A2(new_n703), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n622), .A2(new_n528), .A3(new_n648), .ZN(new_n705));
  OAI21_X1  g0505(.A(G330), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n686), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n672), .B1(new_n708), .B2(G1), .ZN(G364));
  AOI21_X1  g0509(.A(new_n443), .B1(new_n641), .B2(G45), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n667), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n712), .B1(new_n651), .B2(G330), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n651), .A2(G330), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(G13), .A2(G33), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(G20), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT95), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n651), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n221), .B1(G20), .B2(new_n291), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OR3_X1    g0522(.A1(KEYINPUT98), .A2(G179), .A3(G200), .ZN(new_n723));
  OAI21_X1  g0523(.A(KEYINPUT98), .B1(G179), .B2(G200), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n607), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(new_n222), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n508), .ZN(new_n727));
  NAND2_X1  g0527(.A1(G20), .A2(G179), .ZN(new_n728));
  XOR2_X1   g0528(.A(new_n728), .B(KEYINPUT96), .Z(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G190), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n329), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n222), .A2(G190), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n734), .B1(new_n723), .B2(new_n724), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G159), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT32), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n732), .A2(new_n311), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n729), .A2(new_n607), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n329), .ZN(new_n742));
  AOI211_X1 g0542(.A(new_n727), .B(new_n740), .C1(G68), .C2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n329), .A2(G179), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(G20), .A3(G190), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G87), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n733), .A2(new_n744), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G107), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n747), .A2(new_n750), .A3(new_n278), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n751), .B1(new_n738), .B2(new_n739), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n730), .A2(G200), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n741), .A2(G200), .ZN(new_n754));
  AOI22_X1  g0554(.A1(G58), .A2(new_n753), .B1(new_n754), .B2(G77), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT97), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n743), .A2(new_n752), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g0557(.A(KEYINPUT33), .B(G317), .ZN(new_n758));
  AOI22_X1  g0558(.A1(G322), .A2(new_n753), .B1(new_n742), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n754), .A2(G311), .ZN(new_n760));
  INV_X1    g0560(.A(G303), .ZN(new_n761));
  INV_X1    g0561(.A(G283), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n745), .A2(new_n761), .B1(new_n748), .B2(new_n762), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n278), .B(new_n763), .C1(G329), .C2(new_n735), .ZN(new_n764));
  INV_X1    g0564(.A(new_n726), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n731), .A2(G326), .B1(new_n765), .B2(G294), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n759), .A2(new_n760), .A3(new_n764), .A4(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n722), .B1(new_n757), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n719), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n721), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT94), .ZN(new_n772));
  INV_X1    g0572(.A(new_n240), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n772), .B1(new_n773), .B2(new_n247), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n240), .A2(KEYINPUT94), .A3(G45), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n225), .A2(new_n247), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n380), .A2(new_n666), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n774), .A2(new_n775), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n495), .A2(new_n666), .ZN(new_n779));
  INV_X1    g0579(.A(G116), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n779), .A2(G355), .B1(new_n780), .B2(new_n666), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n771), .B1(new_n778), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n712), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n768), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n713), .A2(new_n715), .B1(new_n720), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(G396));
  OAI21_X1  g0586(.A(new_n358), .B1(new_n357), .B2(new_n653), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n365), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n363), .A2(new_n653), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n673), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n648), .B1(new_n635), .B2(new_n636), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n792), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n712), .B1(new_n797), .B2(new_n706), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(new_n706), .B2(new_n797), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n722), .A2(new_n717), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT99), .Z(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n783), .B1(new_n802), .B2(new_n202), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G116), .A2(new_n754), .B1(new_n742), .B2(G283), .ZN(new_n804));
  INV_X1    g0604(.A(G294), .ZN(new_n805));
  INV_X1    g0605(.A(new_n753), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n804), .B1(new_n805), .B2(new_n806), .C1(new_n761), .C2(new_n732), .ZN(new_n807));
  INV_X1    g0607(.A(G311), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n736), .A2(new_n808), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n495), .B1(new_n587), .B2(new_n748), .C1(new_n338), .C2(new_n745), .ZN(new_n810));
  NOR4_X1   g0610(.A1(new_n807), .A2(new_n727), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G58), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n726), .A2(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n746), .A2(G50), .B1(new_n749), .B2(G68), .ZN(new_n814));
  INV_X1    g0614(.A(G132), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n814), .B(new_n380), .C1(new_n815), .C2(new_n736), .ZN(new_n816));
  AOI22_X1  g0616(.A1(G143), .A2(new_n753), .B1(new_n742), .B2(G150), .ZN(new_n817));
  INV_X1    g0617(.A(G137), .ZN(new_n818));
  INV_X1    g0618(.A(new_n754), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n817), .B1(new_n818), .B2(new_n732), .C1(new_n737), .C2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT34), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n813), .B(new_n816), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n811), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n803), .B1(new_n722), .B2(new_n824), .C1(new_n792), .C2(new_n717), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n799), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G384));
  NOR2_X1   g0627(.A1(new_n536), .A2(new_n537), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT35), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n831), .A2(G116), .A3(new_n223), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT100), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n833), .B2(new_n832), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT36), .ZN(new_n836));
  OAI21_X1  g0636(.A(G77), .B1(new_n812), .B2(new_n309), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n837), .A2(new_n224), .B1(G50), .B2(new_n309), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n838), .A2(G1), .A3(new_n320), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT101), .Z(new_n840));
  AOI21_X1  g0640(.A(KEYINPUT7), .B1(new_n495), .B2(new_n222), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n374), .A2(new_n375), .ZN(new_n842));
  OAI21_X1  g0642(.A(G68), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(KEYINPUT16), .B1(new_n843), .B2(new_n370), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n388), .A2(new_n317), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n394), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n409), .A2(new_n408), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n848), .A2(new_n406), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT37), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n846), .A2(new_n646), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n849), .A2(KEYINPUT103), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n403), .A2(new_n405), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n846), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n854), .A2(new_n851), .A3(new_n850), .A4(new_n410), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT103), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n852), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT16), .B1(new_n387), .B2(new_n370), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n394), .B1(new_n845), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT102), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT102), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n862), .B(new_n394), .C1(new_n845), .C2(new_n859), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n861), .A2(new_n646), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n861), .A2(new_n853), .A3(new_n863), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n864), .A2(new_n865), .A3(new_n410), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT37), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n858), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n407), .A2(new_n411), .ZN(new_n869));
  INV_X1    g0669(.A(new_n864), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n868), .A2(KEYINPUT38), .A3(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n854), .A2(new_n851), .A3(new_n410), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n852), .A2(new_n857), .B1(KEYINPUT37), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n851), .B1(new_n407), .B2(new_n411), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n873), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n700), .A2(new_n702), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n792), .B1(new_n705), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n653), .A2(new_n326), .ZN(new_n882));
  AOI221_X4 g0682(.A(new_n882), .B1(new_n331), .B2(new_n332), .C1(new_n307), .C2(new_n327), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n307), .A2(new_n327), .A3(new_n648), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n878), .B(new_n881), .C1(new_n883), .C2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n882), .ZN(new_n887));
  INV_X1    g0687(.A(new_n288), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n287), .B1(new_n301), .B2(new_n258), .ZN(new_n889));
  OAI21_X1  g0689(.A(G169), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT14), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n289), .A2(new_n245), .A3(G169), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n303), .A2(G179), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT78), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n303), .A2(new_n294), .A3(G179), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n893), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n333), .B(new_n887), .C1(new_n897), .C2(new_n326), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n880), .B1(new_n898), .B2(new_n884), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n852), .A2(new_n857), .B1(new_n866), .B2(KEYINPUT37), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n864), .B1(new_n407), .B2(new_n411), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n873), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT40), .B1(new_n872), .B2(new_n902), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n886), .A2(KEYINPUT40), .B1(new_n899), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n705), .A2(new_n879), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n904), .A2(new_n442), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n899), .A2(new_n903), .ZN(new_n907));
  AOI221_X4 g0707(.A(new_n880), .B1(new_n872), .B2(new_n877), .C1(new_n898), .C2(new_n884), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT40), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(G330), .ZN(new_n911));
  AOI221_X4 g0711(.A(new_n440), .B1(new_n331), .B2(new_n332), .C1(new_n307), .C2(new_n327), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n912), .B(G330), .C1(new_n705), .C2(new_n879), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n906), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n407), .A2(new_n646), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n872), .A2(new_n902), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT39), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT39), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n872), .A2(new_n877), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n307), .A2(new_n327), .A3(new_n653), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT104), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n307), .A2(KEYINPUT104), .A3(new_n327), .A4(new_n653), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n915), .B1(new_n920), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n791), .B1(new_n795), .B2(new_n792), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n898), .B2(new_n884), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n916), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n914), .B(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT29), .B1(new_n637), .B2(new_n653), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n571), .A2(new_n611), .A3(new_n621), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n933), .A2(new_n528), .B1(new_n680), .B2(new_n681), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n648), .B1(new_n934), .B2(new_n683), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n932), .B1(new_n935), .B2(KEYINPUT29), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n936), .A2(new_n912), .A3(KEYINPUT105), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT105), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n686), .B2(new_n442), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n940), .A2(new_n628), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n931), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n443), .B2(new_n641), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n931), .A2(new_n941), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n836), .B(new_n840), .C1(new_n943), .C2(new_n944), .ZN(G367));
  AOI21_X1  g0745(.A(new_n771), .B1(new_n666), .B2(new_n347), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n235), .A2(new_n777), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n783), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n653), .A2(new_n601), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(new_n603), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n746), .A2(G58), .B1(new_n749), .B2(G77), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n952), .B(new_n278), .C1(new_n818), .C2(new_n736), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n731), .A2(G143), .B1(new_n765), .B2(G68), .ZN(new_n954));
  INV_X1    g0754(.A(new_n742), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n954), .B1(new_n415), .B2(new_n806), .C1(new_n737), .C2(new_n955), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n953), .B(new_n956), .C1(G50), .C2(new_n754), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT110), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n761), .A2(new_n806), .B1(new_n732), .B2(new_n808), .ZN(new_n959));
  INV_X1    g0759(.A(G317), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n736), .A2(new_n960), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n385), .B1(KEYINPUT109), .B2(KEYINPUT46), .C1(new_n508), .C2(new_n748), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n746), .A2(G116), .ZN(new_n963));
  NAND2_X1  g0763(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n963), .B(new_n964), .ZN(new_n965));
  NOR4_X1   g0765(.A1(new_n959), .A2(new_n961), .A3(new_n962), .A4(new_n965), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n754), .A2(G283), .B1(new_n765), .B2(G107), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n966), .B(new_n967), .C1(new_n805), .C2(new_n955), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n958), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n970), .A2(KEYINPUT47), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n721), .B1(new_n970), .B2(KEYINPUT47), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n948), .B1(new_n719), .B2(new_n951), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n632), .B1(new_n618), .B2(new_n620), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n662), .A2(new_n974), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n975), .A2(KEYINPUT42), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(KEYINPUT42), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n974), .B1(new_n556), .B2(new_n653), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n570), .A2(new_n648), .A3(new_n552), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n632), .B1(new_n980), .B2(new_n657), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n976), .B(new_n977), .C1(new_n648), .C2(new_n981), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n982), .A2(KEYINPUT106), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(KEYINPUT106), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n985), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n983), .A2(new_n986), .A3(new_n984), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n989), .A2(new_n660), .A3(new_n980), .A4(new_n990), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n991), .A2(KEYINPUT107), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n989), .A2(new_n990), .ZN(new_n993));
  INV_X1    g0793(.A(new_n660), .ZN(new_n994));
  INV_X1    g0794(.A(new_n980), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n993), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n991), .A2(KEYINPUT107), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n992), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n664), .A2(new_n995), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT44), .Z(new_n1000));
  NOR2_X1   g0800(.A1(new_n664), .A2(new_n995), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT45), .ZN(new_n1002));
  AND3_X1   g0802(.A1(new_n1000), .A2(new_n994), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n994), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(KEYINPUT108), .B1(new_n659), .B2(new_n661), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n652), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n652), .A2(new_n1007), .ZN(new_n1009));
  AND3_X1   g0809(.A1(new_n1008), .A2(new_n662), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n662), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n708), .B1(new_n1006), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n667), .B(KEYINPUT41), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n711), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n973), .B1(new_n998), .B2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT111), .Z(G387));
  INV_X1    g0817(.A(new_n777), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n231), .B2(G45), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n669), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1019), .B1(new_n1020), .B2(new_n779), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n344), .A2(G50), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT112), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n1023), .A2(KEYINPUT50), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1023), .A2(KEYINPUT50), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n669), .B(new_n247), .C1(new_n309), .C2(new_n202), .ZN(new_n1026));
  NOR3_X1   g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n1021), .A2(new_n1027), .B1(G107), .B2(new_n206), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n783), .B1(new_n1028), .B2(new_n770), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n765), .A2(new_n347), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n806), .B2(new_n311), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT113), .ZN(new_n1032));
  AND2_X1   g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n745), .A2(new_n202), .B1(new_n748), .B2(new_n508), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n385), .B(new_n1035), .C1(G150), .C2(new_n735), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n737), .B2(new_n732), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n309), .A2(new_n819), .B1(new_n955), .B2(new_n392), .ZN(new_n1038));
  NOR4_X1   g0838(.A1(new_n1033), .A2(new_n1034), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G303), .A2(new_n754), .B1(new_n731), .B2(G322), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n808), .B2(new_n955), .C1(new_n960), .C2(new_n806), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT48), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n762), .B2(new_n726), .C1(new_n805), .C2(new_n745), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT49), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n735), .A2(G326), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1046), .B(new_n385), .C1(new_n780), .C2(new_n748), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1039), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1029), .B1(new_n1049), .B2(new_n722), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n659), .B2(new_n769), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1012), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1051), .B1(new_n1052), .B2(new_n711), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1012), .A2(new_n707), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n667), .B(KEYINPUT114), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1052), .A2(new_n708), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1053), .B1(new_n1058), .B2(new_n1059), .ZN(G393));
  OAI211_X1 g0860(.A(new_n495), .B(new_n750), .C1(new_n762), .C2(new_n745), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n726), .A2(new_n780), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(G322), .C2(new_n735), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1063), .B1(new_n805), .B2(new_n819), .C1(new_n761), .C2(new_n955), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G311), .A2(new_n753), .B1(new_n731), .B2(G317), .ZN(new_n1065));
  XOR2_X1   g0865(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n1066));
  XNOR2_X1  g0866(.A(new_n1065), .B(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1069), .A2(KEYINPUT116), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT116), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n380), .B1(new_n309), .B2(new_n745), .C1(new_n587), .C2(new_n748), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n955), .A2(new_n311), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1072), .B(new_n1073), .C1(G143), .C2(new_n735), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n415), .A2(new_n732), .B1(new_n806), .B2(new_n737), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT51), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n726), .A2(new_n202), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n344), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1078), .B1(new_n1079), .B2(new_n754), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1074), .A2(new_n1077), .A3(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n1068), .A2(new_n1071), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n721), .B1(new_n1070), .B2(new_n1083), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n770), .B1(new_n508), .B2(new_n206), .C1(new_n243), .C2(new_n1018), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1084), .A2(new_n712), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n995), .B2(new_n769), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n1005), .B2(new_n711), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1057), .B1(new_n1006), .B2(new_n1055), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1005), .A2(new_n1054), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(G390));
  NAND2_X1  g0891(.A1(new_n898), .A2(new_n884), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n684), .A2(new_n653), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n790), .B1(new_n1093), .B2(new_n789), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n923), .A2(new_n924), .A3(new_n878), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n872), .A2(new_n877), .A3(new_n918), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n918), .B1(new_n872), .B2(new_n902), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n928), .B2(new_n925), .ZN(new_n1101));
  OAI211_X1 g0901(.A(G330), .B(new_n792), .C1(new_n704), .C2(new_n705), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1092), .A2(new_n1103), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n1097), .A2(new_n1101), .A3(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1092), .A2(G330), .A3(new_n881), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n711), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(G97), .A2(new_n754), .B1(new_n742), .B2(G107), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1110), .B1(new_n780), .B2(new_n806), .C1(new_n762), .C2(new_n732), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n736), .A2(new_n805), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n747), .B(new_n495), .C1(new_n309), .C2(new_n748), .ZN(new_n1113));
  NOR4_X1   g0913(.A1(new_n1111), .A2(new_n1078), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  XOR2_X1   g0914(.A(KEYINPUT54), .B(G143), .Z(new_n1115));
  AOI22_X1  g0915(.A1(G128), .A2(new_n731), .B1(new_n754), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n818), .B2(new_n955), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n745), .A2(new_n415), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT53), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n735), .A2(G125), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n495), .B1(G50), .B2(new_n749), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n806), .A2(new_n815), .B1(new_n737), .B2(new_n726), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n1117), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n721), .B1(new_n1114), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n783), .B1(new_n802), .B2(new_n392), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1125), .B(new_n1126), .C1(new_n920), .C2(new_n717), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1109), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT117), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1102), .A2(new_n898), .A3(new_n884), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1106), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n927), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n307), .A2(new_n327), .B1(new_n331), .B2(new_n332), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n307), .A2(new_n327), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1134), .A2(new_n887), .B1(new_n1135), .B2(new_n648), .ZN(new_n1136));
  OAI211_X1 g0936(.A(G330), .B(new_n792), .C1(new_n705), .C2(new_n879), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1094), .B1(new_n1092), .B2(new_n1103), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1132), .A2(new_n1133), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n940), .A2(new_n628), .A3(new_n913), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1130), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1139), .A2(new_n1138), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(G330), .A2(new_n899), .B1(new_n1136), .B2(new_n1102), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1143), .B1(new_n1144), .B2(new_n927), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n940), .A2(new_n628), .A3(new_n913), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1145), .A2(new_n1146), .A3(KEYINPUT117), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1108), .B1(new_n1142), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1141), .B1(new_n1149), .B2(new_n1143), .ZN(new_n1150));
  AOI21_X1  g0950(.A(KEYINPUT118), .B1(new_n1108), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1057), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  AOI211_X1 g0952(.A(KEYINPUT118), .B(new_n1108), .C1(new_n1142), .C2(new_n1147), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1129), .B1(new_n1152), .B2(new_n1153), .ZN(G378));
  AOI21_X1  g0954(.A(KEYINPUT122), .B1(new_n926), .B2(new_n929), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n439), .B(KEYINPUT55), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n418), .A2(new_n646), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1157), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1163), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1157), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n1165), .A2(new_n1166), .A3(new_n1161), .ZN(new_n1167));
  OR2_X1    g0967(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n910), .B2(G330), .ZN(new_n1169));
  INV_X1    g0969(.A(G330), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n904), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1156), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1171), .B1(new_n904), .B2(new_n1170), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n907), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n909), .B1(new_n899), .B2(new_n878), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1168), .B(G330), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1174), .A2(new_n1155), .A3(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1173), .A2(new_n711), .A3(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(G97), .A2(new_n742), .B1(new_n754), .B2(new_n347), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT119), .Z(new_n1181));
  NOR2_X1   g0981(.A1(new_n748), .A2(new_n812), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(G77), .B2(new_n746), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n380), .A2(G41), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(new_n762), .C2(new_n736), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n731), .A2(G116), .B1(new_n765), .B2(G68), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n338), .B2(new_n806), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n1181), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT120), .Z(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(KEYINPUT58), .ZN(new_n1190));
  AOI211_X1 g0990(.A(G50), .B(new_n1184), .C1(new_n263), .C2(new_n246), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n263), .B(new_n246), .C1(new_n748), .C2(new_n737), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(G128), .A2(new_n753), .B1(new_n754), .B2(G137), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n731), .A2(G125), .B1(new_n746), .B2(new_n1115), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n742), .A2(G132), .B1(new_n765), .B2(G150), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n1196), .A2(KEYINPUT59), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1192), .B(new_n1197), .C1(G124), .C2(new_n735), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1196), .A2(KEYINPUT59), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1191), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1190), .A2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1189), .A2(KEYINPUT58), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n721), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n783), .B1(new_n802), .B2(new_n311), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(new_n1168), .C2(new_n717), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1179), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1106), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1133), .B1(new_n883), .B2(new_n885), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n923), .A2(new_n924), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n920), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n923), .A2(new_n924), .A3(new_n878), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1208), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1097), .A2(new_n1101), .A3(new_n1104), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1146), .B1(new_n1216), .B2(new_n1140), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n930), .ZN(new_n1218));
  AND3_X1   g1018(.A1(new_n1174), .A2(new_n1218), .A3(new_n1177), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1218), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1217), .B(KEYINPUT57), .C1(new_n1219), .C2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n1057), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1174), .A2(new_n1155), .A3(new_n1177), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1155), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(KEYINPUT57), .B1(new_n1225), .B2(new_n1217), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1207), .B1(new_n1222), .B2(new_n1226), .ZN(G375));
  NAND2_X1  g1027(.A1(new_n1142), .A2(new_n1147), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1228), .A2(new_n1014), .A3(new_n1229), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(G283), .A2(new_n753), .B1(new_n731), .B2(G294), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1231), .B1(new_n338), .B2(new_n819), .C1(new_n780), .C2(new_n955), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n735), .A2(G303), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n746), .A2(G97), .B1(new_n749), .B2(G77), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1030), .A2(new_n495), .A3(new_n1233), .A4(new_n1234), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n731), .A2(G132), .B1(new_n765), .B2(G50), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n818), .B2(new_n806), .C1(new_n415), .C2(new_n819), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n742), .A2(new_n1115), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n735), .A2(G128), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1182), .B1(G159), .B2(new_n746), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1238), .A2(new_n380), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n1232), .A2(new_n1235), .B1(new_n1237), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n721), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1243), .B(new_n712), .C1(G68), .C2(new_n801), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n1136), .B2(new_n716), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(new_n1145), .B2(new_n711), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1230), .A2(new_n1246), .ZN(G381));
  OAI211_X1 g1047(.A(new_n785), .B(new_n1053), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1248));
  OR2_X1    g1048(.A1(new_n1248), .A2(G384), .ZN(new_n1249));
  NOR4_X1   g1049(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(G375), .A2(G378), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(G407));
  INV_X1    g1052(.A(G343), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(G213), .ZN(new_n1254));
  XOR2_X1   g1054(.A(new_n1254), .B(KEYINPUT123), .Z(new_n1255));
  NAND2_X1  g1055(.A1(new_n1251), .A2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(G407), .A2(G213), .A3(new_n1256), .ZN(G409));
  NAND2_X1  g1057(.A1(G393), .A2(G396), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1248), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(G390), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT111), .B1(new_n1258), .B2(new_n1248), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1260), .B1(new_n1261), .B2(G390), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1016), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1016), .B(new_n1260), .C1(G390), .C2(new_n1261), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n711), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1205), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT125), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1217), .A2(new_n1178), .A3(new_n1173), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n1268), .A2(new_n1269), .B1(new_n1270), .B2(new_n1014), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1267), .A2(KEYINPUT125), .A3(new_n1205), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1228), .A2(new_n1216), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1145), .A2(new_n1214), .A3(new_n1146), .A4(new_n1215), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT118), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1056), .B1(new_n1274), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1148), .A2(new_n1276), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1128), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1273), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT124), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n930), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1174), .A2(new_n1218), .A3(new_n1177), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT57), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1286), .B1(new_n1275), .B2(new_n1146), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1056), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1217), .A2(new_n1173), .A3(new_n1178), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1286), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  AND4_X1   g1091(.A1(new_n1282), .A2(G378), .A3(new_n1291), .A4(new_n1207), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1206), .B1(new_n1288), .B2(new_n1290), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1282), .B1(new_n1293), .B2(G378), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1281), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1255), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT126), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1229), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(KEYINPUT60), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT60), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1229), .A2(new_n1297), .A3(new_n1300), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1150), .A2(new_n1056), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1299), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1303), .A2(G384), .A3(new_n1246), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(G384), .B1(new_n1303), .B2(new_n1246), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1295), .A2(new_n1296), .A3(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(KEYINPUT62), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT62), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1295), .A2(new_n1310), .A3(new_n1296), .A4(new_n1307), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1309), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1303), .A2(new_n1246), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n826), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1255), .A2(G2897), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1314), .A2(new_n1304), .A3(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1315), .B1(new_n1314), .B2(new_n1304), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(G378), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1319));
  OAI21_X1  g1119(.A(KEYINPUT124), .B1(G375), .B2(new_n1280), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1293), .A2(new_n1282), .A3(G378), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1319), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1318), .B1(new_n1322), .B2(new_n1255), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT61), .ZN(new_n1324));
  AOI21_X1  g1124(.A(KEYINPUT127), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1266), .B1(new_n1312), .B2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1308), .A2(KEYINPUT63), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1266), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT63), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1295), .A2(new_n1329), .A3(new_n1296), .A4(new_n1307), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1327), .A2(new_n1328), .A3(new_n1330), .ZN(new_n1331));
  OR2_X1    g1131(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1332), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1333));
  AOI21_X1  g1133(.A(KEYINPUT127), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1334));
  NOR3_X1   g1134(.A1(new_n1333), .A2(new_n1334), .A3(KEYINPUT61), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1331), .A2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1326), .A2(new_n1336), .ZN(G405));
  NAND2_X1  g1137(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(G375), .A2(new_n1280), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  XNOR2_X1  g1140(.A(new_n1340), .B(new_n1307), .ZN(new_n1341));
  XNOR2_X1  g1141(.A(new_n1341), .B(new_n1266), .ZN(G402));
endmodule


