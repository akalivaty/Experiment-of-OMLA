//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  XNOR2_X1  g000(.A(KEYINPUT2), .B(G113), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(G116), .B(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  XOR2_X1   g004(.A(G116), .B(G119), .Z(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(new_n187), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G143), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G146), .ZN(new_n197));
  AND2_X1   g011(.A1(KEYINPUT0), .A2(G128), .ZN(new_n198));
  AND3_X1   g012(.A1(new_n195), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n200), .B1(new_n196), .B2(G146), .ZN(new_n201));
  NOR3_X1   g015(.A1(new_n194), .A2(KEYINPUT64), .A3(G143), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n195), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT0), .A2(G128), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n198), .A2(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n199), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT11), .ZN(new_n207));
  INV_X1    g021(.A(G134), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(G137), .ZN(new_n209));
  INV_X1    g023(.A(G137), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT11), .A3(G134), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n208), .A2(G137), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G131), .ZN(new_n214));
  AOI21_X1  g028(.A(G131), .B1(new_n208), .B2(G137), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n209), .A2(new_n215), .A3(new_n211), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n193), .B1(new_n206), .B2(new_n217), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n209), .A2(new_n215), .A3(new_n211), .ZN(new_n219));
  INV_X1    g033(.A(G131), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n210), .A2(G134), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(new_n212), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G128), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(new_n195), .A3(new_n197), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n196), .A2(G146), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT64), .B1(new_n194), .B2(G143), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n200), .A2(new_n196), .A3(G146), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n224), .B1(new_n195), .B2(KEYINPUT1), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n226), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n223), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(KEYINPUT28), .B1(new_n218), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n235), .B1(new_n219), .B2(new_n222), .ZN(new_n236));
  INV_X1    g050(.A(new_n222), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(new_n216), .A3(KEYINPUT65), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n232), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n206), .A2(new_n217), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n193), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n225), .A2(new_n195), .A3(new_n197), .ZN(new_n243));
  INV_X1    g057(.A(new_n231), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n243), .B1(new_n203), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n237), .A2(new_n216), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT67), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT67), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n223), .A2(new_n232), .A3(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n218), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n242), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n234), .B1(new_n251), .B2(KEYINPUT28), .ZN(new_n252));
  NOR2_X1   g066(.A1(G237), .A2(G953), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G210), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n254), .B(KEYINPUT27), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT26), .B(G101), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n255), .B(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT66), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT30), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n260), .B1(new_n241), .B2(new_n261), .ZN(new_n262));
  AOI211_X1 g076(.A(KEYINPUT66), .B(KEYINPUT30), .C1(new_n239), .C2(new_n240), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n247), .A2(KEYINPUT30), .A3(new_n240), .A4(new_n249), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n193), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT68), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n265), .A2(new_n193), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT68), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n268), .B(new_n269), .C1(new_n263), .C2(new_n262), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n250), .A2(KEYINPUT69), .A3(new_n257), .ZN(new_n272));
  AOI21_X1  g086(.A(KEYINPUT69), .B1(new_n250), .B2(new_n257), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT31), .B1(new_n271), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT31), .ZN(new_n277));
  AOI211_X1 g091(.A(new_n277), .B(new_n274), .C1(new_n267), .C2(new_n270), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n259), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(G472), .A2(G902), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT32), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT29), .B1(new_n252), .B2(new_n257), .ZN(new_n284));
  INV_X1    g098(.A(new_n250), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n285), .B1(new_n267), .B2(new_n270), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n284), .B1(new_n286), .B2(new_n257), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n247), .A2(new_n240), .A3(new_n249), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n193), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n250), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n234), .B1(new_n290), .B2(KEYINPUT28), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n257), .A2(KEYINPUT29), .ZN(new_n292));
  AOI21_X1  g106(.A(G902), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n287), .A2(new_n293), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n279), .A2(new_n283), .B1(new_n294), .B2(G472), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT30), .B1(new_n239), .B2(new_n240), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n296), .B(new_n260), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n269), .B1(new_n297), .B2(new_n268), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n264), .A2(KEYINPUT68), .A3(new_n266), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n275), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n277), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n274), .B1(new_n267), .B2(new_n270), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT31), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n258), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n282), .B1(new_n304), .B2(new_n281), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n295), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(G214), .B1(G237), .B2(G902), .ZN(new_n307));
  INV_X1    g121(.A(G953), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n308), .A2(G952), .ZN(new_n309));
  NAND2_X1  g123(.A1(G234), .A2(G237), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n310), .A2(G902), .A3(G953), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT21), .B(G898), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n312), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(G110), .B(G122), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n318), .B(KEYINPUT78), .ZN(new_n319));
  INV_X1    g133(.A(G104), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G107), .ZN(new_n321));
  INV_X1    g135(.A(G107), .ZN(new_n322));
  AND3_X1   g136(.A1(new_n322), .A2(KEYINPUT3), .A3(G104), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT3), .B1(new_n322), .B2(G104), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n321), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G101), .ZN(new_n326));
  INV_X1    g140(.A(G101), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n327), .B(new_n321), .C1(new_n323), .C2(new_n324), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n326), .A2(KEYINPUT4), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT77), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT4), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n325), .A2(new_n331), .A3(G101), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n329), .A2(new_n330), .A3(new_n193), .A4(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT73), .B1(new_n322), .B2(G104), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT73), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(new_n320), .A3(G107), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n322), .A2(G104), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n334), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G101), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n339), .A2(new_n328), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT5), .ZN(new_n341));
  INV_X1    g155(.A(G119), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n342), .A3(G116), .ZN(new_n343));
  OAI211_X1 g157(.A(G113), .B(new_n343), .C1(new_n191), .C2(new_n341), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n340), .A2(new_n190), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n333), .A2(new_n345), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n193), .A2(new_n332), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n330), .B1(new_n347), .B2(new_n329), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n319), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n328), .A2(KEYINPUT4), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT3), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n337), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n322), .A2(KEYINPUT3), .A3(G104), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n327), .B1(new_n354), .B2(new_n321), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n193), .B(new_n332), .C1(new_n350), .C2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT77), .ZN(new_n357));
  INV_X1    g171(.A(new_n319), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n357), .A2(new_n333), .A3(new_n358), .A4(new_n345), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n349), .A2(KEYINPUT6), .A3(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(G143), .B(G146), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n198), .ZN(new_n362));
  OR2_X1    g176(.A1(new_n198), .A2(new_n204), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n362), .B1(new_n230), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT79), .B1(new_n364), .B2(G125), .ZN(new_n365));
  INV_X1    g179(.A(G125), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n366), .B(new_n226), .C1(new_n230), .C2(new_n231), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n367), .B1(new_n206), .B2(new_n366), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n365), .B1(new_n368), .B2(KEYINPUT79), .ZN(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT80), .B(G224), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n308), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT81), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n370), .A2(KEYINPUT81), .A3(new_n308), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n369), .B(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT6), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n378), .B(new_n319), .C1(new_n346), .C2(new_n348), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n360), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G902), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n373), .A2(KEYINPUT7), .A3(new_n374), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT82), .B1(new_n369), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT79), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n364), .A2(G125), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n385), .B1(new_n386), .B2(new_n367), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT82), .ZN(new_n388));
  NOR4_X1   g202(.A1(new_n387), .A2(new_n388), .A3(new_n365), .A4(new_n382), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  XOR2_X1   g204(.A(new_n319), .B(KEYINPUT8), .Z(new_n391));
  NAND2_X1  g205(.A1(new_n344), .A2(new_n190), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n339), .A2(new_n328), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n345), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n382), .B1(new_n387), .B2(new_n365), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n359), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n381), .B1(new_n390), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(G210), .B1(G237), .B2(G902), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n380), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n400), .B(KEYINPUT83), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  OR2_X1    g218(.A1(new_n384), .A2(new_n389), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n359), .A2(new_n396), .A3(new_n397), .ZN(new_n406));
  AOI21_X1  g220(.A(G902), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n360), .A2(new_n377), .A3(new_n379), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n404), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n307), .B(new_n317), .C1(new_n402), .C2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(G128), .A3(new_n196), .ZN(new_n412));
  XNOR2_X1  g226(.A(G128), .B(G143), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n412), .B(G134), .C1(new_n414), .C2(new_n411), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n208), .ZN(new_n416));
  XNOR2_X1  g230(.A(G116), .B(G122), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n417), .B(new_n322), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n415), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n413), .B(new_n208), .ZN(new_n420));
  INV_X1    g234(.A(G116), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(KEYINPUT14), .A3(G122), .ZN(new_n422));
  INV_X1    g236(.A(new_n417), .ZN(new_n423));
  OAI211_X1 g237(.A(G107), .B(new_n422), .C1(new_n423), .C2(KEYINPUT14), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n417), .A2(new_n322), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n420), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n419), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT9), .B(G234), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(G217), .A3(new_n308), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n427), .A2(new_n430), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n381), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AND2_X1   g247(.A1(KEYINPUT92), .A2(KEYINPUT15), .ZN(new_n434));
  NOR2_X1   g248(.A1(KEYINPUT92), .A2(KEYINPUT15), .ZN(new_n435));
  OAI21_X1  g249(.A(G478), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n433), .B(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G237), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(new_n308), .A3(G214), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n196), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n253), .A2(G143), .A3(G214), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT86), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(new_n444), .A3(G131), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n444), .B1(new_n443), .B2(G131), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT17), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n440), .A2(new_n196), .ZN(new_n449));
  AOI21_X1  g263(.A(G143), .B1(new_n253), .B2(G214), .ZN(new_n450));
  OAI21_X1  g264(.A(G131), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT86), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n441), .A2(new_n220), .A3(new_n442), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT17), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n452), .A2(new_n453), .A3(new_n454), .A4(new_n445), .ZN(new_n455));
  INV_X1    g269(.A(G140), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(G125), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n366), .A2(G140), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT16), .ZN(new_n459));
  OR3_X1    g273(.A1(new_n366), .A2(KEYINPUT16), .A3(G140), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n194), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n459), .A2(new_n460), .A3(G146), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n448), .A2(new_n455), .A3(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(G113), .B(G122), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(new_n320), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n457), .A2(new_n458), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G146), .ZN(new_n470));
  XNOR2_X1  g284(.A(G125), .B(G140), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n194), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT84), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n470), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n473), .B1(new_n470), .B2(new_n472), .ZN(new_n475));
  OR2_X1    g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT85), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n441), .A2(new_n477), .A3(new_n442), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(KEYINPUT18), .A3(G131), .ZN(new_n479));
  NAND2_X1  g293(.A1(KEYINPUT18), .A2(G131), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n441), .A2(new_n477), .A3(new_n442), .A4(new_n480), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n466), .A2(new_n468), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n474), .A2(new_n475), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n479), .A2(new_n481), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n452), .A2(new_n445), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n464), .B1(new_n489), .B2(KEYINPUT17), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n488), .B1(new_n490), .B2(new_n455), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT90), .B1(new_n491), .B2(new_n468), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n466), .A2(new_n483), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT90), .ZN(new_n494));
  INV_X1    g308(.A(new_n468), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n485), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(G475), .B1(new_n497), .B2(G902), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT88), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT19), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n469), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(KEYINPUT19), .B1(new_n457), .B2(new_n458), .ZN(new_n502));
  OAI211_X1 g316(.A(KEYINPUT87), .B(new_n194), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n463), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n469), .A2(new_n500), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n471), .A2(KEYINPUT19), .ZN(new_n506));
  AOI21_X1  g320(.A(G146), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n507), .A2(KEYINPUT87), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n452), .A2(new_n453), .A3(new_n445), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n509), .A2(new_n510), .B1(new_n476), .B2(new_n482), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n499), .B1(new_n511), .B2(new_n468), .ZN(new_n512));
  OR2_X1    g326(.A1(new_n507), .A2(KEYINPUT87), .ZN(new_n513));
  INV_X1    g327(.A(new_n463), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n514), .B1(new_n507), .B2(KEYINPUT87), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n513), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n483), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n517), .A2(KEYINPUT88), .A3(new_n495), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n512), .A2(new_n484), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT20), .ZN(new_n520));
  NOR2_X1   g334(.A1(G475), .A2(G902), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(KEYINPUT89), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n520), .B1(new_n519), .B2(new_n522), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n498), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n410), .A2(new_n438), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n342), .A2(G128), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n224), .A2(KEYINPUT23), .A3(G119), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n342), .A2(G128), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n527), .B(new_n528), .C1(new_n529), .C2(KEYINPUT23), .ZN(new_n530));
  XOR2_X1   g344(.A(KEYINPUT24), .B(G110), .Z(new_n531));
  XNOR2_X1  g345(.A(G119), .B(G128), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n530), .A2(G110), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n464), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT70), .B(G110), .ZN(new_n535));
  OAI22_X1  g349(.A1(new_n530), .A2(new_n535), .B1(new_n531), .B2(new_n532), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(new_n463), .A3(new_n472), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT22), .B(G137), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n308), .A2(G221), .A3(G234), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n538), .B(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT71), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT25), .ZN(new_n544));
  AOI21_X1  g358(.A(G902), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n543), .A2(new_n544), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(G234), .ZN(new_n549));
  OAI21_X1  g363(.A(G217), .B1(new_n549), .B2(G902), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n550), .B1(new_n546), .B2(new_n547), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n542), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n550), .A2(new_n381), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(G221), .B1(new_n428), .B2(G902), .ZN(new_n557));
  XOR2_X1   g371(.A(new_n557), .B(KEYINPUT72), .Z(new_n558));
  INV_X1    g372(.A(G469), .ZN(new_n559));
  XNOR2_X1  g373(.A(G110), .B(G140), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n308), .A2(G227), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n560), .B(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n206), .B(new_n332), .C1(new_n355), .C2(new_n350), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n226), .B1(new_n231), .B2(new_n361), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(new_n339), .A3(new_n328), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT10), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n232), .A2(KEYINPUT10), .A3(new_n328), .A4(new_n339), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n564), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n217), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT75), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT75), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n570), .A2(new_n573), .A3(new_n217), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n217), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n564), .A2(new_n576), .A3(new_n568), .A4(new_n569), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n563), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n566), .B1(new_n340), .B2(new_n232), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n576), .A2(KEYINPUT74), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT12), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT12), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n579), .A2(new_n580), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n577), .A2(new_n563), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n559), .B(new_n381), .C1(new_n578), .C2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT76), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n570), .A2(new_n573), .A3(new_n217), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n573), .B1(new_n570), .B2(new_n217), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n577), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n562), .ZN(new_n594));
  INV_X1    g408(.A(new_n587), .ZN(new_n595));
  AOI21_X1  g409(.A(G902), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(KEYINPUT76), .A3(new_n559), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n590), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n586), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n575), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n577), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n562), .B1(new_n585), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(G469), .B1(new_n604), .B2(G902), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n558), .B1(new_n598), .B2(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n306), .A2(new_n526), .A3(new_n556), .A4(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT93), .B(G101), .Z(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G3));
  NAND2_X1  g423(.A1(new_n279), .A2(new_n381), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n610), .A2(G472), .B1(new_n280), .B2(new_n279), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n606), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n612), .A2(new_n555), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n307), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n401), .B1(new_n380), .B2(new_n399), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n407), .A2(new_n408), .A3(new_n400), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n317), .ZN(new_n619));
  INV_X1    g433(.A(G478), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n433), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT95), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT94), .B1(new_n431), .B2(new_n432), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT33), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI211_X1 g439(.A(KEYINPUT94), .B(KEYINPUT33), .C1(new_n431), .C2(new_n432), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n627), .A2(G478), .A3(new_n381), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n622), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n525), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n619), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n614), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT34), .B(G104), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  OAI211_X1 g448(.A(new_n498), .B(new_n438), .C1(new_n523), .C2(new_n524), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n619), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n614), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT35), .B(G107), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G9));
  INV_X1    g453(.A(KEYINPUT36), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n541), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT96), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT97), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n642), .A2(KEYINPUT97), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n538), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OR2_X1    g460(.A1(new_n642), .A2(KEYINPUT97), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n647), .A2(new_n534), .A3(new_n537), .A4(new_n643), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n554), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n552), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n611), .A2(new_n526), .A3(new_n606), .A4(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  NAND2_X1  g469(.A1(new_n518), .A2(new_n484), .ZN(new_n656));
  AOI21_X1  g470(.A(KEYINPUT88), .B1(new_n517), .B2(new_n495), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n522), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT20), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(G900), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n314), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n311), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n661), .A2(new_n438), .A3(new_n498), .A4(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n400), .B1(new_n407), .B2(new_n408), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n307), .B1(new_n402), .B2(new_n666), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n665), .A2(new_n667), .A3(KEYINPUT98), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(KEYINPUT98), .B1(new_n665), .B2(new_n667), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n671), .A2(new_n306), .A3(new_n606), .A4(new_n652), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT99), .B(G128), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G30));
  NAND2_X1  g488(.A1(new_n279), .A2(new_n283), .ZN(new_n675));
  INV_X1    g489(.A(new_n257), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n290), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT101), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n381), .B1(new_n678), .B2(new_n302), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(G472), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(KEYINPUT32), .B1(new_n279), .B2(new_n280), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n402), .A2(new_n409), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n437), .B1(new_n661), .B2(new_n498), .ZN(new_n687));
  INV_X1    g501(.A(new_n652), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n687), .A2(new_n307), .A3(new_n688), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n683), .A2(new_n686), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n664), .B(KEYINPUT39), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n606), .A2(new_n691), .ZN(new_n692));
  OR2_X1    g506(.A1(new_n692), .A2(KEYINPUT40), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(KEYINPUT40), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n690), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT102), .B(G143), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G45));
  OAI211_X1 g511(.A(new_n652), .B(new_n307), .C1(new_n402), .C2(new_n666), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n525), .A2(new_n629), .A3(new_n664), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n284), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n250), .B1(new_n298), .B2(new_n299), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n701), .B1(new_n702), .B2(new_n676), .ZN(new_n703));
  INV_X1    g517(.A(new_n293), .ZN(new_n704));
  OAI21_X1  g518(.A(G472), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n675), .A2(new_n705), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n700), .B(new_n606), .C1(new_n706), .C2(new_n682), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G146), .ZN(G48));
  AOI21_X1  g522(.A(new_n555), .B1(new_n295), .B2(new_n305), .ZN(new_n709));
  INV_X1    g523(.A(new_n558), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n587), .B1(new_n562), .B2(new_n593), .ZN(new_n711));
  OAI21_X1  g525(.A(G469), .B1(new_n711), .B2(G902), .ZN(new_n712));
  AOI21_X1  g526(.A(KEYINPUT76), .B1(new_n596), .B2(new_n559), .ZN(new_n713));
  NOR4_X1   g527(.A1(new_n711), .A2(new_n589), .A3(G469), .A4(G902), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n710), .B(new_n712), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n709), .A2(new_n631), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  NAND4_X1  g533(.A1(new_n306), .A2(new_n716), .A3(new_n636), .A4(new_n556), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT103), .B(G116), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G18));
  NOR2_X1   g536(.A1(new_n715), .A2(new_n667), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n525), .A2(new_n438), .A3(new_n316), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n306), .A2(new_n723), .A3(new_n652), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G119), .ZN(G21));
  OR2_X1    g540(.A1(new_n291), .A2(KEYINPUT104), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n291), .A2(KEYINPUT104), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n676), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n729), .B1(new_n276), .B2(new_n278), .ZN(new_n730));
  AOI22_X1  g544(.A1(new_n610), .A2(G472), .B1(new_n280), .B2(new_n730), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n687), .A2(new_n317), .A3(new_n618), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n731), .A2(new_n732), .A3(new_n556), .A4(new_n716), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G122), .ZN(G24));
  NAND2_X1  g548(.A1(new_n610), .A2(G472), .ZN(new_n735));
  INV_X1    g549(.A(new_n699), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n730), .A2(new_n280), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n735), .A2(new_n736), .A3(new_n652), .A4(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n723), .ZN(new_n739));
  OR2_X1    g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G125), .ZN(G27));
  OAI211_X1 g555(.A(new_n556), .B(new_n606), .C1(new_n706), .C2(new_n682), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n684), .A2(new_n307), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(KEYINPUT42), .A3(new_n736), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT42), .ZN(new_n746));
  INV_X1    g560(.A(new_n743), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n306), .A2(new_n556), .A3(new_n606), .A4(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n746), .B1(new_n748), .B2(new_n699), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G131), .ZN(G33));
  NOR2_X1   g565(.A1(new_n748), .A2(new_n665), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n208), .ZN(G36));
  INV_X1    g567(.A(new_n629), .ZN(new_n754));
  OR3_X1    g568(.A1(new_n754), .A2(KEYINPUT43), .A3(new_n525), .ZN(new_n755));
  OAI21_X1  g569(.A(KEYINPUT43), .B1(new_n754), .B2(new_n525), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n612), .A2(KEYINPUT106), .A3(new_n652), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT106), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n759), .B1(new_n611), .B2(new_n688), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n757), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n761), .A2(KEYINPUT44), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(KEYINPUT44), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n559), .A2(new_n381), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n603), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT105), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n559), .B1(new_n603), .B2(new_n765), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n764), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n598), .B1(new_n770), .B2(KEYINPUT46), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT46), .ZN(new_n772));
  AOI211_X1 g586(.A(new_n772), .B(new_n764), .C1(new_n768), .C2(new_n769), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n710), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n691), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n762), .A2(new_n763), .A3(new_n743), .A4(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(new_n210), .ZN(G39));
  NOR4_X1   g592(.A1(new_n306), .A2(new_n556), .A3(new_n699), .A4(new_n743), .ZN(new_n779));
  XOR2_X1   g593(.A(new_n779), .B(KEYINPUT108), .Z(new_n780));
  XNOR2_X1  g594(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n710), .B(new_n781), .C1(new_n771), .C2(new_n773), .ZN(new_n782));
  INV_X1    g596(.A(new_n781), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n774), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n780), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(new_n456), .ZN(G42));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n787));
  NOR2_X1   g601(.A1(G952), .A2(G953), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n715), .A2(new_n743), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n683), .A2(new_n312), .A3(new_n556), .A4(new_n789), .ZN(new_n790));
  OR3_X1    g604(.A1(new_n790), .A2(new_n525), .A3(new_n629), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n735), .A2(new_n737), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n688), .ZN(new_n793));
  INV_X1    g607(.A(new_n757), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n793), .A2(new_n794), .A3(new_n312), .A4(new_n789), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n791), .A2(new_n795), .A3(KEYINPUT51), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n794), .A2(new_n312), .A3(new_n556), .A4(new_n731), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n686), .A2(new_n615), .A3(new_n716), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NOR4_X1   g614(.A1(new_n757), .A2(new_n792), .A3(new_n311), .A4(new_n555), .ZN(new_n801));
  INV_X1    g615(.A(new_n799), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(KEYINPUT50), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n798), .A2(new_n743), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n598), .A2(new_n558), .A3(new_n712), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n784), .A2(new_n782), .A3(new_n807), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n796), .B(new_n804), .C1(new_n806), .C2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT114), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT51), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n791), .A2(new_n795), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n812), .B1(new_n804), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n814), .B1(new_n813), .B2(new_n804), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n784), .A2(KEYINPUT112), .A3(new_n782), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n816), .A2(new_n807), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n784), .A2(new_n782), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT112), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n806), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n811), .B1(new_n815), .B2(new_n821), .ZN(new_n822));
  OAI221_X1 g636(.A(new_n309), .B1(new_n630), .B2(new_n790), .C1(new_n798), .C2(new_n739), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n794), .A2(new_n312), .A3(new_n709), .A4(new_n789), .ZN(new_n827));
  XOR2_X1   g641(.A(new_n827), .B(KEYINPUT48), .Z(new_n828));
  NOR3_X1   g642(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n810), .A2(new_n822), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n832));
  INV_X1    g646(.A(new_n664), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n652), .A2(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n687), .A2(new_n834), .A3(new_n618), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n835), .B(new_n606), .C1(new_n681), .C2(new_n682), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n836), .A2(new_n707), .A3(KEYINPUT52), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n837), .A2(new_n672), .A3(KEYINPUT111), .A4(new_n740), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT98), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n635), .A2(new_n833), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n840), .B1(new_n841), .B2(new_n618), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n606), .B1(new_n842), .B2(new_n668), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n652), .B1(new_n706), .B2(new_n682), .ZN(new_n844));
  OAI22_X1  g658(.A1(new_n843), .A2(new_n844), .B1(new_n739), .B2(new_n738), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n836), .A2(new_n707), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n839), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT111), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n836), .A2(new_n707), .A3(KEYINPUT52), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n848), .B1(new_n845), .B2(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n838), .A2(new_n847), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n410), .B1(new_n630), .B2(new_n635), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n611), .A2(new_n556), .A3(new_n852), .A4(new_n606), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n717), .A2(new_n720), .A3(new_n725), .A4(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n607), .A2(new_n733), .A3(new_n653), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n606), .A2(new_n747), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n525), .A2(new_n438), .A3(new_n833), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n652), .B(new_n857), .C1(new_n706), .C2(new_n682), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n856), .B1(new_n858), .B2(new_n738), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n854), .A2(new_n855), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n752), .B1(new_n745), .B2(new_n749), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n832), .B1(new_n851), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n752), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT42), .B1(new_n744), .B2(new_n736), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n748), .A2(new_n746), .A3(new_n699), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n607), .A2(new_n733), .A3(new_n653), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n725), .A2(new_n853), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n709), .B(new_n716), .C1(new_n631), .C2(new_n636), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n858), .A2(new_n738), .ZN(new_n871));
  INV_X1    g685(.A(new_n856), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n868), .A2(new_n869), .A3(new_n870), .A4(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n837), .A2(new_n672), .A3(new_n740), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n847), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n875), .A2(KEYINPUT53), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n831), .B1(new_n863), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(KEYINPUT53), .B1(new_n851), .B2(new_n862), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n875), .A2(new_n832), .A3(new_n877), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT54), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n788), .B1(new_n830), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n598), .A2(new_n712), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n885), .A2(KEYINPUT49), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT109), .Z(new_n887));
  INV_X1    g701(.A(new_n525), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n555), .A2(new_n615), .A3(new_n558), .ZN(new_n889));
  AND4_X1   g703(.A1(new_n888), .A2(new_n686), .A3(new_n629), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n885), .A2(KEYINPUT49), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n887), .A2(new_n890), .A3(new_n683), .A4(new_n891), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT110), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n787), .B1(new_n884), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n893), .ZN(new_n895));
  AND4_X1   g709(.A1(new_n883), .A2(new_n822), .A3(new_n810), .A4(new_n829), .ZN(new_n896));
  OAI211_X1 g710(.A(KEYINPUT116), .B(new_n895), .C1(new_n896), .C2(new_n788), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n894), .A2(new_n897), .ZN(G75));
  NAND2_X1  g712(.A1(new_n880), .A2(new_n881), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n899), .A2(new_n381), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT56), .B1(new_n900), .B2(G210), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n360), .A2(new_n379), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n377), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT55), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n308), .A2(G952), .ZN(new_n906));
  NOR2_X1   g720(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n907));
  AND2_X1   g721(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n904), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n909), .B1(new_n900), .B2(new_n403), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n905), .A2(new_n906), .A3(new_n910), .ZN(G51));
  NAND3_X1  g725(.A1(new_n838), .A2(new_n847), .A3(new_n850), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n832), .B1(new_n875), .B2(new_n912), .ZN(new_n913));
  AND4_X1   g727(.A1(new_n832), .A2(new_n877), .A3(new_n861), .A4(new_n860), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n831), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT118), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g731(.A(KEYINPUT118), .B(new_n831), .C1(new_n913), .C2(new_n914), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n880), .A2(new_n881), .A3(KEYINPUT54), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n764), .B(KEYINPUT57), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n922), .B1(new_n578), .B2(new_n587), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n900), .A2(new_n768), .A3(new_n769), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n906), .B1(new_n923), .B2(new_n924), .ZN(G54));
  NAND2_X1  g739(.A1(KEYINPUT58), .A2(G475), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n880), .A2(new_n881), .A3(G902), .A4(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n519), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT119), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n928), .A2(new_n929), .ZN(new_n933));
  INV_X1    g747(.A(new_n906), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n928), .A2(KEYINPUT119), .A3(new_n929), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n932), .A2(new_n933), .A3(new_n934), .A4(new_n935), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT120), .Z(G60));
  NAND2_X1  g751(.A1(G478), .A2(G902), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT59), .Z(new_n939));
  AOI21_X1  g753(.A(KEYINPUT53), .B1(new_n875), .B2(new_n912), .ZN(new_n940));
  AND4_X1   g754(.A1(KEYINPUT53), .A2(new_n877), .A3(new_n861), .A4(new_n860), .ZN(new_n941));
  OAI21_X1  g755(.A(KEYINPUT54), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n939), .B1(new_n942), .B2(new_n915), .ZN(new_n943));
  OAI21_X1  g757(.A(KEYINPUT121), .B1(new_n943), .B2(new_n627), .ZN(new_n944));
  INV_X1    g758(.A(new_n939), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(new_n879), .B2(new_n882), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT121), .ZN(new_n947));
  INV_X1    g761(.A(new_n627), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n939), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n918), .A2(new_n919), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT118), .B1(new_n899), .B2(new_n831), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n944), .A2(new_n949), .A3(new_n934), .A4(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT122), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n906), .B1(new_n920), .B2(new_n950), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n957), .A2(KEYINPUT122), .A3(new_n944), .A4(new_n949), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n956), .A2(new_n958), .ZN(G63));
  NAND2_X1  g773(.A1(G217), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT60), .Z(new_n961));
  NAND3_X1  g775(.A1(new_n880), .A2(new_n881), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n906), .B1(new_n962), .B2(new_n553), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n649), .B(KEYINPUT123), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n963), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT61), .Z(G66));
  INV_X1    g780(.A(new_n315), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n308), .B1(new_n967), .B2(new_n370), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n854), .A2(new_n855), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n968), .B1(new_n970), .B2(new_n308), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n902), .B1(G898), .B2(new_n308), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT124), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT125), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n971), .B(new_n974), .ZN(G69));
  NOR2_X1   g789(.A1(new_n777), .A2(new_n785), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n709), .A2(new_n618), .A3(new_n687), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n776), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n672), .A2(new_n740), .A3(new_n707), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n978), .A2(new_n867), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n976), .A2(new_n308), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(new_n662), .B2(new_n308), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n297), .A2(new_n265), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT126), .Z(new_n984));
  NAND2_X1  g798(.A1(new_n505), .A2(new_n506), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n984), .B(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n982), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(G227), .A2(G900), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(G953), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n987), .A2(G953), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n630), .A2(new_n635), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n709), .A2(new_n747), .A3(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n976), .B1(new_n692), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n979), .A2(new_n695), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT62), .Z(new_n996));
  OAI21_X1  g810(.A(new_n991), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  AND3_X1   g811(.A1(new_n988), .A2(new_n990), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n990), .B1(new_n988), .B2(new_n997), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n998), .A2(new_n999), .ZN(G72));
  NOR3_X1   g814(.A1(new_n994), .A2(new_n970), .A3(new_n996), .ZN(new_n1001));
  NAND2_X1  g815(.A1(G472), .A2(G902), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT63), .Z(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n257), .B(new_n702), .C1(new_n1001), .C2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n976), .A2(new_n980), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1003), .B1(new_n1006), .B2(new_n970), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n286), .A2(new_n676), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT127), .Z(new_n1009));
  NAND2_X1  g823(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n300), .B1(new_n257), .B2(new_n286), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n1003), .B(new_n1011), .C1(new_n940), .C2(new_n941), .ZN(new_n1012));
  AND4_X1   g826(.A1(new_n934), .A2(new_n1005), .A3(new_n1010), .A4(new_n1012), .ZN(G57));
endmodule


