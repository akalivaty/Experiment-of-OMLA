//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT74), .A3(G128), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G119), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  XOR2_X1   g009(.A(KEYINPUT24), .B(G110), .Z(new_n196));
  INV_X1    g010(.A(KEYINPUT75), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT74), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n198), .B1(new_n193), .B2(G119), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n195), .A2(new_n196), .A3(new_n197), .A4(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n194), .A3(new_n192), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT24), .B(G110), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT75), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(KEYINPUT23), .B1(new_n193), .B2(G119), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n193), .A2(G119), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n193), .A2(KEYINPUT23), .A3(G119), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AOI22_X1  g022(.A1(new_n200), .A2(new_n203), .B1(G110), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  OR2_X1    g024(.A1(KEYINPUT16), .A2(G140), .ZN(new_n211));
  INV_X1    g025(.A(G125), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT76), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT76), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G125), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n211), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(G125), .A2(G140), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT76), .B(G125), .ZN(new_n219));
  INV_X1    g033(.A(G140), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI211_X1 g035(.A(new_n210), .B(new_n216), .C1(new_n221), .C2(KEYINPUT16), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n220), .B1(new_n213), .B2(new_n215), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT16), .B1(new_n223), .B2(new_n217), .ZN(new_n224));
  INV_X1    g038(.A(new_n216), .ZN(new_n225));
  AOI21_X1  g039(.A(G146), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n209), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n212), .A2(new_n220), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n210), .B1(new_n228), .B2(new_n217), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT77), .B(G110), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n206), .A2(new_n207), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n201), .A2(new_n202), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n230), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n224), .A2(G146), .A3(new_n225), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n227), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT22), .B(G137), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT78), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n238), .B(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G953), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT67), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G953), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G221), .ZN(new_n246));
  INV_X1    g060(.A(G234), .ZN(new_n247));
  NOR3_X1   g061(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n240), .B(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n237), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n227), .A2(new_n249), .A3(new_n236), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(new_n188), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT25), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n251), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n252), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n190), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n227), .A2(new_n236), .A3(new_n249), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n249), .B1(new_n227), .B2(new_n236), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n189), .A2(G902), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n257), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT70), .B(KEYINPUT32), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n191), .A2(G116), .ZN(new_n265));
  INV_X1    g079(.A(G116), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G119), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  XOR2_X1   g082(.A(KEYINPUT2), .B(G113), .Z(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n265), .A2(new_n267), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT2), .B(G113), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G143), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT1), .B1(new_n275), .B2(G146), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(G146), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n210), .A2(G143), .ZN(new_n278));
  OAI211_X1 g092(.A(G128), .B(new_n276), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n210), .A2(G143), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n275), .A2(G146), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n280), .B(new_n281), .C1(KEYINPUT1), .C2(new_n193), .ZN(new_n282));
  INV_X1    g096(.A(G134), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(G137), .ZN(new_n284));
  INV_X1    g098(.A(G137), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(G134), .ZN(new_n286));
  OAI21_X1  g100(.A(G131), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n279), .A2(new_n282), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n285), .A2(KEYINPUT11), .A3(G134), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n283), .A2(G137), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT65), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT64), .B(G131), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT11), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n294), .B1(new_n283), .B2(G137), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n291), .A2(new_n292), .A3(new_n293), .A4(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n289), .A3(new_n290), .ZN(new_n297));
  XOR2_X1   g111(.A(KEYINPUT64), .B(G131), .Z(new_n298));
  OAI21_X1  g112(.A(KEYINPUT65), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n288), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n295), .A2(new_n289), .A3(new_n290), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n292), .B1(new_n301), .B2(new_n293), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n297), .A2(new_n298), .A3(KEYINPUT65), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT66), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n297), .A2(new_n304), .A3(G131), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n304), .B1(new_n297), .B2(G131), .ZN(new_n306));
  OAI22_X1  g120(.A1(new_n302), .A2(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AND2_X1   g121(.A1(KEYINPUT0), .A2(G128), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n280), .A2(new_n281), .A3(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(G143), .B(G146), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT0), .B(G128), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n300), .B1(new_n307), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT30), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G131), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT66), .B1(new_n301), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n297), .A2(new_n304), .A3(G131), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n296), .A2(new_n299), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n312), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NOR3_X1   g136(.A1(new_n322), .A2(KEYINPUT30), .A3(new_n300), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n274), .B1(new_n316), .B2(new_n323), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n279), .A2(new_n282), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n321), .A2(new_n325), .A3(new_n287), .ZN(new_n326));
  INV_X1    g140(.A(new_n274), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n318), .A2(new_n319), .B1(new_n296), .B2(new_n299), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n326), .B(new_n327), .C1(new_n328), .C2(new_n312), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT67), .B(G953), .ZN(new_n330));
  INV_X1    g144(.A(G237), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(G210), .A3(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(KEYINPUT27), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT26), .B(G101), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n333), .B(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT68), .B(KEYINPUT31), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n324), .A2(new_n329), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n335), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n274), .B1(new_n322), .B2(new_n300), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n340), .B1(new_n341), .B2(new_n329), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT28), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n329), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n338), .B1(new_n342), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT30), .B1(new_n322), .B2(new_n300), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n326), .B(new_n315), .C1(new_n328), .C2(new_n312), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n327), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NOR3_X1   g163(.A1(new_n322), .A2(new_n274), .A3(new_n300), .ZN(new_n350));
  NOR3_X1   g164(.A1(new_n349), .A2(new_n350), .A3(new_n338), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT31), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n337), .B(new_n346), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(G472), .A2(G902), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n264), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n353), .A2(new_n354), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n355), .B1(KEYINPUT32), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n344), .B(KEYINPUT73), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n335), .A2(KEYINPUT29), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT71), .B1(new_n341), .B2(new_n329), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT71), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n361), .B1(new_n314), .B2(new_n327), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT28), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT72), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT72), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n365), .B(KEYINPUT28), .C1(new_n360), .C2(new_n362), .ZN(new_n366));
  AOI211_X1 g180(.A(new_n358), .B(new_n359), .C1(new_n364), .C2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n314), .A2(new_n327), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n339), .B1(new_n368), .B2(new_n350), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(new_n344), .A3(new_n335), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n338), .B1(new_n349), .B2(new_n350), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n188), .ZN(new_n374));
  OAI21_X1  g188(.A(G472), .B1(new_n367), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n263), .B1(new_n357), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(G210), .B1(G237), .B2(G902), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n279), .A2(new_n282), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n219), .ZN(new_n380));
  INV_X1    g194(.A(new_n219), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n312), .A2(KEYINPUT81), .A3(new_n381), .ZN(new_n382));
  AND2_X1   g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n312), .A2(new_n381), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT81), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G224), .ZN(new_n387));
  OAI21_X1  g201(.A(KEYINPUT7), .B1(new_n387), .B2(G953), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n383), .A2(KEYINPUT83), .A3(new_n386), .A4(new_n389), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n386), .A2(new_n380), .A3(new_n382), .A4(new_n389), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT83), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n384), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n381), .B1(new_n279), .B2(new_n282), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n388), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G104), .ZN(new_n398));
  OAI21_X1  g212(.A(KEYINPUT3), .B1(new_n398), .B2(G107), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT3), .ZN(new_n400));
  INV_X1    g214(.A(G107), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(new_n401), .A3(G104), .ZN(new_n402));
  INV_X1    g216(.A(G101), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n398), .A2(G107), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n399), .A2(new_n402), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n398), .A2(G107), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n401), .A2(G104), .ZN(new_n407));
  OAI21_X1  g221(.A(G101), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(G113), .B1(new_n265), .B2(KEYINPUT5), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT82), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI211_X1 g226(.A(KEYINPUT82), .B(G113), .C1(new_n265), .C2(KEYINPUT5), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT5), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n412), .B(new_n413), .C1(new_n414), .C2(new_n271), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n409), .B1(new_n415), .B2(new_n270), .ZN(new_n416));
  XNOR2_X1  g230(.A(G110), .B(G122), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n417), .B(KEYINPUT8), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n271), .A2(new_n414), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n270), .B1(new_n419), .B2(new_n410), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n405), .A2(new_n408), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n418), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n397), .B1(new_n416), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT84), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n394), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n399), .A2(new_n402), .A3(new_n404), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G101), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(KEYINPUT4), .A3(new_n405), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT4), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n427), .A2(new_n430), .A3(G101), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n429), .A2(new_n274), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT80), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT80), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n429), .A2(new_n434), .A3(new_n274), .A4(new_n431), .ZN(new_n435));
  OR2_X1    g249(.A1(new_n420), .A2(new_n409), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n433), .A2(new_n417), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n426), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n423), .B1(new_n390), .B2(new_n393), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n439), .A2(new_n425), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n188), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n433), .A2(new_n435), .A3(new_n436), .ZN(new_n442));
  INV_X1    g256(.A(new_n417), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(KEYINPUT6), .A3(new_n437), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT6), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n442), .A2(new_n446), .A3(new_n443), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n383), .A2(new_n386), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n387), .A2(G953), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n448), .B(new_n449), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n445), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n378), .B1(new_n441), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n437), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(new_n439), .B2(new_n425), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n394), .A2(new_n424), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT84), .ZN(new_n456));
  AOI21_X1  g270(.A(G902), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n445), .A2(new_n447), .A3(new_n450), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n458), .A3(new_n377), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n452), .A2(KEYINPUT85), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT85), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n457), .A2(new_n461), .A3(new_n458), .A4(new_n377), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n241), .A2(G952), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n463), .B1(G234), .B2(G237), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n245), .B(G902), .C1(new_n247), .C2(new_n331), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(KEYINPUT96), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(G898), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(G214), .B1(G237), .B2(G902), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n460), .A2(new_n462), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n242), .A2(new_n244), .A3(G214), .A4(new_n331), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n275), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n330), .A2(G143), .A3(G214), .A4(new_n331), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n298), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT88), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n474), .A2(new_n475), .A3(new_n293), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT17), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT88), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n476), .A2(new_n481), .A3(new_n298), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n478), .A2(new_n479), .A3(new_n480), .A4(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n222), .A2(new_n226), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n481), .B1(new_n476), .B2(new_n298), .ZN(new_n485));
  AOI211_X1 g299(.A(KEYINPUT88), .B(new_n293), .C1(new_n474), .C2(new_n475), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT17), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n483), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(G113), .B(G122), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(new_n398), .ZN(new_n490));
  NAND2_X1  g304(.A1(KEYINPUT18), .A2(G131), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n476), .B(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n223), .A2(new_n217), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT86), .ZN(new_n494));
  AOI22_X1  g308(.A1(new_n493), .A2(G146), .B1(new_n494), .B2(new_n229), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n221), .A2(KEYINPUT86), .A3(new_n210), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT87), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  OAI22_X1  g312(.A1(new_n230), .A2(KEYINPUT86), .B1(new_n221), .B2(new_n210), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n493), .A2(new_n494), .A3(G146), .ZN(new_n500));
  AOI21_X1  g314(.A(KEYINPUT87), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n492), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n488), .A2(new_n490), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT90), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n488), .A2(KEYINPUT90), .A3(new_n502), .A4(new_n490), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n478), .A2(new_n482), .A3(new_n479), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT89), .ZN(new_n509));
  OR2_X1    g323(.A1(new_n509), .A2(KEYINPUT19), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(KEYINPUT19), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n510), .B(new_n511), .C1(new_n228), .C2(new_n217), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n513), .B1(KEYINPUT19), .B2(new_n493), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n222), .B1(new_n210), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n508), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n502), .ZN(new_n517));
  INV_X1    g331(.A(new_n490), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n507), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT20), .ZN(new_n521));
  NOR2_X1   g335(.A1(G475), .A2(G902), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n505), .A2(new_n506), .B1(new_n518), .B2(new_n517), .ZN(new_n524));
  INV_X1    g338(.A(new_n522), .ZN(new_n525));
  OAI21_X1  g339(.A(KEYINPUT20), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n490), .B1(new_n488), .B2(new_n502), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n528), .B1(new_n505), .B2(new_n506), .ZN(new_n529));
  OAI21_X1  g343(.A(G475), .B1(new_n529), .B2(G902), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n275), .A2(KEYINPUT13), .A3(G128), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n193), .A2(G143), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n275), .A2(G128), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT13), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n531), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n536), .A2(G134), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n533), .A2(new_n532), .A3(new_n283), .ZN(new_n538));
  INV_X1    g352(.A(G122), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(G116), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n266), .A2(G122), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n541), .A3(new_n401), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n401), .B1(new_n540), .B2(new_n541), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n538), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n537), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT93), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT14), .B1(new_n539), .B2(G116), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT92), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT92), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n541), .A2(new_n550), .A3(KEYINPUT14), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT14), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(new_n266), .A3(G122), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n549), .A2(new_n551), .A3(new_n540), .A4(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n547), .B1(new_n554), .B2(G107), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n542), .A2(KEYINPUT91), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT91), .ZN(new_n557));
  XNOR2_X1  g371(.A(G116), .B(G122), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n557), .B1(new_n558), .B2(new_n401), .ZN(new_n559));
  INV_X1    g373(.A(new_n538), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n283), .B1(new_n533), .B2(new_n532), .ZN(new_n561));
  OAI22_X1  g375(.A1(new_n556), .A2(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n554), .A2(new_n547), .A3(G107), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n546), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT9), .B(G234), .ZN(new_n566));
  NOR3_X1   g380(.A1(new_n566), .A2(new_n187), .A3(G953), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT95), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n554), .A2(G107), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT93), .ZN(new_n570));
  OR2_X1    g384(.A1(new_n560), .A2(new_n561), .ZN(new_n571));
  OR2_X1    g385(.A1(new_n556), .A2(new_n559), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n570), .A2(new_n564), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n546), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT95), .ZN(new_n576));
  INV_X1    g390(.A(new_n567), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(KEYINPUT94), .B1(new_n565), .B2(new_n567), .ZN(new_n579));
  AND4_X1   g393(.A1(KEYINPUT94), .A2(new_n573), .A3(new_n574), .A4(new_n567), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n568), .B(new_n578), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n188), .ZN(new_n582));
  INV_X1    g396(.A(G478), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(KEYINPUT15), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n582), .B(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n527), .A2(new_n530), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n330), .A2(G227), .ZN(new_n588));
  XOR2_X1   g402(.A(G110), .B(G140), .Z(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n279), .A2(new_n405), .A3(new_n408), .A4(new_n282), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(KEYINPUT10), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n429), .A2(new_n313), .A3(new_n431), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n328), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT10), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n325), .A2(new_n421), .A3(KEYINPUT10), .ZN(new_n597));
  AND4_X1   g411(.A1(new_n328), .A2(new_n593), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n590), .B1(new_n594), .B2(new_n598), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n328), .A2(new_n593), .A3(new_n596), .A4(new_n597), .ZN(new_n600));
  INV_X1    g414(.A(new_n590), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n379), .A2(new_n409), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n591), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n307), .A2(KEYINPUT12), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT12), .B1(new_n307), .B2(new_n603), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n600), .B(new_n601), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n599), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(G469), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(new_n608), .A3(new_n188), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT79), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n610), .B1(new_n598), .B2(new_n590), .ZN(new_n611));
  INV_X1    g425(.A(new_n594), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n600), .A2(KEYINPUT79), .A3(new_n601), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n600), .B1(new_n604), .B2(new_n605), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n590), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(G469), .A3(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n608), .A2(new_n188), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n609), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n566), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n246), .B1(new_n621), .B2(new_n188), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n587), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n376), .A2(new_n472), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT97), .B(G101), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G3));
  INV_X1    g442(.A(G472), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n353), .B2(new_n188), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n356), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n632), .A2(new_n263), .A3(new_n624), .ZN(new_n633));
  OR2_X1    g447(.A1(new_n529), .A2(G902), .ZN(new_n634));
  AOI22_X1  g448(.A1(new_n526), .A2(new_n523), .B1(new_n634), .B2(G475), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n441), .A2(new_n451), .A3(new_n378), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n377), .B1(new_n457), .B2(new_n458), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n469), .B(new_n470), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n582), .A2(new_n583), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n575), .A2(new_n577), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n565), .A2(new_n567), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT33), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n579), .A2(new_n580), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n568), .A2(new_n578), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT98), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n581), .A2(KEYINPUT98), .A3(new_n643), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n644), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n583), .A2(G902), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n640), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n635), .A2(new_n638), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n633), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT34), .B(G104), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT99), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n655), .B(new_n657), .ZN(G6));
  XNOR2_X1  g472(.A(new_n582), .B(new_n584), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n521), .B1(new_n520), .B2(new_n522), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n524), .A2(KEYINPUT20), .A3(new_n525), .ZN(new_n661));
  OAI211_X1 g475(.A(new_n530), .B(new_n659), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n638), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n633), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n664), .B(KEYINPUT100), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT101), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT35), .B(G107), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  AOI21_X1  g482(.A(KEYINPUT25), .B1(new_n260), .B2(new_n188), .ZN(new_n669));
  INV_X1    g483(.A(new_n256), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n189), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT36), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n249), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(new_n237), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n261), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n671), .A2(new_n672), .A3(new_n676), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n675), .A2(new_n261), .ZN(new_n678));
  OAI21_X1  g492(.A(KEYINPUT102), .B1(new_n257), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n625), .A2(new_n472), .A3(new_n631), .A4(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT37), .B(G110), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G12));
  AOI22_X1  g497(.A1(new_n357), .A2(new_n375), .B1(new_n679), .B2(new_n677), .ZN(new_n684));
  INV_X1    g498(.A(G900), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n466), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(new_n464), .ZN(new_n687));
  OAI21_X1  g501(.A(KEYINPUT103), .B1(new_n662), .B2(new_n687), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n659), .A2(new_n530), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT103), .ZN(new_n690));
  INV_X1    g504(.A(new_n687), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n689), .A2(new_n690), .A3(new_n527), .A4(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n470), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n452), .B2(new_n459), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n623), .A3(new_n620), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n684), .A2(new_n688), .A3(new_n692), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G128), .ZN(G30));
  XOR2_X1   g512(.A(new_n687), .B(KEYINPUT39), .Z(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n624), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n702), .A2(KEYINPUT40), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(KEYINPUT40), .ZN(new_n704));
  NOR4_X1   g518(.A1(new_n703), .A2(new_n704), .A3(new_n693), .A4(new_n680), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n460), .A2(new_n462), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT38), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n353), .A2(new_n354), .ZN(new_n709));
  INV_X1    g523(.A(new_n264), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n353), .A2(KEYINPUT32), .A3(new_n354), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n360), .A2(new_n362), .ZN(new_n714));
  AOI21_X1  g528(.A(G902), .B1(new_n714), .B2(new_n338), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n324), .A2(new_n329), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n335), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n629), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n713), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n635), .A2(new_n586), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n705), .A2(new_n708), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G143), .ZN(G45));
  NOR3_X1   g536(.A1(new_n635), .A2(new_n653), .A3(new_n687), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n684), .A2(new_n723), .A3(new_n696), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G146), .ZN(G48));
  INV_X1    g539(.A(new_n609), .ZN(new_n726));
  AOI21_X1  g540(.A(G902), .B1(new_n599), .B2(new_n606), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n608), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n726), .A2(new_n728), .A3(new_n622), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n654), .A2(new_n376), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT41), .B(G113), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G15));
  NAND3_X1  g546(.A1(new_n376), .A2(new_n663), .A3(new_n729), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G116), .ZN(G18));
  INV_X1    g548(.A(new_n587), .ZN(new_n735));
  INV_X1    g549(.A(new_n729), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n638), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n358), .B1(new_n364), .B2(new_n366), .ZN(new_n738));
  INV_X1    g552(.A(new_n359), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n374), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n712), .B(new_n711), .C1(new_n740), .C2(new_n629), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n735), .A2(new_n737), .A3(new_n741), .A4(new_n680), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  OAI21_X1  g557(.A(KEYINPUT31), .B1(new_n716), .B2(new_n338), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n744), .B(new_n337), .C1(new_n738), .C2(new_n335), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n630), .B1(new_n745), .B2(new_n354), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n720), .A2(new_n746), .A3(new_n737), .A4(new_n262), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G122), .ZN(G24));
  INV_X1    g562(.A(new_n630), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n744), .A2(new_n337), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n364), .A2(new_n366), .ZN(new_n751));
  INV_X1    g565(.A(new_n358), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n750), .B1(new_n753), .B2(new_n338), .ZN(new_n754));
  INV_X1    g568(.A(new_n354), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n749), .B(new_n680), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n530), .B1(new_n660), .B2(new_n661), .ZN(new_n757));
  INV_X1    g571(.A(new_n644), .ZN(new_n758));
  INV_X1    g572(.A(new_n650), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT98), .B1(new_n581), .B2(new_n643), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n758), .B(new_n652), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n639), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n757), .A2(new_n762), .A3(new_n691), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n756), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n694), .A2(new_n729), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G125), .ZN(G27));
  INV_X1    g582(.A(KEYINPUT32), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n709), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n712), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n738), .A2(new_n739), .ZN(new_n772));
  INV_X1    g586(.A(new_n374), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n629), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n262), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT105), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n375), .A2(new_n712), .A3(new_n770), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT105), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n778), .A3(new_n262), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n693), .B1(new_n460), .B2(new_n462), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n618), .B1(new_n727), .B2(new_n608), .ZN(new_n782));
  AOI211_X1 g596(.A(KEYINPUT104), .B(new_n622), .C1(new_n782), .C2(new_n617), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT104), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n784), .B1(new_n620), .B2(new_n623), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n781), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n757), .A2(new_n762), .A3(KEYINPUT42), .A4(new_n691), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n786), .A2(new_n706), .A3(new_n470), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n790), .A2(new_n376), .A3(new_n723), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT42), .ZN(new_n792));
  AOI22_X1  g606(.A1(new_n780), .A2(new_n789), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(new_n317), .ZN(G33));
  AND2_X1   g608(.A1(new_n688), .A2(new_n692), .ZN(new_n795));
  AND4_X1   g609(.A1(new_n741), .A2(new_n262), .A3(new_n781), .A4(new_n786), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G134), .ZN(G36));
  INV_X1    g612(.A(KEYINPUT43), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n799), .B1(new_n757), .B2(KEYINPUT106), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n757), .A2(new_n653), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n632), .A3(new_n680), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT44), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT45), .B1(new_n614), .B2(new_n616), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n608), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n614), .A2(KEYINPUT45), .A3(new_n616), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(new_n618), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n811), .A2(KEYINPUT46), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n609), .B1(new_n811), .B2(KEYINPUT46), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n623), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OR2_X1    g628(.A1(new_n814), .A2(new_n700), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n805), .A2(new_n781), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n803), .A2(new_n804), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(new_n285), .ZN(G39));
  INV_X1    g634(.A(KEYINPUT47), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n814), .A2(new_n821), .ZN(new_n822));
  OAI211_X1 g636(.A(KEYINPUT47), .B(new_n623), .C1(new_n812), .C2(new_n813), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n781), .ZN(new_n825));
  NOR4_X1   g639(.A1(new_n825), .A2(new_n763), .A3(new_n741), .A4(new_n262), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G140), .ZN(G42));
  NAND3_X1  g642(.A1(new_n262), .A2(new_n470), .A3(new_n623), .ZN(new_n829));
  XOR2_X1   g643(.A(new_n829), .B(KEYINPUT107), .Z(new_n830));
  NOR2_X1   g644(.A1(new_n726), .A2(new_n728), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT49), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR4_X1   g647(.A1(new_n830), .A2(new_n757), .A3(new_n653), .A4(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT108), .ZN(new_n835));
  INV_X1    g649(.A(new_n708), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n719), .B1(new_n832), .B2(new_n831), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n719), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n825), .A2(new_n736), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n839), .A2(new_n840), .A3(new_n262), .A4(new_n464), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n635), .A2(new_n653), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  OAI211_X1 g657(.A(G952), .B(new_n241), .C1(new_n841), .C2(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n802), .A2(new_n464), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n746), .A2(new_n262), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n844), .B1(new_n847), .B2(new_n766), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT48), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n845), .A2(new_n840), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n849), .B1(new_n850), .B2(new_n780), .ZN(new_n851));
  AND4_X1   g665(.A1(new_n849), .A2(new_n845), .A3(new_n780), .A4(new_n840), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n848), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n708), .A2(new_n470), .A3(new_n736), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n854), .A2(new_n802), .A3(new_n464), .A4(new_n846), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT117), .B1(new_n855), .B2(KEYINPUT116), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT50), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n831), .A2(new_n622), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n822), .A2(new_n823), .A3(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n860), .A2(new_n845), .A3(new_n846), .A4(new_n781), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT116), .B1(KEYINPUT117), .B2(KEYINPUT50), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n855), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n756), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n845), .A2(new_n865), .A3(new_n840), .ZN(new_n866));
  OR3_X1    g680(.A1(new_n841), .A2(new_n757), .A3(new_n762), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n861), .A2(new_n864), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n858), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT51), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n853), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n858), .A2(new_n868), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT118), .B1(new_n872), .B2(KEYINPUT51), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n874));
  NOR4_X1   g688(.A1(new_n858), .A2(new_n868), .A3(new_n874), .A4(new_n870), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n871), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(KEYINPUT119), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n871), .B(new_n878), .C1(new_n873), .C2(new_n875), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n775), .A2(KEYINPUT105), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n778), .B1(new_n777), .B2(new_n262), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n789), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n791), .A2(new_n792), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AND4_X1   g698(.A1(new_n730), .A2(new_n733), .A3(new_n742), .A4(new_n747), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR4_X1   g700(.A1(new_n624), .A2(new_n257), .A3(new_n678), .A4(new_n687), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n719), .A2(new_n887), .A3(new_n694), .A4(new_n720), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n767), .A2(new_n697), .A3(new_n888), .A4(new_n724), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT52), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n886), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT109), .ZN(new_n894));
  OR3_X1    g708(.A1(new_n471), .A2(new_n662), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n894), .B1(new_n471), .B2(new_n662), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n895), .A2(new_n633), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n633), .A2(new_n472), .A3(new_n842), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n897), .A2(new_n626), .A3(new_n898), .A4(new_n681), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT111), .ZN(new_n900));
  AOI211_X1 g714(.A(new_n622), .B(new_n687), .C1(new_n782), .C2(new_n617), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n680), .A2(new_n901), .A3(new_n586), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n741), .A2(new_n902), .A3(new_n635), .A4(new_n781), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT110), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n680), .A2(new_n901), .A3(new_n586), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(new_n757), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT110), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n906), .A2(new_n907), .A3(new_n741), .A4(new_n781), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n865), .A2(new_n723), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n688), .A2(new_n692), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n741), .A2(new_n262), .A3(new_n781), .A4(new_n786), .ZN(new_n912));
  OAI22_X1  g726(.A1(new_n910), .A2(new_n787), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n900), .B1(new_n909), .B2(new_n913), .ZN(new_n914));
  AOI22_X1  g728(.A1(new_n795), .A2(new_n796), .B1(new_n764), .B2(new_n790), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n904), .A2(new_n908), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n915), .A2(KEYINPUT111), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n899), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n893), .A2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT53), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n889), .B(KEYINPUT52), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n920), .B1(new_n921), .B2(KEYINPUT112), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n919), .B(new_n922), .Z(new_n923));
  AOI21_X1  g737(.A(KEYINPUT53), .B1(new_n893), .B2(new_n918), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT113), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n914), .A2(new_n917), .ZN(new_n926));
  INV_X1    g740(.A(new_n899), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI211_X1 g742(.A(KEYINPUT113), .B(new_n899), .C1(new_n914), .C2(new_n917), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT114), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n730), .A2(new_n733), .A3(new_n742), .A4(new_n747), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n931), .B1(new_n793), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n884), .A2(new_n885), .A3(KEYINPUT114), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n933), .A2(new_n934), .A3(KEYINPUT53), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n935), .A2(new_n921), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n924), .B1(new_n930), .B2(new_n936), .ZN(new_n937));
  XOR2_X1   g751(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n938));
  AOI22_X1  g752(.A1(new_n923), .A2(KEYINPUT54), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n877), .A2(new_n879), .A3(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(G952), .A2(G953), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n838), .B1(new_n940), .B2(new_n941), .ZN(G75));
  INV_X1    g756(.A(KEYINPUT56), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n909), .A2(new_n913), .A3(new_n900), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT111), .B1(new_n915), .B2(new_n916), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n927), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT113), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n918), .A2(new_n925), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n936), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n919), .A2(new_n920), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(G902), .ZN(new_n952));
  INV_X1    g766(.A(G210), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n943), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n445), .A2(new_n447), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n955), .A2(new_n450), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n956), .A2(new_n451), .ZN(new_n957));
  XOR2_X1   g771(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n954), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n954), .A2(new_n960), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n330), .A2(G952), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(G51));
  INV_X1    g778(.A(new_n938), .ZN(new_n965));
  OAI21_X1  g779(.A(KEYINPUT121), .B1(new_n951), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n951), .A2(new_n965), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT121), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n949), .A2(new_n950), .A3(new_n968), .A4(new_n938), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n966), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n618), .B(KEYINPUT57), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n607), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n937), .A2(new_n188), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n974), .A2(KEYINPUT122), .A3(new_n810), .ZN(new_n975));
  AOI21_X1  g789(.A(KEYINPUT122), .B1(new_n974), .B2(new_n810), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n963), .B1(new_n973), .B2(new_n977), .ZN(G54));
  NAND3_X1  g792(.A1(new_n974), .A2(KEYINPUT58), .A3(G475), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n979), .A2(new_n524), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(new_n524), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n980), .A2(new_n981), .A3(new_n963), .ZN(G60));
  INV_X1    g796(.A(new_n651), .ZN(new_n983));
  NAND2_X1  g797(.A1(G478), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT59), .Z(new_n985));
  OAI21_X1  g799(.A(new_n983), .B1(new_n939), .B2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n963), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n983), .A2(new_n985), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n970), .A2(new_n988), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n986), .A2(new_n987), .A3(new_n989), .ZN(G63));
  XOR2_X1   g804(.A(new_n675), .B(KEYINPUT124), .Z(new_n991));
  INV_X1    g805(.A(KEYINPUT123), .ZN(new_n992));
  NAND2_X1  g806(.A1(G217), .A2(G902), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT60), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n992), .B1(new_n951), .B2(new_n995), .ZN(new_n996));
  AOI211_X1 g810(.A(KEYINPUT123), .B(new_n994), .C1(new_n949), .C2(new_n950), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n991), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(KEYINPUT123), .B1(new_n937), .B2(new_n994), .ZN(new_n999));
  INV_X1    g813(.A(new_n260), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n951), .A2(new_n992), .A3(new_n995), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n998), .A2(new_n1002), .A3(new_n987), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT61), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n998), .A2(new_n1002), .A3(KEYINPUT61), .A4(new_n987), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1005), .A2(new_n1006), .ZN(G66));
  OAI21_X1  g821(.A(G953), .B1(new_n467), .B2(new_n387), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n899), .A2(new_n932), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1008), .B1(new_n1009), .B2(new_n245), .ZN(new_n1010));
  INV_X1    g824(.A(G898), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n955), .B1(new_n1011), .B2(new_n245), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1010), .B(new_n1012), .Z(G69));
  AOI21_X1  g827(.A(new_n330), .B1(G227), .B2(G900), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n347), .A2(new_n348), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n1015), .B(new_n514), .Z(new_n1016));
  AND2_X1   g830(.A1(new_n697), .A2(new_n724), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n1017), .A2(new_n767), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(new_n721), .ZN(new_n1019));
  OR2_X1    g833(.A1(new_n1019), .A2(KEYINPUT62), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n843), .A2(new_n662), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n1021), .A2(new_n376), .A3(new_n701), .A4(new_n781), .ZN(new_n1022));
  AND2_X1   g836(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n827), .B1(new_n817), .B2(new_n818), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1019), .A2(KEYINPUT62), .ZN(new_n1026));
  AND3_X1   g840(.A1(new_n1023), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1016), .B1(new_n1027), .B2(new_n245), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1016), .B1(G900), .B2(new_n245), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n780), .A2(new_n694), .A3(new_n720), .ZN(new_n1030));
  OR2_X1    g844(.A1(new_n815), .A2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g845(.A1(new_n1031), .A2(new_n884), .A3(new_n1018), .A4(new_n797), .ZN(new_n1032));
  OR2_X1    g846(.A1(new_n1024), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1029), .B1(new_n1033), .B2(new_n245), .ZN(new_n1034));
  INV_X1    g848(.A(KEYINPUT126), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1028), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g851(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n1014), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  XOR2_X1   g853(.A(new_n1014), .B(KEYINPUT125), .Z(new_n1040));
  NAND3_X1  g854(.A1(new_n1028), .A2(new_n1034), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1039), .A2(new_n1041), .ZN(G72));
  NAND2_X1  g856(.A1(G472), .A2(G902), .ZN(new_n1043));
  XOR2_X1   g857(.A(new_n1043), .B(KEYINPUT63), .Z(new_n1044));
  XNOR2_X1  g858(.A(new_n716), .B(new_n338), .ZN(new_n1045));
  AND3_X1   g859(.A1(new_n923), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  NAND4_X1  g860(.A1(new_n1023), .A2(new_n1009), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n717), .B1(new_n1047), .B2(new_n1044), .ZN(new_n1048));
  INV_X1    g862(.A(new_n1009), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1044), .B1(new_n1033), .B2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g864(.A1(new_n716), .A2(new_n335), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n1052), .A2(new_n987), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1053), .A2(KEYINPUT127), .ZN(new_n1054));
  INV_X1    g868(.A(KEYINPUT127), .ZN(new_n1055));
  NAND3_X1  g869(.A1(new_n1052), .A2(new_n1055), .A3(new_n987), .ZN(new_n1056));
  AOI211_X1 g870(.A(new_n1046), .B(new_n1048), .C1(new_n1054), .C2(new_n1056), .ZN(G57));
endmodule


