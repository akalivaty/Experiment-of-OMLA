//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 1 1 0 0 0 1 0 1 0 0 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n850, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1032, new_n1033, new_n1034, new_n1035, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1043, new_n1044,
    new_n1045, new_n1046;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(KEYINPUT94), .B(G36gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT95), .ZN(new_n209));
  INV_X1    g008(.A(G29gat), .ZN(new_n210));
  OR3_X1    g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n209), .B1(new_n208), .B2(new_n210), .ZN(new_n212));
  NOR2_X1   g011(.A1(G29gat), .A2(G36gat), .ZN(new_n213));
  XOR2_X1   g012(.A(new_n213), .B(KEYINPUT14), .Z(new_n214));
  NAND3_X1  g013(.A1(new_n211), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT15), .ZN(new_n216));
  XNOR2_X1  g015(.A(G43gat), .B(G50gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT93), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(new_n218), .B2(new_n217), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT96), .ZN(new_n222));
  INV_X1    g021(.A(G50gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(G43gat), .ZN(new_n224));
  INV_X1    g023(.A(G43gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(KEYINPUT96), .A3(G50gat), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n224), .B(new_n226), .C1(new_n225), .C2(G50gat), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n227), .A2(new_n216), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n220), .B1(new_n215), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n221), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT17), .ZN(new_n231));
  XNOR2_X1  g030(.A(G15gat), .B(G22gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT16), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n232), .B1(new_n233), .B2(G1gat), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(G1gat), .B2(new_n232), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n235), .B(G8gat), .Z(new_n236));
  INV_X1    g035(.A(KEYINPUT17), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n237), .A3(new_n229), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n231), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G229gat), .A2(G233gat), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n221), .A2(new_n229), .ZN(new_n241));
  INV_X1    g040(.A(new_n236), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n239), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT18), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n236), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n240), .B(KEYINPUT13), .Z(new_n248));
  AOI22_X1  g047(.A1(new_n244), .A2(new_n245), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n239), .A2(KEYINPUT18), .A3(new_n240), .A4(new_n243), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n207), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n249), .A2(new_n207), .A3(new_n250), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G183gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT27), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT27), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(G183gat), .ZN(new_n259));
  INV_X1    g058(.A(G190gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT28), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT27), .B(G183gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n264), .A2(KEYINPUT28), .A3(new_n260), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(G169gat), .A2(G176gat), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(G169gat), .A2(G176gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT26), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n269), .A2(new_n272), .B1(G183gat), .B2(G190gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n266), .A2(new_n273), .ZN(new_n274));
  XOR2_X1   g073(.A(KEYINPUT65), .B(KEYINPUT25), .Z(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n270), .A2(KEYINPUT23), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(new_n268), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT23), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT66), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT66), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT23), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n270), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n278), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT24), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(G183gat), .A3(G190gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n256), .A2(G190gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n260), .A2(G183gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n287), .B1(new_n290), .B2(KEYINPUT24), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n276), .B1(new_n284), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G183gat), .B(G190gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n286), .B1(new_n293), .B2(new_n285), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT67), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n268), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n277), .A2(KEYINPUT25), .A3(new_n296), .A4(new_n297), .ZN(new_n298));
  NOR3_X1   g097(.A1(new_n294), .A2(new_n298), .A3(new_n283), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n274), .B1(new_n292), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT29), .ZN(new_n301));
  NAND2_X1  g100(.A1(G226gat), .A2(G233gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(KEYINPUT66), .B(KEYINPUT23), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n277), .B(new_n268), .C1(new_n304), .C2(new_n270), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n275), .B1(new_n305), .B2(new_n294), .ZN(new_n306));
  INV_X1    g105(.A(new_n298), .ZN(new_n307));
  INV_X1    g106(.A(new_n283), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n291), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT68), .ZN(new_n311));
  AND3_X1   g110(.A1(new_n266), .A2(new_n311), .A3(new_n273), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n311), .B1(new_n266), .B2(new_n273), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n310), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n303), .B1(new_n302), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT77), .ZN(new_n316));
  XNOR2_X1  g115(.A(G197gat), .B(G204gat), .ZN(new_n317));
  INV_X1    g116(.A(G211gat), .ZN(new_n318));
  OR2_X1    g117(.A1(KEYINPUT75), .A2(G218gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(KEYINPUT75), .A2(G218gat), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT22), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT74), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT74), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT22), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n317), .B1(new_n321), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n318), .A2(G218gat), .ZN(new_n328));
  INV_X1    g127(.A(G218gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n329), .A2(G211gat), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT76), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(G211gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n318), .A2(G218gat), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT76), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n327), .A2(new_n336), .ZN(new_n337));
  AND2_X1   g136(.A1(KEYINPUT75), .A2(G218gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(KEYINPUT75), .A2(G218gat), .ZN(new_n339));
  OAI21_X1  g138(.A(G211gat), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(KEYINPUT74), .B(KEYINPUT22), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n342), .A2(new_n317), .B1(new_n331), .B2(new_n335), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n316), .B1(new_n337), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n336), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n342), .A2(new_n317), .A3(new_n331), .A4(new_n335), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n346), .A3(KEYINPUT77), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n315), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT80), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT80), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n315), .A2(new_n351), .A3(new_n348), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G8gat), .B(G36gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(G64gat), .B(G92gat), .ZN(new_n355));
  XOR2_X1   g154(.A(new_n354), .B(new_n355), .Z(new_n356));
  AOI22_X1  g155(.A1(new_n306), .A2(new_n309), .B1(new_n266), .B2(new_n273), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT78), .B1(new_n357), .B2(new_n302), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT28), .B1(new_n264), .B2(new_n260), .ZN(new_n359));
  AND4_X1   g158(.A1(KEYINPUT28), .A2(new_n257), .A3(new_n259), .A4(new_n260), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n272), .A2(new_n268), .A3(new_n267), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n362), .B1(new_n256), .B2(new_n260), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT68), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n266), .A2(new_n311), .A3(new_n273), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT29), .B1(new_n366), .B2(new_n310), .ZN(new_n367));
  INV_X1    g166(.A(new_n302), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n358), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n364), .A2(new_n365), .B1(new_n309), .B2(new_n306), .ZN(new_n370));
  OAI211_X1 g169(.A(KEYINPUT78), .B(new_n302), .C1(new_n370), .C2(KEYINPUT29), .ZN(new_n371));
  AOI211_X1 g170(.A(KEYINPUT79), .B(new_n348), .C1(new_n369), .C2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT79), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n368), .B1(new_n314), .B2(new_n301), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n375), .B1(new_n300), .B2(new_n368), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n371), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n348), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n373), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n353), .B(new_n356), .C1(new_n372), .C2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT30), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n314), .A2(new_n301), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n376), .B1(new_n383), .B2(new_n302), .ZN(new_n384));
  AOI211_X1 g183(.A(new_n375), .B(new_n368), .C1(new_n314), .C2(new_n301), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n378), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT79), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n377), .A2(new_n373), .A3(new_n378), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n389), .A2(KEYINPUT30), .A3(new_n353), .A4(new_n356), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n353), .B1(new_n372), .B2(new_n379), .ZN(new_n391));
  INV_X1    g190(.A(new_n356), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n382), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(G1gat), .B(G29gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n395), .B(KEYINPUT0), .ZN(new_n396));
  XNOR2_X1  g195(.A(G57gat), .B(G85gat), .ZN(new_n397));
  XOR2_X1   g196(.A(new_n396), .B(new_n397), .Z(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  OR2_X1    g198(.A1(G141gat), .A2(G148gat), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT2), .ZN(new_n401));
  NAND2_X1  g200(.A1(G141gat), .A2(G148gat), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(G162gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(G155gat), .ZN(new_n405));
  INV_X1    g204(.A(G155gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(G162gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n403), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT81), .B(G162gat), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n401), .B1(new_n410), .B2(G155gat), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n400), .A2(new_n405), .A3(new_n407), .A4(new_n402), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AND2_X1   g212(.A1(G113gat), .A2(G120gat), .ZN(new_n414));
  NOR2_X1   g213(.A1(G113gat), .A2(G120gat), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AND2_X1   g215(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n417));
  NOR2_X1   g216(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G127gat), .B(G134gat), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n416), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(G113gat), .ZN(new_n422));
  INV_X1    g221(.A(G120gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT1), .ZN(new_n425));
  NAND2_X1  g224(.A1(G113gat), .A2(G120gat), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(G134gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(G127gat), .ZN(new_n429));
  INV_X1    g228(.A(G127gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(G134gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n421), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT84), .B1(new_n413), .B2(new_n434), .ZN(new_n435));
  AND2_X1   g234(.A1(KEYINPUT81), .A2(G162gat), .ZN(new_n436));
  NOR2_X1   g235(.A1(KEYINPUT81), .A2(G162gat), .ZN(new_n437));
  OAI21_X1  g236(.A(G155gat), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT2), .ZN(new_n439));
  AND4_X1   g238(.A1(new_n405), .A2(new_n400), .A3(new_n407), .A4(new_n402), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n439), .A2(new_n440), .B1(new_n408), .B2(new_n403), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n421), .A2(new_n433), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT84), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n435), .A2(new_n444), .B1(new_n413), .B2(new_n434), .ZN(new_n445));
  NAND2_X1  g244(.A1(G225gat), .A2(G233gat), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT5), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n446), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n442), .B1(KEYINPUT3), .B2(new_n413), .ZN(new_n449));
  XNOR2_X1  g248(.A(KEYINPUT82), .B(KEYINPUT3), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n441), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n448), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT70), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n434), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n421), .A2(new_n433), .A3(KEYINPUT70), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(new_n441), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT83), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT4), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT4), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n435), .A2(new_n444), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n457), .B1(new_n456), .B2(KEYINPUT4), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n452), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT85), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(KEYINPUT85), .B(new_n452), .C1(new_n461), .C2(new_n462), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n447), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT5), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n456), .A2(new_n459), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n435), .A2(new_n444), .A3(KEYINPUT4), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n452), .A2(new_n468), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n399), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n445), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT39), .B1(new_n474), .B2(new_n448), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n449), .A2(new_n451), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n470), .A2(new_n476), .A3(new_n469), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n475), .B1(new_n448), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n448), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n398), .B1(new_n479), .B2(KEYINPUT39), .ZN(new_n480));
  NOR2_X1   g279(.A1(KEYINPUT90), .A2(KEYINPUT40), .ZN(new_n481));
  OR3_X1    g280(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n481), .B1(new_n478), .B2(new_n480), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n473), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n394), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(G228gat), .A2(G233gat), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n450), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n301), .B1(new_n413), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n344), .A2(new_n347), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT29), .B1(new_n345), .B2(new_n346), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n413), .B1(new_n491), .B2(new_n488), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n487), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(KEYINPUT87), .ZN(new_n494));
  INV_X1    g293(.A(G22gat), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n413), .B1(new_n491), .B2(KEYINPUT3), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n490), .A2(new_n496), .A3(new_n487), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n494), .A2(KEYINPUT88), .A3(new_n495), .A4(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n493), .A2(KEYINPUT87), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT87), .ZN(new_n500));
  AOI211_X1 g299(.A(new_n500), .B(new_n487), .C1(new_n490), .C2(new_n492), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n495), .B(new_n497), .C1(new_n499), .C2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT88), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n497), .B1(new_n499), .B2(new_n501), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(G22gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n498), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G78gat), .B(G106gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT31), .B(G50gat), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n508), .B(new_n509), .Z(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT86), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n510), .B1(new_n505), .B2(G22gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n502), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT38), .ZN(new_n516));
  XOR2_X1   g315(.A(KEYINPUT91), .B(KEYINPUT37), .Z(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n353), .B(new_n518), .C1(new_n372), .C2(new_n379), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n519), .A2(new_n392), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n391), .A2(KEYINPUT37), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n516), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n447), .ZN(new_n523));
  INV_X1    g322(.A(new_n466), .ZN(new_n524));
  AND3_X1   g323(.A1(new_n421), .A2(new_n433), .A3(KEYINPUT70), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT70), .B1(new_n421), .B2(new_n433), .ZN(new_n526));
  NOR3_X1   g325(.A1(new_n525), .A2(new_n526), .A3(new_n413), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT83), .B1(new_n527), .B2(new_n459), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n528), .A2(new_n460), .A3(new_n458), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT85), .B1(new_n529), .B2(new_n452), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n523), .B1(new_n524), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n531), .A2(new_n398), .A3(new_n471), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT6), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n473), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  OAI211_X1 g333(.A(KEYINPUT6), .B(new_n399), .C1(new_n467), .C2(new_n472), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n377), .A2(new_n348), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT37), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n537), .B1(new_n315), .B2(new_n378), .ZN(new_n538));
  AOI211_X1 g337(.A(KEYINPUT38), .B(new_n356), .C1(new_n536), .C2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n519), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n534), .A2(new_n535), .A3(new_n380), .A4(new_n540), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n485), .B(new_n515), .C1(new_n522), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT92), .ZN(new_n543));
  INV_X1    g342(.A(new_n521), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n519), .A2(new_n392), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT38), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n534), .A2(new_n535), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n540), .A2(new_n380), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n507), .A2(new_n511), .B1(new_n513), .B2(new_n502), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n550), .B1(new_n394), .B2(new_n484), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT92), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n549), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n543), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n550), .B1(new_n547), .B2(new_n394), .ZN(new_n555));
  INV_X1    g354(.A(G227gat), .ZN(new_n556));
  INV_X1    g355(.A(G233gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT64), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n525), .A2(new_n526), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n314), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n560), .B1(new_n366), .B2(new_n310), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n559), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT33), .ZN(new_n565));
  XNOR2_X1  g364(.A(G15gat), .B(G43gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(G71gat), .B(G99gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n564), .B(KEYINPUT32), .C1(new_n565), .C2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n568), .B1(new_n564), .B2(new_n565), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT71), .ZN(new_n572));
  INV_X1    g371(.A(new_n559), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n370), .A2(new_n560), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n314), .A2(new_n561), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT32), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n572), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n564), .A2(KEYINPUT71), .A3(KEYINPUT32), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n571), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT72), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT72), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n571), .A2(new_n578), .A3(new_n579), .A4(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n570), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n562), .A2(new_n563), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n559), .A2(KEYINPUT34), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n574), .B(new_n575), .C1(new_n556), .C2(new_n557), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT73), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n588), .A2(new_n589), .A3(KEYINPUT34), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n589), .B1(new_n588), .B2(KEYINPUT34), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n587), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n584), .A2(new_n593), .ZN(new_n594));
  AOI211_X1 g393(.A(new_n570), .B(new_n592), .C1(new_n581), .C2(new_n583), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT36), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n583), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n569), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(new_n592), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT36), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n593), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n555), .A2(new_n596), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT89), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT89), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n555), .A2(new_n605), .A3(new_n596), .A4(new_n602), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n554), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n599), .A2(new_n515), .A3(new_n601), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n382), .A2(new_n390), .A3(new_n393), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n534), .A2(new_n535), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(KEYINPUT35), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n394), .B1(new_n535), .B2(new_n534), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n594), .A2(new_n595), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT35), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n613), .A2(new_n614), .A3(new_n615), .A4(new_n515), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n255), .B1(new_n607), .B2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT97), .B(G57gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(G64gat), .ZN(new_n621));
  INV_X1    g420(.A(G64gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(G57gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(G71gat), .ZN(new_n625));
  INV_X1    g424(.A(G78gat), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(G71gat), .A2(G78gat), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n627), .B1(KEYINPUT9), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n623), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n622), .A2(G57gat), .ZN(new_n632));
  OAI21_X1  g431(.A(KEYINPUT9), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n627), .A2(new_n628), .ZN(new_n634));
  AOI22_X1  g433(.A1(new_n624), .A2(new_n630), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT98), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n634), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n631), .B1(new_n620), .B2(G64gat), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n638), .B1(new_n639), .B2(new_n629), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(KEYINPUT98), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n242), .B1(new_n642), .B2(KEYINPUT21), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT101), .B(KEYINPUT20), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n642), .ZN(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT99), .B(KEYINPUT21), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(G231gat), .A2(G233gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n650), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n649), .B(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n652), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(G127gat), .B(G155gat), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g459(.A(G183gat), .B(G211gat), .Z(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n659), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n653), .A2(new_n657), .A3(new_n663), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n660), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n662), .B1(new_n660), .B2(new_n664), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n646), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n660), .A2(new_n664), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n661), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n660), .A2(new_n662), .A3(new_n664), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n669), .A2(new_n645), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(G134gat), .B(G162gat), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT102), .B(KEYINPUT7), .ZN(new_n678));
  NAND2_X1  g477(.A1(G85gat), .A2(G92gat), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  NAND2_X1  g480(.A1(G99gat), .A2(G106gat), .ZN(new_n682));
  INV_X1    g481(.A(G85gat), .ZN(new_n683));
  INV_X1    g482(.A(G92gat), .ZN(new_n684));
  AOI22_X1  g483(.A1(KEYINPUT8), .A2(new_n682), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n680), .A2(new_n681), .A3(new_n685), .ZN(new_n686));
  XOR2_X1   g485(.A(G99gat), .B(G106gat), .Z(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n687), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n680), .A2(new_n689), .A3(new_n681), .A4(new_n685), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n231), .A2(new_n238), .A3(new_n691), .ZN(new_n692));
  AND3_X1   g491(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n688), .A2(new_n690), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n693), .B1(new_n241), .B2(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(G190gat), .B(G218gat), .Z(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n692), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n697), .B1(new_n692), .B2(new_n695), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n677), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n700), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n702), .A2(new_n676), .A3(new_n698), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(G230gat), .A2(G233gat), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(new_n642), .B2(new_n694), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n691), .A2(KEYINPUT103), .A3(new_n637), .A4(new_n641), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT10), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n694), .A2(new_n712), .A3(new_n635), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT104), .B1(new_n691), .B2(new_n640), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n710), .A2(new_n711), .A3(new_n715), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n647), .A2(new_n711), .A3(new_n691), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n706), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(G120gat), .B(G148gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(G176gat), .B(G204gat), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n719), .B(new_n720), .Z(new_n721));
  AOI22_X1  g520(.A1(new_n708), .A2(new_n709), .B1(new_n713), .B2(new_n714), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n718), .B(new_n721), .C1(new_n706), .C2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n721), .ZN(new_n724));
  INV_X1    g523(.A(new_n706), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n722), .A2(new_n711), .ZN(new_n726));
  INV_X1    g525(.A(new_n717), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n722), .A2(new_n706), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n724), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n723), .A2(new_n730), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n673), .A2(new_n705), .A3(new_n731), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n619), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n547), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g534(.A1(new_n619), .A2(new_n732), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(new_n609), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT105), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT105), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(new_n736), .B2(new_n609), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n738), .A2(G8gat), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(KEYINPUT16), .B(G8gat), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT42), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n737), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n742), .B1(new_n738), .B2(new_n740), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n741), .B(new_n745), .C1(new_n746), .C2(KEYINPUT42), .ZN(G1325gat));
  NAND2_X1  g546(.A1(new_n602), .A2(new_n596), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(G15gat), .B1(new_n736), .B2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n614), .ZN(new_n751));
  OR2_X1    g550(.A1(new_n751), .A2(G15gat), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n736), .B2(new_n752), .ZN(G1326gat));
  NAND2_X1  g552(.A1(new_n733), .A2(new_n550), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT106), .ZN(new_n755));
  XNOR2_X1  g554(.A(KEYINPUT43), .B(G22gat), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n754), .A2(KEYINPUT106), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n754), .A2(KEYINPUT106), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n759), .A2(new_n760), .A3(new_n756), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n758), .A2(new_n761), .ZN(G1327gat));
  INV_X1    g561(.A(new_n731), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n673), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n704), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n619), .A2(new_n765), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n766), .A2(G29gat), .A3(new_n610), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n767), .B(KEYINPUT45), .Z(new_n768));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n705), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n603), .B1(new_n543), .B2(new_n553), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n617), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n555), .A2(new_n596), .A3(new_n602), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n542), .A2(KEYINPUT92), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n552), .B1(new_n549), .B2(new_n551), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT108), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n770), .B1(new_n773), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n607), .A2(new_n618), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n705), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT44), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT107), .ZN(new_n785));
  INV_X1    g584(.A(new_n253), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n786), .B2(new_n251), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n252), .A2(KEYINPUT107), .A3(new_n253), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n764), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n784), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(G29gat), .B1(new_n792), .B2(new_n610), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n768), .A2(new_n793), .ZN(G1328gat));
  INV_X1    g593(.A(new_n791), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n795), .B1(new_n780), .B2(new_n783), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n208), .B1(new_n796), .B2(new_n394), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n619), .A2(new_n208), .A3(new_n394), .A4(new_n765), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT46), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT109), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT46), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n798), .B(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT109), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n769), .B1(new_n781), .B2(new_n705), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n394), .B(new_n791), .C1(new_n804), .C2(new_n779), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n802), .B(new_n803), .C1(new_n806), .C2(new_n208), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n800), .A2(new_n807), .ZN(G1329gat));
  NAND4_X1  g607(.A1(new_n784), .A2(G43gat), .A3(new_n748), .A4(new_n791), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT47), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT110), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n810), .A2(KEYINPUT110), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n619), .A2(new_n614), .A3(new_n765), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n812), .B1(new_n813), .B2(new_n225), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n809), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n811), .B1(new_n809), .B2(new_n814), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(G1330gat));
  OAI21_X1  g616(.A(new_n223), .B1(new_n766), .B2(new_n515), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n515), .A2(new_n223), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n818), .B1(new_n792), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT48), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT48), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n823), .B(new_n818), .C1(new_n792), .C2(new_n820), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(G1331gat));
  NAND4_X1  g624(.A1(new_n672), .A2(new_n704), .A3(new_n731), .A4(new_n790), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n618), .B1(new_n777), .B2(KEYINPUT108), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n771), .A2(new_n772), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(new_n610), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(new_n620), .ZN(G1332gat));
  NAND2_X1  g631(.A1(new_n830), .A2(KEYINPUT111), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n773), .A2(new_n778), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT111), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n835), .A3(new_n827), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  OAI22_X1  g636(.A1(new_n837), .A2(new_n609), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n838));
  XNOR2_X1  g637(.A(KEYINPUT49), .B(G64gat), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n833), .A2(new_n394), .A3(new_n836), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(G1333gat));
  INV_X1    g640(.A(KEYINPUT50), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n833), .A2(new_n748), .A3(new_n836), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(G71gat), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n830), .A2(G71gat), .A3(new_n751), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n842), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  AOI211_X1 g646(.A(KEYINPUT50), .B(new_n845), .C1(new_n843), .C2(G71gat), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(G1334gat));
  NOR2_X1   g648(.A1(new_n837), .A2(new_n515), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(new_n626), .ZN(G1335gat));
  OR3_X1    g650(.A1(new_n672), .A2(KEYINPUT112), .A3(new_n789), .ZN(new_n852));
  OAI21_X1  g651(.A(KEYINPUT112), .B1(new_n672), .B2(new_n789), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n731), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n784), .A2(new_n547), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(G85gat), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n704), .B1(new_n852), .B2(new_n853), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n834), .A2(new_n859), .A3(KEYINPUT51), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT51), .B1(new_n834), .B2(new_n859), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n547), .A2(new_n731), .A3(new_n683), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n858), .B1(new_n862), .B2(new_n863), .ZN(G1336gat));
  OAI211_X1 g663(.A(new_n394), .B(new_n856), .C1(new_n804), .C2(new_n779), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(G92gat), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT113), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n609), .A2(new_n763), .A3(G92gat), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n868), .B1(new_n860), .B2(new_n861), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n867), .A2(new_n870), .A3(KEYINPUT52), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n866), .B(new_n869), .C1(KEYINPUT113), .C2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(G1337gat));
  OAI211_X1 g673(.A(new_n748), .B(new_n856), .C1(new_n804), .C2(new_n779), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT114), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(G99gat), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n875), .A2(KEYINPUT114), .ZN(new_n878));
  OR3_X1    g677(.A1(new_n751), .A2(G99gat), .A3(new_n763), .ZN(new_n879));
  OAI22_X1  g678(.A1(new_n877), .A2(new_n878), .B1(new_n862), .B2(new_n879), .ZN(G1338gat));
  NOR3_X1   g679(.A1(new_n515), .A2(new_n763), .A3(G106gat), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n881), .B1(new_n860), .B2(new_n861), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n550), .B(new_n856), .C1(new_n804), .C2(new_n779), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(G106gat), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(KEYINPUT53), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n882), .B(new_n888), .C1(new_n884), .C2(new_n885), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(G1339gat));
  AND4_X1   g689(.A1(new_n672), .A2(new_n704), .A3(new_n763), .A4(new_n790), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT115), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n892), .B1(new_n247), .B2(new_n248), .ZN(new_n893));
  INV_X1    g692(.A(new_n248), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n243), .A2(KEYINPUT115), .A3(new_n246), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n240), .B1(new_n239), .B2(new_n243), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n205), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AND4_X1   g697(.A1(new_n253), .A2(new_n898), .A3(new_n703), .A4(new_n701), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT55), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n726), .A2(new_n725), .A3(new_n727), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n718), .A2(KEYINPUT54), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n724), .B1(new_n718), .B2(KEYINPUT54), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT54), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n721), .B1(new_n728), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n718), .A2(new_n901), .A3(KEYINPUT54), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT55), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n899), .A2(new_n904), .A3(new_n723), .A4(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT116), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n908), .A2(new_n723), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT116), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n911), .A2(new_n912), .A3(new_n904), .A4(new_n899), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n731), .A2(new_n253), .A3(new_n898), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n908), .A2(new_n723), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT55), .B1(new_n906), .B2(new_n907), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n915), .B1(new_n918), .B2(new_n789), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n910), .B(new_n913), .C1(new_n919), .C2(new_n705), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n891), .B1(new_n920), .B2(new_n673), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n921), .A2(new_n608), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n610), .A2(new_n394), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n924), .A2(new_n422), .A3(new_n255), .ZN(new_n925));
  INV_X1    g724(.A(new_n924), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n789), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n925), .B1(new_n422), .B2(new_n927), .ZN(G1340gat));
  OAI21_X1  g727(.A(G120gat), .B1(new_n924), .B2(new_n763), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n929), .A2(KEYINPUT117), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n929), .A2(KEYINPUT117), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n731), .A2(new_n423), .ZN(new_n932));
  XOR2_X1   g731(.A(new_n932), .B(KEYINPUT118), .Z(new_n933));
  OAI22_X1  g732(.A1(new_n930), .A2(new_n931), .B1(new_n924), .B2(new_n933), .ZN(G1341gat));
  NOR2_X1   g733(.A1(new_n924), .A2(new_n673), .ZN(new_n935));
  XNOR2_X1  g734(.A(KEYINPUT119), .B(G127gat), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n935), .B(new_n936), .ZN(G1342gat));
  AOI211_X1 g736(.A(new_n704), .B(new_n924), .C1(KEYINPUT56), .C2(G134gat), .ZN(new_n938));
  NOR2_X1   g737(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n938), .B(new_n939), .ZN(G1343gat));
  INV_X1    g739(.A(KEYINPUT120), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n789), .A2(new_n911), .A3(new_n904), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n705), .B1(new_n942), .B2(new_n914), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n910), .A2(new_n913), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n673), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n672), .A2(new_n704), .A3(new_n763), .A4(new_n790), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n515), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n941), .B1(new_n947), .B2(KEYINPUT57), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT57), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n515), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n904), .A2(new_n254), .A3(new_n723), .A4(new_n908), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(new_n914), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT121), .B1(new_n952), .B2(new_n704), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n953), .A2(new_n944), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n705), .B1(new_n951), .B2(new_n914), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(KEYINPUT121), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n672), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n950), .B1(new_n957), .B2(new_n891), .ZN(new_n958));
  OAI211_X1 g757(.A(KEYINPUT120), .B(new_n949), .C1(new_n921), .C2(new_n515), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n948), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n749), .A2(new_n923), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n960), .A2(new_n254), .A3(new_n962), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n963), .A2(G141gat), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n945), .A2(new_n946), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(new_n550), .ZN(new_n966));
  NOR4_X1   g765(.A1(new_n966), .A2(G141gat), .A3(new_n255), .A4(new_n961), .ZN(new_n967));
  XNOR2_X1  g766(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n960), .A2(new_n789), .A3(new_n962), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n967), .B1(new_n970), .B2(G141gat), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT58), .ZN(new_n972));
  OAI22_X1  g771(.A1(new_n964), .A2(new_n969), .B1(new_n971), .B2(new_n972), .ZN(G1344gat));
  INV_X1    g772(.A(G148gat), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n974), .A2(KEYINPUT59), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n962), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n975), .B1(new_n976), .B2(new_n763), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n966), .A2(KEYINPUT57), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n732), .A2(new_n255), .ZN(new_n979));
  INV_X1    g778(.A(new_n909), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n673), .B1(new_n955), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n982), .A2(new_n949), .A3(new_n550), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n978), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n962), .A2(new_n731), .ZN(new_n985));
  OAI21_X1  g784(.A(G148gat), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(KEYINPUT59), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n977), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n966), .A2(new_n961), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n989), .A2(new_n974), .A3(new_n731), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n988), .A2(new_n990), .ZN(G1345gat));
  OAI21_X1  g790(.A(G155gat), .B1(new_n976), .B2(new_n673), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n989), .A2(new_n406), .A3(new_n672), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n992), .A2(new_n993), .ZN(G1346gat));
  OAI21_X1  g793(.A(new_n410), .B1(new_n976), .B2(new_n704), .ZN(new_n995));
  INV_X1    g794(.A(new_n410), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n989), .A2(new_n996), .A3(new_n705), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n995), .A2(new_n997), .ZN(G1347gat));
  NOR2_X1   g797(.A1(new_n547), .A2(new_n609), .ZN(new_n999));
  AND2_X1   g798(.A1(new_n922), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g799(.A(G169gat), .B1(new_n1000), .B2(new_n789), .ZN(new_n1001));
  AND2_X1   g800(.A1(new_n254), .A2(G169gat), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n1001), .B1(new_n1000), .B2(new_n1002), .ZN(G1348gat));
  NAND2_X1  g802(.A1(new_n1000), .A2(new_n731), .ZN(new_n1004));
  XNOR2_X1  g803(.A(new_n1004), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g804(.A1(new_n1000), .A2(new_n264), .A3(new_n672), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1006), .A2(KEYINPUT123), .ZN(new_n1007));
  AOI21_X1  g806(.A(new_n256), .B1(new_n1000), .B2(new_n672), .ZN(new_n1008));
  OAI21_X1  g807(.A(KEYINPUT60), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g808(.A(new_n1008), .ZN(new_n1010));
  INV_X1    g809(.A(KEYINPUT60), .ZN(new_n1011));
  NAND4_X1  g810(.A1(new_n1010), .A2(KEYINPUT123), .A3(new_n1011), .A4(new_n1006), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1009), .A2(new_n1012), .ZN(G1350gat));
  NAND2_X1  g812(.A1(new_n1000), .A2(new_n705), .ZN(new_n1014));
  INV_X1    g813(.A(KEYINPUT124), .ZN(new_n1015));
  AOI21_X1  g814(.A(new_n260), .B1(new_n1015), .B2(KEYINPUT61), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g816(.A(KEYINPUT61), .ZN(new_n1018));
  NAND3_X1  g817(.A1(new_n1017), .A2(KEYINPUT124), .A3(new_n1018), .ZN(new_n1019));
  OAI211_X1 g818(.A(new_n1014), .B(new_n1016), .C1(new_n1015), .C2(KEYINPUT61), .ZN(new_n1020));
  OAI211_X1 g819(.A(new_n1019), .B(new_n1020), .C1(G190gat), .C2(new_n1014), .ZN(G1351gat));
  NAND2_X1  g820(.A1(new_n749), .A2(new_n999), .ZN(new_n1022));
  INV_X1    g821(.A(new_n1022), .ZN(new_n1023));
  NAND3_X1  g822(.A1(new_n978), .A2(new_n983), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g823(.A(G197gat), .B1(new_n1024), .B2(new_n255), .ZN(new_n1025));
  INV_X1    g824(.A(KEYINPUT125), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n947), .A2(new_n1023), .ZN(new_n1027));
  OR3_X1    g826(.A1(new_n1027), .A2(G197gat), .A3(new_n790), .ZN(new_n1028));
  AND3_X1   g827(.A1(new_n1025), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g828(.A(new_n1026), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1030));
  NOR2_X1   g829(.A1(new_n1029), .A2(new_n1030), .ZN(G1352gat));
  XOR2_X1   g830(.A(KEYINPUT126), .B(G204gat), .Z(new_n1032));
  NOR3_X1   g831(.A1(new_n1027), .A2(new_n763), .A3(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g832(.A(new_n1033), .B(KEYINPUT62), .ZN(new_n1034));
  OAI21_X1  g833(.A(new_n1032), .B1(new_n1024), .B2(new_n763), .ZN(new_n1035));
  NAND2_X1  g834(.A1(new_n1034), .A2(new_n1035), .ZN(G1353gat));
  NAND4_X1  g835(.A1(new_n978), .A2(new_n983), .A3(new_n672), .A4(new_n1023), .ZN(new_n1037));
  NAND3_X1  g836(.A1(new_n1037), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1038));
  INV_X1    g837(.A(new_n1038), .ZN(new_n1039));
  AOI21_X1  g838(.A(KEYINPUT63), .B1(new_n1037), .B2(G211gat), .ZN(new_n1040));
  NAND2_X1  g839(.A1(new_n672), .A2(new_n318), .ZN(new_n1041));
  OAI22_X1  g840(.A1(new_n1039), .A2(new_n1040), .B1(new_n1027), .B2(new_n1041), .ZN(G1354gat));
  OAI21_X1  g841(.A(new_n329), .B1(new_n1027), .B2(new_n704), .ZN(new_n1043));
  OAI21_X1  g842(.A(new_n705), .B1(new_n339), .B2(new_n338), .ZN(new_n1044));
  XNOR2_X1  g843(.A(new_n1044), .B(KEYINPUT127), .ZN(new_n1045));
  OAI21_X1  g844(.A(new_n1043), .B1(new_n1024), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g845(.A(new_n1046), .ZN(G1355gat));
endmodule


