

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U552 ( .A(KEYINPUT66), .B(n522), .ZN(n653) );
  NOR2_X2 U553 ( .A1(n818), .A2(n817), .ZN(n820) );
  BUF_X2 U554 ( .A(n748), .Z(n517) );
  XOR2_X1 U555 ( .A(KEYINPUT17), .B(n615), .Z(n518) );
  NOR2_X2 U556 ( .A1(G2105), .A2(G2104), .ZN(n615) );
  NOR2_X2 U557 ( .A1(n693), .A2(n788), .ZN(n695) );
  NOR2_X2 U558 ( .A1(G164), .A2(G1384), .ZN(n789) );
  XNOR2_X2 U559 ( .A(n552), .B(n551), .ZN(G164) );
  NAND2_X1 U560 ( .A1(n720), .A2(n721), .ZN(n710) );
  XNOR2_X1 U561 ( .A(n591), .B(KEYINPUT15), .ZN(n720) );
  NOR2_X1 U562 ( .A1(G651), .A2(n638), .ZN(n660) );
  NOR2_X1 U563 ( .A1(n638), .A2(n527), .ZN(n656) );
  XNOR2_X1 U564 ( .A(n586), .B(KEYINPUT75), .ZN(n519) );
  INV_X1 U565 ( .A(KEYINPUT99), .ZN(n732) );
  NOR2_X1 U566 ( .A1(n719), .A2(n718), .ZN(n723) );
  NOR2_X1 U567 ( .A1(G168), .A2(n736), .ZN(n737) );
  INV_X1 U568 ( .A(KEYINPUT31), .ZN(n741) );
  INV_X1 U569 ( .A(KEYINPUT32), .ZN(n761) );
  XNOR2_X1 U570 ( .A(n762), .B(n761), .ZN(n763) );
  NAND2_X1 U571 ( .A1(n748), .A2(G8), .ZN(n731) );
  INV_X1 U572 ( .A(G651), .ZN(n527) );
  NOR2_X2 U573 ( .A1(G2105), .A2(n538), .ZN(n894) );
  INV_X1 U574 ( .A(n720), .ZN(n975) );
  NOR2_X1 U575 ( .A1(n543), .A2(n542), .ZN(G160) );
  XNOR2_X1 U576 ( .A(G543), .B(KEYINPUT0), .ZN(n520) );
  XNOR2_X1 U577 ( .A(n520), .B(KEYINPUT65), .ZN(n638) );
  NAND2_X1 U578 ( .A1(G51), .A2(n660), .ZN(n524) );
  NOR2_X1 U579 ( .A1(G543), .A2(n527), .ZN(n521) );
  XOR2_X1 U580 ( .A(KEYINPUT1), .B(n521), .Z(n522) );
  NAND2_X1 U581 ( .A1(G63), .A2(n653), .ZN(n523) );
  NAND2_X1 U582 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U583 ( .A(KEYINPUT6), .B(n525), .ZN(n533) );
  NOR2_X1 U584 ( .A1(G651), .A2(G543), .ZN(n652) );
  NAND2_X1 U585 ( .A1(n652), .A2(G89), .ZN(n526) );
  XNOR2_X1 U586 ( .A(n526), .B(KEYINPUT4), .ZN(n529) );
  NAND2_X1 U587 ( .A1(G76), .A2(n656), .ZN(n528) );
  NAND2_X1 U588 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U589 ( .A(KEYINPUT77), .B(n530), .ZN(n531) );
  XNOR2_X1 U590 ( .A(KEYINPUT5), .B(n531), .ZN(n532) );
  NOR2_X1 U591 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U592 ( .A(KEYINPUT7), .B(n534), .Z(G168) );
  INV_X1 U593 ( .A(G2104), .ZN(n538) );
  AND2_X1 U594 ( .A1(n538), .A2(G2105), .ZN(n897) );
  NAND2_X1 U595 ( .A1(G125), .A2(n897), .ZN(n536) );
  AND2_X1 U596 ( .A1(G2105), .A2(G2104), .ZN(n898) );
  NAND2_X1 U597 ( .A1(G113), .A2(n898), .ZN(n535) );
  NAND2_X1 U598 ( .A1(n536), .A2(n535), .ZN(n543) );
  NAND2_X1 U599 ( .A1(G137), .A2(n518), .ZN(n537) );
  XNOR2_X1 U600 ( .A(n537), .B(KEYINPUT64), .ZN(n541) );
  NAND2_X1 U601 ( .A1(G101), .A2(n894), .ZN(n539) );
  XOR2_X1 U602 ( .A(KEYINPUT23), .B(n539), .Z(n540) );
  NAND2_X1 U603 ( .A1(n541), .A2(n540), .ZN(n542) );
  INV_X1 U604 ( .A(KEYINPUT89), .ZN(n552) );
  NAND2_X1 U605 ( .A1(G102), .A2(n894), .ZN(n545) );
  NAND2_X1 U606 ( .A1(G138), .A2(n518), .ZN(n544) );
  NAND2_X1 U607 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U608 ( .A(n546), .B(KEYINPUT88), .ZN(n550) );
  NAND2_X1 U609 ( .A1(G126), .A2(n897), .ZN(n548) );
  NAND2_X1 U610 ( .A1(G114), .A2(n898), .ZN(n547) );
  NAND2_X1 U611 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U612 ( .A1(n550), .A2(n549), .ZN(n551) );
  NAND2_X1 U613 ( .A1(G52), .A2(n660), .ZN(n554) );
  NAND2_X1 U614 ( .A1(G64), .A2(n653), .ZN(n553) );
  NAND2_X1 U615 ( .A1(n554), .A2(n553), .ZN(n560) );
  NAND2_X1 U616 ( .A1(n656), .A2(G77), .ZN(n555) );
  XNOR2_X1 U617 ( .A(n555), .B(KEYINPUT68), .ZN(n557) );
  NAND2_X1 U618 ( .A1(G90), .A2(n652), .ZN(n556) );
  NAND2_X1 U619 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U620 ( .A(KEYINPUT9), .B(n558), .Z(n559) );
  NOR2_X1 U621 ( .A1(n560), .A2(n559), .ZN(G171) );
  XOR2_X1 U622 ( .A(G2438), .B(G2454), .Z(n562) );
  XNOR2_X1 U623 ( .A(G2435), .B(G2430), .ZN(n561) );
  XNOR2_X1 U624 ( .A(n562), .B(n561), .ZN(n563) );
  XOR2_X1 U625 ( .A(n563), .B(G2427), .Z(n565) );
  INV_X1 U626 ( .A(G1341), .ZN(n1010) );
  XOR2_X1 U627 ( .A(n1010), .B(G1348), .Z(n564) );
  XNOR2_X1 U628 ( .A(n565), .B(n564), .ZN(n569) );
  XOR2_X1 U629 ( .A(G2443), .B(G2446), .Z(n567) );
  XNOR2_X1 U630 ( .A(KEYINPUT106), .B(G2451), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n567), .B(n566), .ZN(n568) );
  XOR2_X1 U632 ( .A(n569), .B(n568), .Z(n570) );
  AND2_X1 U633 ( .A1(G14), .A2(n570), .ZN(G401) );
  AND2_X1 U634 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U635 ( .A(G132), .ZN(G219) );
  INV_X1 U636 ( .A(G82), .ZN(G220) );
  INV_X1 U637 ( .A(G57), .ZN(G237) );
  XOR2_X1 U638 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U639 ( .A(KEYINPUT72), .B(KEYINPUT11), .Z(n574) );
  XOR2_X1 U640 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n572) );
  NAND2_X1 U641 ( .A1(G7), .A2(G661), .ZN(n571) );
  XOR2_X1 U642 ( .A(n572), .B(n571), .Z(n922) );
  NAND2_X1 U643 ( .A1(G567), .A2(n922), .ZN(n573) );
  XNOR2_X1 U644 ( .A(n574), .B(n573), .ZN(G234) );
  NAND2_X1 U645 ( .A1(n653), .A2(G56), .ZN(n575) );
  XOR2_X1 U646 ( .A(KEYINPUT14), .B(n575), .Z(n581) );
  NAND2_X1 U647 ( .A1(n652), .A2(G81), .ZN(n576) );
  XNOR2_X1 U648 ( .A(n576), .B(KEYINPUT12), .ZN(n578) );
  NAND2_X1 U649 ( .A1(G68), .A2(n656), .ZN(n577) );
  NAND2_X1 U650 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U651 ( .A(KEYINPUT13), .B(n579), .Z(n580) );
  NOR2_X1 U652 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U653 ( .A1(n660), .A2(G43), .ZN(n582) );
  NAND2_X1 U654 ( .A1(n583), .A2(n582), .ZN(n983) );
  XNOR2_X1 U655 ( .A(G860), .B(KEYINPUT73), .ZN(n605) );
  OR2_X1 U656 ( .A1(n983), .A2(n605), .ZN(G153) );
  XOR2_X1 U657 ( .A(G171), .B(KEYINPUT74), .Z(G301) );
  NAND2_X1 U658 ( .A1(G868), .A2(G301), .ZN(n593) );
  NAND2_X1 U659 ( .A1(n652), .A2(G92), .ZN(n585) );
  NAND2_X1 U660 ( .A1(G66), .A2(n653), .ZN(n584) );
  NAND2_X1 U661 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U662 ( .A1(G54), .A2(n660), .ZN(n587) );
  NAND2_X1 U663 ( .A1(n519), .A2(n587), .ZN(n590) );
  NAND2_X1 U664 ( .A1(n656), .A2(G79), .ZN(n588) );
  XOR2_X1 U665 ( .A(KEYINPUT76), .B(n588), .Z(n589) );
  NOR2_X1 U666 ( .A1(n590), .A2(n589), .ZN(n591) );
  INV_X1 U667 ( .A(G868), .ZN(n602) );
  NAND2_X1 U668 ( .A1(n720), .A2(n602), .ZN(n592) );
  NAND2_X1 U669 ( .A1(n593), .A2(n592), .ZN(G284) );
  NAND2_X1 U670 ( .A1(G53), .A2(n660), .ZN(n595) );
  NAND2_X1 U671 ( .A1(G65), .A2(n653), .ZN(n594) );
  NAND2_X1 U672 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U673 ( .A(KEYINPUT70), .B(n596), .ZN(n599) );
  NAND2_X1 U674 ( .A1(G91), .A2(n652), .ZN(n597) );
  XNOR2_X1 U675 ( .A(KEYINPUT69), .B(n597), .ZN(n598) );
  NOR2_X1 U676 ( .A1(n599), .A2(n598), .ZN(n601) );
  NAND2_X1 U677 ( .A1(n656), .A2(G78), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n601), .A2(n600), .ZN(G299) );
  NOR2_X1 U679 ( .A1(G286), .A2(n602), .ZN(n604) );
  NOR2_X1 U680 ( .A1(G868), .A2(G299), .ZN(n603) );
  NOR2_X1 U681 ( .A1(n604), .A2(n603), .ZN(G297) );
  NAND2_X1 U682 ( .A1(n605), .A2(G559), .ZN(n606) );
  NAND2_X1 U683 ( .A1(n606), .A2(n975), .ZN(n607) );
  XNOR2_X1 U684 ( .A(n607), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U685 ( .A1(n975), .A2(G868), .ZN(n608) );
  NOR2_X1 U686 ( .A1(G559), .A2(n608), .ZN(n609) );
  XNOR2_X1 U687 ( .A(n609), .B(KEYINPUT78), .ZN(n611) );
  NOR2_X1 U688 ( .A1(n983), .A2(G868), .ZN(n610) );
  NOR2_X1 U689 ( .A1(n611), .A2(n610), .ZN(G282) );
  NAND2_X1 U690 ( .A1(G123), .A2(n897), .ZN(n612) );
  XNOR2_X1 U691 ( .A(n612), .B(KEYINPUT18), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n894), .A2(G99), .ZN(n613) );
  NAND2_X1 U693 ( .A1(n614), .A2(n613), .ZN(n619) );
  XOR2_X1 U694 ( .A(KEYINPUT17), .B(n615), .Z(n893) );
  NAND2_X1 U695 ( .A1(G135), .A2(n893), .ZN(n617) );
  NAND2_X1 U696 ( .A1(G111), .A2(n898), .ZN(n616) );
  NAND2_X1 U697 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U698 ( .A1(n619), .A2(n618), .ZN(n924) );
  XNOR2_X1 U699 ( .A(n924), .B(G2096), .ZN(n620) );
  INV_X1 U700 ( .A(G2100), .ZN(n856) );
  NAND2_X1 U701 ( .A1(n620), .A2(n856), .ZN(G156) );
  NAND2_X1 U702 ( .A1(G55), .A2(n660), .ZN(n622) );
  NAND2_X1 U703 ( .A1(G67), .A2(n653), .ZN(n621) );
  NAND2_X1 U704 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U705 ( .A1(G93), .A2(n652), .ZN(n624) );
  NAND2_X1 U706 ( .A1(G80), .A2(n656), .ZN(n623) );
  NAND2_X1 U707 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U708 ( .A1(n626), .A2(n625), .ZN(n664) );
  NAND2_X1 U709 ( .A1(G559), .A2(n975), .ZN(n627) );
  XNOR2_X1 U710 ( .A(n627), .B(KEYINPUT79), .ZN(n671) );
  XOR2_X1 U711 ( .A(n671), .B(KEYINPUT80), .Z(n628) );
  XNOR2_X1 U712 ( .A(n983), .B(n628), .ZN(n629) );
  NOR2_X1 U713 ( .A1(G860), .A2(n629), .ZN(n630) );
  XNOR2_X1 U714 ( .A(n664), .B(n630), .ZN(G145) );
  NAND2_X1 U715 ( .A1(n652), .A2(G88), .ZN(n631) );
  XNOR2_X1 U716 ( .A(n631), .B(KEYINPUT82), .ZN(n633) );
  NAND2_X1 U717 ( .A1(G75), .A2(n656), .ZN(n632) );
  NAND2_X1 U718 ( .A1(n633), .A2(n632), .ZN(n637) );
  NAND2_X1 U719 ( .A1(G50), .A2(n660), .ZN(n635) );
  NAND2_X1 U720 ( .A1(G62), .A2(n653), .ZN(n634) );
  NAND2_X1 U721 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U722 ( .A1(n637), .A2(n636), .ZN(G166) );
  INV_X1 U723 ( .A(G166), .ZN(G303) );
  NAND2_X1 U724 ( .A1(G49), .A2(n660), .ZN(n640) );
  NAND2_X1 U725 ( .A1(G87), .A2(n638), .ZN(n639) );
  NAND2_X1 U726 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U727 ( .A1(n653), .A2(n641), .ZN(n644) );
  NAND2_X1 U728 ( .A1(G74), .A2(G651), .ZN(n642) );
  XOR2_X1 U729 ( .A(KEYINPUT81), .B(n642), .Z(n643) );
  NAND2_X1 U730 ( .A1(n644), .A2(n643), .ZN(G288) );
  NAND2_X1 U731 ( .A1(G85), .A2(n652), .ZN(n646) );
  NAND2_X1 U732 ( .A1(G72), .A2(n656), .ZN(n645) );
  NAND2_X1 U733 ( .A1(n646), .A2(n645), .ZN(n649) );
  NAND2_X1 U734 ( .A1(G47), .A2(n660), .ZN(n647) );
  XNOR2_X1 U735 ( .A(KEYINPUT67), .B(n647), .ZN(n648) );
  NOR2_X1 U736 ( .A1(n649), .A2(n648), .ZN(n651) );
  NAND2_X1 U737 ( .A1(G60), .A2(n653), .ZN(n650) );
  NAND2_X1 U738 ( .A1(n651), .A2(n650), .ZN(G290) );
  NAND2_X1 U739 ( .A1(n652), .A2(G86), .ZN(n655) );
  NAND2_X1 U740 ( .A1(G61), .A2(n653), .ZN(n654) );
  NAND2_X1 U741 ( .A1(n655), .A2(n654), .ZN(n659) );
  NAND2_X1 U742 ( .A1(n656), .A2(G73), .ZN(n657) );
  XOR2_X1 U743 ( .A(KEYINPUT2), .B(n657), .Z(n658) );
  NOR2_X1 U744 ( .A1(n659), .A2(n658), .ZN(n662) );
  NAND2_X1 U745 ( .A1(n660), .A2(G48), .ZN(n661) );
  NAND2_X1 U746 ( .A1(n662), .A2(n661), .ZN(G305) );
  NOR2_X1 U747 ( .A1(G868), .A2(n664), .ZN(n663) );
  XNOR2_X1 U748 ( .A(n663), .B(KEYINPUT83), .ZN(n674) );
  XOR2_X1 U749 ( .A(KEYINPUT19), .B(n664), .Z(n665) );
  XNOR2_X1 U750 ( .A(G288), .B(n665), .ZN(n666) );
  XOR2_X1 U751 ( .A(G303), .B(n666), .Z(n669) );
  XNOR2_X1 U752 ( .A(G290), .B(G305), .ZN(n667) );
  XNOR2_X1 U753 ( .A(n667), .B(n983), .ZN(n668) );
  XNOR2_X1 U754 ( .A(n669), .B(n668), .ZN(n670) );
  XOR2_X1 U755 ( .A(G299), .B(n670), .Z(n911) );
  XNOR2_X1 U756 ( .A(n911), .B(n671), .ZN(n672) );
  NAND2_X1 U757 ( .A1(G868), .A2(n672), .ZN(n673) );
  NAND2_X1 U758 ( .A1(n674), .A2(n673), .ZN(G295) );
  NAND2_X1 U759 ( .A1(G2078), .A2(G2084), .ZN(n675) );
  XOR2_X1 U760 ( .A(KEYINPUT20), .B(n675), .Z(n676) );
  NAND2_X1 U761 ( .A1(G2090), .A2(n676), .ZN(n677) );
  XNOR2_X1 U762 ( .A(KEYINPUT21), .B(n677), .ZN(n678) );
  NAND2_X1 U763 ( .A1(n678), .A2(G2072), .ZN(n679) );
  XNOR2_X1 U764 ( .A(KEYINPUT84), .B(n679), .ZN(G158) );
  XOR2_X1 U765 ( .A(KEYINPUT85), .B(G44), .Z(n680) );
  XNOR2_X1 U766 ( .A(KEYINPUT3), .B(n680), .ZN(G218) );
  NAND2_X1 U767 ( .A1(G120), .A2(G69), .ZN(n681) );
  NOR2_X1 U768 ( .A1(G237), .A2(n681), .ZN(n682) );
  XNOR2_X1 U769 ( .A(KEYINPUT86), .B(n682), .ZN(n683) );
  NAND2_X1 U770 ( .A1(n683), .A2(G108), .ZN(n842) );
  NAND2_X1 U771 ( .A1(G567), .A2(n842), .ZN(n684) );
  XNOR2_X1 U772 ( .A(n684), .B(KEYINPUT87), .ZN(n689) );
  NOR2_X1 U773 ( .A1(G220), .A2(G219), .ZN(n685) );
  XNOR2_X1 U774 ( .A(KEYINPUT22), .B(n685), .ZN(n686) );
  NAND2_X1 U775 ( .A1(n686), .A2(G96), .ZN(n687) );
  OR2_X1 U776 ( .A1(G218), .A2(n687), .ZN(n843) );
  AND2_X1 U777 ( .A1(G2106), .A2(n843), .ZN(n688) );
  NOR2_X1 U778 ( .A1(n689), .A2(n688), .ZN(G319) );
  INV_X1 U779 ( .A(G319), .ZN(n691) );
  NAND2_X1 U780 ( .A1(G661), .A2(G483), .ZN(n690) );
  NOR2_X1 U781 ( .A1(n691), .A2(n690), .ZN(n841) );
  NAND2_X1 U782 ( .A1(n841), .A2(G36), .ZN(G176) );
  INV_X1 U783 ( .A(n789), .ZN(n693) );
  NAND2_X1 U784 ( .A1(G160), .A2(G40), .ZN(n788) );
  INV_X1 U785 ( .A(n695), .ZN(n748) );
  INV_X1 U786 ( .A(n731), .ZN(n768) );
  INV_X1 U787 ( .A(n768), .ZN(n785) );
  NOR2_X1 U788 ( .A1(G1976), .A2(G288), .ZN(n766) );
  NAND2_X1 U789 ( .A1(n766), .A2(KEYINPUT33), .ZN(n694) );
  NOR2_X1 U790 ( .A1(n785), .A2(n694), .ZN(n773) );
  XNOR2_X1 U791 ( .A(G1961), .B(KEYINPUT93), .ZN(n1008) );
  NAND2_X1 U792 ( .A1(n517), .A2(n1008), .ZN(n697) );
  BUF_X2 U793 ( .A(n695), .Z(n707) );
  XNOR2_X1 U794 ( .A(KEYINPUT25), .B(G2078), .ZN(n957) );
  NAND2_X1 U795 ( .A1(n707), .A2(n957), .ZN(n696) );
  NAND2_X1 U796 ( .A1(n697), .A2(n696), .ZN(n738) );
  NAND2_X1 U797 ( .A1(n738), .A2(G171), .ZN(n730) );
  NAND2_X1 U798 ( .A1(G2072), .A2(n707), .ZN(n698) );
  XNOR2_X1 U799 ( .A(n698), .B(KEYINPUT27), .ZN(n699) );
  XNOR2_X1 U800 ( .A(KEYINPUT94), .B(n699), .ZN(n701) );
  XNOR2_X1 U801 ( .A(G1956), .B(KEYINPUT95), .ZN(n1009) );
  NOR2_X1 U802 ( .A1(n707), .A2(n1009), .ZN(n700) );
  NOR2_X1 U803 ( .A1(n701), .A2(n700), .ZN(n705) );
  INV_X1 U804 ( .A(G299), .ZN(n704) );
  NOR2_X1 U805 ( .A1(n705), .A2(n704), .ZN(n703) );
  XOR2_X1 U806 ( .A(KEYINPUT28), .B(KEYINPUT96), .Z(n702) );
  XNOR2_X1 U807 ( .A(n703), .B(n702), .ZN(n727) );
  NAND2_X1 U808 ( .A1(n705), .A2(n704), .ZN(n725) );
  XNOR2_X1 U809 ( .A(G1996), .B(KEYINPUT97), .ZN(n713) );
  INV_X1 U810 ( .A(n713), .ZN(n952) );
  XNOR2_X1 U811 ( .A(KEYINPUT26), .B(KEYINPUT98), .ZN(n714) );
  NOR2_X1 U812 ( .A1(n952), .A2(n714), .ZN(n706) );
  NOR2_X1 U813 ( .A1(n706), .A2(n983), .ZN(n711) );
  NAND2_X1 U814 ( .A1(G1348), .A2(n517), .ZN(n709) );
  NAND2_X1 U815 ( .A1(G2067), .A2(n707), .ZN(n708) );
  NAND2_X1 U816 ( .A1(n709), .A2(n708), .ZN(n721) );
  NAND2_X1 U817 ( .A1(n711), .A2(n710), .ZN(n719) );
  NAND2_X1 U818 ( .A1(n1010), .A2(n714), .ZN(n712) );
  NAND2_X1 U819 ( .A1(n712), .A2(n517), .ZN(n717) );
  NOR2_X1 U820 ( .A1(n517), .A2(n713), .ZN(n715) );
  NAND2_X1 U821 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U822 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U823 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U824 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U825 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U826 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U827 ( .A(KEYINPUT29), .B(n728), .Z(n729) );
  NAND2_X1 U828 ( .A1(n730), .A2(n729), .ZN(n754) );
  NOR2_X1 U829 ( .A1(n731), .A2(G1966), .ZN(n746) );
  NOR2_X1 U830 ( .A1(G2084), .A2(n517), .ZN(n743) );
  NOR2_X1 U831 ( .A1(n746), .A2(n743), .ZN(n733) );
  XNOR2_X1 U832 ( .A(n733), .B(n732), .ZN(n734) );
  NAND2_X1 U833 ( .A1(n734), .A2(G8), .ZN(n735) );
  XNOR2_X1 U834 ( .A(n735), .B(KEYINPUT30), .ZN(n736) );
  XNOR2_X1 U835 ( .A(n737), .B(KEYINPUT100), .ZN(n740) );
  NOR2_X1 U836 ( .A1(n738), .A2(G171), .ZN(n739) );
  NOR2_X1 U837 ( .A1(n740), .A2(n739), .ZN(n742) );
  XNOR2_X1 U838 ( .A(n742), .B(n741), .ZN(n756) );
  NAND2_X1 U839 ( .A1(n754), .A2(n756), .ZN(n745) );
  NAND2_X1 U840 ( .A1(G8), .A2(n743), .ZN(n744) );
  NAND2_X1 U841 ( .A1(n745), .A2(n744), .ZN(n747) );
  NOR2_X1 U842 ( .A1(n747), .A2(n746), .ZN(n764) );
  INV_X1 U843 ( .A(G8), .ZN(n753) );
  NOR2_X1 U844 ( .A1(G1971), .A2(n785), .ZN(n750) );
  NOR2_X1 U845 ( .A1(G2090), .A2(n517), .ZN(n749) );
  NOR2_X1 U846 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U847 ( .A1(n751), .A2(G303), .ZN(n752) );
  OR2_X1 U848 ( .A1(n753), .A2(n752), .ZN(n757) );
  AND2_X1 U849 ( .A1(n754), .A2(n757), .ZN(n755) );
  NAND2_X1 U850 ( .A1(n756), .A2(n755), .ZN(n760) );
  INV_X1 U851 ( .A(n757), .ZN(n758) );
  OR2_X1 U852 ( .A1(n758), .A2(G286), .ZN(n759) );
  NAND2_X1 U853 ( .A1(n760), .A2(n759), .ZN(n762) );
  NOR2_X2 U854 ( .A1(n764), .A2(n763), .ZN(n775) );
  NOR2_X1 U855 ( .A1(G1971), .A2(G303), .ZN(n765) );
  NOR2_X1 U856 ( .A1(n766), .A2(n765), .ZN(n985) );
  XNOR2_X1 U857 ( .A(KEYINPUT101), .B(n985), .ZN(n767) );
  NOR2_X1 U858 ( .A1(n775), .A2(n767), .ZN(n770) );
  NAND2_X1 U859 ( .A1(G1976), .A2(G288), .ZN(n984) );
  NAND2_X1 U860 ( .A1(n984), .A2(n768), .ZN(n769) );
  NOR2_X1 U861 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U862 ( .A1(n771), .A2(KEYINPUT33), .ZN(n772) );
  NOR2_X1 U863 ( .A1(n773), .A2(n772), .ZN(n774) );
  XOR2_X1 U864 ( .A(G1981), .B(G305), .Z(n980) );
  NAND2_X1 U865 ( .A1(n774), .A2(n980), .ZN(n781) );
  INV_X1 U866 ( .A(n775), .ZN(n778) );
  NOR2_X1 U867 ( .A1(G2090), .A2(G303), .ZN(n776) );
  NAND2_X1 U868 ( .A1(G8), .A2(n776), .ZN(n777) );
  NAND2_X1 U869 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U870 ( .A1(n779), .A2(n785), .ZN(n780) );
  NAND2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U872 ( .A(n782), .B(KEYINPUT102), .ZN(n787) );
  NOR2_X1 U873 ( .A1(G1981), .A2(G305), .ZN(n783) );
  XOR2_X1 U874 ( .A(n783), .B(KEYINPUT24), .Z(n784) );
  NOR2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U876 ( .A1(n787), .A2(n786), .ZN(n818) );
  NOR2_X1 U877 ( .A1(n789), .A2(n788), .ZN(n834) );
  XOR2_X1 U878 ( .A(G2067), .B(KEYINPUT37), .Z(n790) );
  XOR2_X1 U879 ( .A(KEYINPUT90), .B(n790), .Z(n821) );
  NAND2_X1 U880 ( .A1(G128), .A2(n897), .ZN(n792) );
  NAND2_X1 U881 ( .A1(G116), .A2(n898), .ZN(n791) );
  NAND2_X1 U882 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U883 ( .A(n793), .B(KEYINPUT35), .ZN(n798) );
  NAND2_X1 U884 ( .A1(G140), .A2(n893), .ZN(n795) );
  NAND2_X1 U885 ( .A1(G104), .A2(n894), .ZN(n794) );
  NAND2_X1 U886 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U887 ( .A(KEYINPUT34), .B(n796), .Z(n797) );
  NAND2_X1 U888 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U889 ( .A(n799), .B(KEYINPUT36), .Z(n905) );
  NOR2_X1 U890 ( .A1(n821), .A2(n905), .ZN(n937) );
  NAND2_X1 U891 ( .A1(n834), .A2(n937), .ZN(n831) );
  NAND2_X1 U892 ( .A1(G129), .A2(n897), .ZN(n801) );
  NAND2_X1 U893 ( .A1(G117), .A2(n898), .ZN(n800) );
  NAND2_X1 U894 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U895 ( .A(KEYINPUT92), .B(n802), .ZN(n805) );
  NAND2_X1 U896 ( .A1(n894), .A2(G105), .ZN(n803) );
  XOR2_X1 U897 ( .A(KEYINPUT38), .B(n803), .Z(n804) );
  NOR2_X1 U898 ( .A1(n805), .A2(n804), .ZN(n807) );
  NAND2_X1 U899 ( .A1(n893), .A2(G141), .ZN(n806) );
  NAND2_X1 U900 ( .A1(n807), .A2(n806), .ZN(n883) );
  NAND2_X1 U901 ( .A1(n883), .A2(G1996), .ZN(n816) );
  NAND2_X1 U902 ( .A1(G131), .A2(n893), .ZN(n809) );
  NAND2_X1 U903 ( .A1(G95), .A2(n894), .ZN(n808) );
  NAND2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n812) );
  NAND2_X1 U905 ( .A1(G119), .A2(n897), .ZN(n810) );
  XNOR2_X1 U906 ( .A(KEYINPUT91), .B(n810), .ZN(n811) );
  NOR2_X1 U907 ( .A1(n812), .A2(n811), .ZN(n814) );
  NAND2_X1 U908 ( .A1(n898), .A2(G107), .ZN(n813) );
  NAND2_X1 U909 ( .A1(n814), .A2(n813), .ZN(n878) );
  NAND2_X1 U910 ( .A1(n878), .A2(G1991), .ZN(n815) );
  NAND2_X1 U911 ( .A1(n816), .A2(n815), .ZN(n930) );
  NAND2_X1 U912 ( .A1(n930), .A2(n834), .ZN(n823) );
  NAND2_X1 U913 ( .A1(n831), .A2(n823), .ZN(n817) );
  XNOR2_X1 U914 ( .A(G1986), .B(G290), .ZN(n977) );
  NAND2_X1 U915 ( .A1(n977), .A2(n834), .ZN(n819) );
  NAND2_X1 U916 ( .A1(n820), .A2(n819), .ZN(n837) );
  AND2_X1 U917 ( .A1(n821), .A2(n905), .ZN(n822) );
  XNOR2_X1 U918 ( .A(n822), .B(KEYINPUT105), .ZN(n944) );
  NOR2_X1 U919 ( .A1(G1996), .A2(n883), .ZN(n932) );
  INV_X1 U920 ( .A(n823), .ZN(n826) );
  NOR2_X1 U921 ( .A1(G1986), .A2(G290), .ZN(n824) );
  NOR2_X1 U922 ( .A1(G1991), .A2(n878), .ZN(n925) );
  NOR2_X1 U923 ( .A1(n824), .A2(n925), .ZN(n825) );
  NOR2_X1 U924 ( .A1(n826), .A2(n825), .ZN(n827) );
  XOR2_X1 U925 ( .A(KEYINPUT103), .B(n827), .Z(n828) );
  NOR2_X1 U926 ( .A1(n932), .A2(n828), .ZN(n829) );
  XNOR2_X1 U927 ( .A(KEYINPUT104), .B(n829), .ZN(n830) );
  XNOR2_X1 U928 ( .A(n830), .B(KEYINPUT39), .ZN(n832) );
  NAND2_X1 U929 ( .A1(n832), .A2(n831), .ZN(n833) );
  NAND2_X1 U930 ( .A1(n944), .A2(n833), .ZN(n835) );
  NAND2_X1 U931 ( .A1(n835), .A2(n834), .ZN(n836) );
  NAND2_X1 U932 ( .A1(n837), .A2(n836), .ZN(n838) );
  XNOR2_X1 U933 ( .A(n838), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n922), .ZN(G217) );
  AND2_X1 U935 ( .A1(G15), .A2(G2), .ZN(n839) );
  NAND2_X1 U936 ( .A1(G661), .A2(n839), .ZN(G259) );
  NAND2_X1 U937 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U938 ( .A1(n841), .A2(n840), .ZN(G188) );
  XNOR2_X1 U939 ( .A(G108), .B(KEYINPUT119), .ZN(G238) );
  INV_X1 U941 ( .A(G120), .ZN(G236) );
  INV_X1 U942 ( .A(G96), .ZN(G221) );
  INV_X1 U943 ( .A(G69), .ZN(G235) );
  NOR2_X1 U944 ( .A1(n843), .A2(n842), .ZN(G325) );
  INV_X1 U945 ( .A(G325), .ZN(G261) );
  XOR2_X1 U946 ( .A(G1976), .B(G1971), .Z(n845) );
  XNOR2_X1 U947 ( .A(G1966), .B(G1956), .ZN(n844) );
  XNOR2_X1 U948 ( .A(n845), .B(n844), .ZN(n855) );
  XOR2_X1 U949 ( .A(G2474), .B(KEYINPUT41), .Z(n847) );
  XNOR2_X1 U950 ( .A(G1991), .B(KEYINPUT110), .ZN(n846) );
  XNOR2_X1 U951 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U952 ( .A(G1961), .B(G1981), .Z(n849) );
  XNOR2_X1 U953 ( .A(G1996), .B(G1986), .ZN(n848) );
  XNOR2_X1 U954 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U955 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U956 ( .A(KEYINPUT111), .B(KEYINPUT109), .ZN(n852) );
  XNOR2_X1 U957 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U958 ( .A(n855), .B(n854), .Z(G229) );
  XNOR2_X1 U959 ( .A(n856), .B(G2678), .ZN(n858) );
  XNOR2_X1 U960 ( .A(KEYINPUT42), .B(KEYINPUT107), .ZN(n857) );
  XNOR2_X1 U961 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U962 ( .A(KEYINPUT108), .B(G2072), .Z(n860) );
  XNOR2_X1 U963 ( .A(G2067), .B(G2090), .ZN(n859) );
  XNOR2_X1 U964 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U965 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U966 ( .A(KEYINPUT43), .B(G2096), .ZN(n863) );
  XNOR2_X1 U967 ( .A(n864), .B(n863), .ZN(n866) );
  XOR2_X1 U968 ( .A(G2078), .B(G2084), .Z(n865) );
  XNOR2_X1 U969 ( .A(n866), .B(n865), .ZN(G227) );
  NAND2_X1 U970 ( .A1(G124), .A2(n897), .ZN(n867) );
  XNOR2_X1 U971 ( .A(n867), .B(KEYINPUT112), .ZN(n868) );
  XNOR2_X1 U972 ( .A(n868), .B(KEYINPUT44), .ZN(n870) );
  NAND2_X1 U973 ( .A1(G100), .A2(n894), .ZN(n869) );
  NAND2_X1 U974 ( .A1(n870), .A2(n869), .ZN(n874) );
  NAND2_X1 U975 ( .A1(G136), .A2(n893), .ZN(n872) );
  NAND2_X1 U976 ( .A1(G112), .A2(n898), .ZN(n871) );
  NAND2_X1 U977 ( .A1(n872), .A2(n871), .ZN(n873) );
  NOR2_X1 U978 ( .A1(n874), .A2(n873), .ZN(G162) );
  XOR2_X1 U979 ( .A(KEYINPUT113), .B(KEYINPUT115), .Z(n876) );
  XNOR2_X1 U980 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n875) );
  XNOR2_X1 U981 ( .A(n876), .B(n875), .ZN(n877) );
  XNOR2_X1 U982 ( .A(G162), .B(n877), .ZN(n880) );
  XNOR2_X1 U983 ( .A(n878), .B(n924), .ZN(n879) );
  XNOR2_X1 U984 ( .A(n880), .B(n879), .ZN(n881) );
  XOR2_X1 U985 ( .A(G160), .B(n881), .Z(n882) );
  XNOR2_X1 U986 ( .A(n883), .B(n882), .ZN(n892) );
  NAND2_X1 U987 ( .A1(G130), .A2(n897), .ZN(n885) );
  NAND2_X1 U988 ( .A1(G118), .A2(n898), .ZN(n884) );
  NAND2_X1 U989 ( .A1(n885), .A2(n884), .ZN(n890) );
  NAND2_X1 U990 ( .A1(G142), .A2(n893), .ZN(n887) );
  NAND2_X1 U991 ( .A1(G106), .A2(n894), .ZN(n886) );
  NAND2_X1 U992 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U993 ( .A(KEYINPUT45), .B(n888), .Z(n889) );
  NOR2_X1 U994 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U995 ( .A(n892), .B(n891), .Z(n907) );
  NAND2_X1 U996 ( .A1(G139), .A2(n893), .ZN(n896) );
  NAND2_X1 U997 ( .A1(G103), .A2(n894), .ZN(n895) );
  NAND2_X1 U998 ( .A1(n896), .A2(n895), .ZN(n903) );
  NAND2_X1 U999 ( .A1(G127), .A2(n897), .ZN(n900) );
  NAND2_X1 U1000 ( .A1(G115), .A2(n898), .ZN(n899) );
  NAND2_X1 U1001 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U1002 ( .A(KEYINPUT47), .B(n901), .Z(n902) );
  NOR2_X1 U1003 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1004 ( .A(KEYINPUT114), .B(n904), .Z(n940) );
  XOR2_X1 U1005 ( .A(n905), .B(n940), .Z(n906) );
  XNOR2_X1 U1006 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1007 ( .A(G164), .B(n908), .Z(n909) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n909), .ZN(G395) );
  XOR2_X1 U1009 ( .A(G286), .B(KEYINPUT116), .Z(n910) );
  XOR2_X1 U1010 ( .A(n975), .B(n910), .Z(n913) );
  XNOR2_X1 U1011 ( .A(G171), .B(n911), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(n913), .B(n912), .ZN(n914) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n914), .ZN(G397) );
  NOR2_X1 U1014 ( .A1(G229), .A2(G227), .ZN(n916) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(KEYINPUT117), .ZN(n915) );
  XNOR2_X1 U1016 ( .A(n916), .B(n915), .ZN(n917) );
  NAND2_X1 U1017 ( .A1(G319), .A2(n917), .ZN(n918) );
  NOR2_X1 U1018 ( .A1(G401), .A2(n918), .ZN(n919) );
  XNOR2_X1 U1019 ( .A(KEYINPUT118), .B(n919), .ZN(n921) );
  NOR2_X1 U1020 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1022 ( .A(G225), .ZN(G308) );
  INV_X1 U1023 ( .A(n922), .ZN(G223) );
  XOR2_X1 U1024 ( .A(G160), .B(G2084), .Z(n923) );
  XNOR2_X1 U1025 ( .A(KEYINPUT120), .B(n923), .ZN(n928) );
  NOR2_X1 U1026 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1027 ( .A(n926), .B(KEYINPUT121), .ZN(n927) );
  NOR2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1029 ( .A(KEYINPUT122), .B(n929), .ZN(n939) );
  INV_X1 U1030 ( .A(n930), .ZN(n935) );
  XOR2_X1 U1031 ( .A(G2090), .B(G162), .Z(n931) );
  NOR2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1033 ( .A(KEYINPUT51), .B(n933), .Z(n934) );
  NAND2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n947) );
  XOR2_X1 U1037 ( .A(G164), .B(G2078), .Z(n942) );
  XNOR2_X1 U1038 ( .A(G2072), .B(n940), .ZN(n941) );
  NOR2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1040 ( .A(n943), .B(KEYINPUT50), .ZN(n945) );
  NAND2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(KEYINPUT52), .B(n948), .ZN(n950) );
  INV_X1 U1044 ( .A(KEYINPUT55), .ZN(n949) );
  NAND2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1046 ( .A1(n951), .A2(G29), .ZN(n973) );
  XNOR2_X1 U1047 ( .A(G1991), .B(G25), .ZN(n962) );
  XOR2_X1 U1048 ( .A(G32), .B(n952), .Z(n956) );
  XNOR2_X1 U1049 ( .A(G2067), .B(G26), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(G33), .B(G2072), .ZN(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n959) );
  XOR2_X1 U1053 ( .A(G27), .B(n957), .Z(n958) );
  NOR2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(KEYINPUT123), .B(n960), .ZN(n961) );
  NOR2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1057 ( .A1(G28), .A2(n963), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(n964), .B(KEYINPUT53), .ZN(n967) );
  XOR2_X1 U1059 ( .A(G2084), .B(G34), .Z(n965) );
  XNOR2_X1 U1060 ( .A(KEYINPUT54), .B(n965), .ZN(n966) );
  NAND2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(G35), .B(G2090), .ZN(n968) );
  NOR2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n1027) );
  INV_X1 U1064 ( .A(n1027), .ZN(n971) );
  NOR2_X1 U1065 ( .A1(G29), .A2(KEYINPUT55), .ZN(n970) );
  NAND2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n1000) );
  XOR2_X1 U1068 ( .A(G16), .B(KEYINPUT56), .Z(n998) );
  XOR2_X1 U1069 ( .A(G1956), .B(G299), .Z(n974) );
  XNOR2_X1 U1070 ( .A(n974), .B(KEYINPUT124), .ZN(n979) );
  XOR2_X1 U1071 ( .A(G1348), .B(n975), .Z(n976) );
  NOR2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n996) );
  XNOR2_X1 U1074 ( .A(G1966), .B(G168), .ZN(n981) );
  NAND2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(n982), .B(KEYINPUT57), .ZN(n994) );
  XOR2_X1 U1077 ( .A(G1341), .B(n983), .Z(n990) );
  AND2_X1 U1078 ( .A1(G303), .A2(G1971), .ZN(n987) );
  NAND2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1081 ( .A(KEYINPUT125), .B(n988), .Z(n989) );
  NAND2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n992) );
  XOR2_X1 U1083 ( .A(G171), .B(G1961), .Z(n991) );
  NOR2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1032) );
  XOR2_X1 U1089 ( .A(KEYINPUT58), .B(KEYINPUT127), .Z(n1007) );
  XNOR2_X1 U1090 ( .A(G1986), .B(G24), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(G1971), .B(G22), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XOR2_X1 U1093 ( .A(G1976), .B(KEYINPUT126), .Z(n1003) );
  XNOR2_X1 U1094 ( .A(G23), .B(n1003), .ZN(n1004) );
  NAND2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1096 ( .A(n1007), .B(n1006), .ZN(n1024) );
  XNOR2_X1 U1097 ( .A(G5), .B(n1008), .ZN(n1022) );
  XNOR2_X1 U1098 ( .A(G20), .B(n1009), .ZN(n1014) );
  XNOR2_X1 U1099 ( .A(G1981), .B(G6), .ZN(n1012) );
  XOR2_X1 U1100 ( .A(n1010), .B(G19), .Z(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1017) );
  XOR2_X1 U1103 ( .A(KEYINPUT59), .B(G1348), .Z(n1015) );
  XNOR2_X1 U1104 ( .A(G4), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1106 ( .A(KEYINPUT60), .B(n1018), .Z(n1020) );
  XNOR2_X1 U1107 ( .A(G1966), .B(G21), .ZN(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1111 ( .A(KEYINPUT61), .B(n1025), .Z(n1026) );
  NOR2_X1 U1112 ( .A1(G16), .A2(n1026), .ZN(n1030) );
  NAND2_X1 U1113 ( .A1(KEYINPUT55), .A2(n1027), .ZN(n1028) );
  NAND2_X1 U1114 ( .A1(G11), .A2(n1028), .ZN(n1029) );
  NOR2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1117 ( .A(KEYINPUT62), .B(n1033), .ZN(G150) );
  INV_X1 U1118 ( .A(G150), .ZN(G311) );
endmodule

