

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588;

  XOR2_X1 U325 ( .A(n299), .B(n347), .Z(n293) );
  XOR2_X1 U326 ( .A(G57GAT), .B(KEYINPUT72), .Z(n294) );
  XNOR2_X1 U327 ( .A(n344), .B(KEYINPUT73), .ZN(n345) );
  XNOR2_X1 U328 ( .A(KEYINPUT117), .B(KEYINPUT48), .ZN(n384) );
  XNOR2_X1 U329 ( .A(n346), .B(n345), .ZN(n349) );
  INV_X1 U330 ( .A(KEYINPUT10), .ZN(n303) );
  XNOR2_X1 U331 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U332 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U333 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U334 ( .A(n306), .B(n305), .ZN(n311) );
  XNOR2_X1 U335 ( .A(n448), .B(G190GAT), .ZN(n449) );
  XNOR2_X1 U336 ( .A(n450), .B(n449), .ZN(G1351GAT) );
  XOR2_X1 U337 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n296) );
  NAND2_X1 U338 ( .A1(G232GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U339 ( .A(n296), .B(n295), .ZN(n299) );
  XOR2_X1 U340 ( .A(G85GAT), .B(KEYINPUT74), .Z(n298) );
  XNOR2_X1 U341 ( .A(G99GAT), .B(G106GAT), .ZN(n297) );
  XNOR2_X1 U342 ( .A(n298), .B(n297), .ZN(n347) );
  XOR2_X1 U343 ( .A(G92GAT), .B(G218GAT), .Z(n301) );
  XNOR2_X1 U344 ( .A(G36GAT), .B(G190GAT), .ZN(n300) );
  XNOR2_X1 U345 ( .A(n301), .B(n300), .ZN(n316) );
  XNOR2_X1 U346 ( .A(G134GAT), .B(n316), .ZN(n302) );
  XNOR2_X1 U347 ( .A(n293), .B(n302), .ZN(n306) );
  XOR2_X1 U348 ( .A(G50GAT), .B(G162GAT), .Z(n392) );
  XNOR2_X1 U349 ( .A(n392), .B(KEYINPUT65), .ZN(n304) );
  XOR2_X1 U350 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n308) );
  XNOR2_X1 U351 ( .A(G43GAT), .B(G29GAT), .ZN(n307) );
  XNOR2_X1 U352 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U353 ( .A(KEYINPUT70), .B(n309), .Z(n338) );
  INV_X1 U354 ( .A(n338), .ZN(n310) );
  XOR2_X1 U355 ( .A(n311), .B(n310), .Z(n563) );
  XNOR2_X1 U356 ( .A(KEYINPUT76), .B(n563), .ZN(n548) );
  XOR2_X1 U357 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n313) );
  XNOR2_X1 U358 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n312) );
  XNOR2_X1 U359 ( .A(n313), .B(n312), .ZN(n442) );
  XOR2_X1 U360 ( .A(G204GAT), .B(G211GAT), .Z(n315) );
  XNOR2_X1 U361 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n314) );
  XNOR2_X1 U362 ( .A(n315), .B(n314), .ZN(n393) );
  XNOR2_X1 U363 ( .A(n442), .B(n393), .ZN(n322) );
  XOR2_X1 U364 ( .A(G8GAT), .B(G183GAT), .Z(n367) );
  XOR2_X1 U365 ( .A(G176GAT), .B(G64GAT), .Z(n351) );
  XNOR2_X1 U366 ( .A(n367), .B(n351), .ZN(n320) );
  XOR2_X1 U367 ( .A(KEYINPUT92), .B(n316), .Z(n318) );
  NAND2_X1 U368 ( .A1(G226GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U370 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n527) );
  XOR2_X1 U372 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n324) );
  XNOR2_X1 U373 ( .A(KEYINPUT67), .B(KEYINPUT29), .ZN(n323) );
  XNOR2_X1 U374 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U375 ( .A(G50GAT), .B(G36GAT), .Z(n326) );
  XOR2_X1 U376 ( .A(G113GAT), .B(G1GAT), .Z(n413) );
  XNOR2_X1 U377 ( .A(n413), .B(KEYINPUT66), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U379 ( .A(n328), .B(n327), .Z(n330) );
  NAND2_X1 U380 ( .A1(G229GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U381 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U382 ( .A(G197GAT), .B(G141GAT), .Z(n332) );
  XNOR2_X1 U383 ( .A(G169GAT), .B(G15GAT), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U385 ( .A(n334), .B(n333), .Z(n340) );
  XOR2_X1 U386 ( .A(KEYINPUT69), .B(KEYINPUT71), .Z(n336) );
  XNOR2_X1 U387 ( .A(G22GAT), .B(G8GAT), .ZN(n335) );
  XNOR2_X1 U388 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U389 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U390 ( .A(n340), .B(n339), .ZN(n576) );
  XNOR2_X1 U391 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n356) );
  XOR2_X1 U392 ( .A(KEYINPUT75), .B(KEYINPUT32), .Z(n342) );
  XNOR2_X1 U393 ( .A(G204GAT), .B(KEYINPUT31), .ZN(n341) );
  XNOR2_X1 U394 ( .A(n342), .B(n341), .ZN(n355) );
  XNOR2_X1 U395 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n343) );
  XNOR2_X1 U396 ( .A(n294), .B(n343), .ZN(n364) );
  XOR2_X1 U397 ( .A(G148GAT), .B(G78GAT), .Z(n390) );
  XNOR2_X1 U398 ( .A(n364), .B(n390), .ZN(n346) );
  AND2_X1 U399 ( .A1(G230GAT), .A2(G233GAT), .ZN(n344) );
  XOR2_X1 U400 ( .A(n347), .B(KEYINPUT33), .Z(n348) );
  XNOR2_X1 U401 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U402 ( .A(G120GAT), .B(G92GAT), .Z(n350) );
  XNOR2_X1 U403 ( .A(n355), .B(n354), .ZN(n580) );
  XNOR2_X1 U404 ( .A(n356), .B(n580), .ZN(n566) );
  NOR2_X1 U405 ( .A1(n576), .A2(n566), .ZN(n357) );
  XNOR2_X1 U406 ( .A(n357), .B(KEYINPUT46), .ZN(n373) );
  XOR2_X1 U407 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n359) );
  NAND2_X1 U408 ( .A1(G231GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U409 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U410 ( .A(KEYINPUT77), .B(n360), .ZN(n372) );
  XOR2_X1 U411 ( .A(KEYINPUT78), .B(G64GAT), .Z(n362) );
  XNOR2_X1 U412 ( .A(G1GAT), .B(KEYINPUT15), .ZN(n361) );
  XNOR2_X1 U413 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U414 ( .A(n364), .B(n363), .Z(n366) );
  XOR2_X1 U415 ( .A(G15GAT), .B(G127GAT), .Z(n432) );
  XOR2_X1 U416 ( .A(G22GAT), .B(G155GAT), .Z(n391) );
  XNOR2_X1 U417 ( .A(n432), .B(n391), .ZN(n365) );
  XNOR2_X1 U418 ( .A(n366), .B(n365), .ZN(n368) );
  XOR2_X1 U419 ( .A(n368), .B(n367), .Z(n370) );
  XNOR2_X1 U420 ( .A(G78GAT), .B(G211GAT), .ZN(n369) );
  XNOR2_X1 U421 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U422 ( .A(n372), .B(n371), .ZN(n583) );
  NOR2_X1 U423 ( .A1(n373), .A2(n583), .ZN(n374) );
  XNOR2_X1 U424 ( .A(n374), .B(KEYINPUT115), .ZN(n376) );
  INV_X1 U425 ( .A(n563), .ZN(n375) );
  NOR2_X1 U426 ( .A1(n376), .A2(n375), .ZN(n377) );
  XNOR2_X1 U427 ( .A(n377), .B(KEYINPUT47), .ZN(n383) );
  INV_X1 U428 ( .A(n583), .ZN(n559) );
  XNOR2_X1 U429 ( .A(KEYINPUT36), .B(n548), .ZN(n483) );
  NOR2_X1 U430 ( .A1(n559), .A2(n483), .ZN(n378) );
  XNOR2_X1 U431 ( .A(KEYINPUT45), .B(n378), .ZN(n379) );
  NAND2_X1 U432 ( .A1(n379), .A2(n576), .ZN(n380) );
  NOR2_X1 U433 ( .A1(n580), .A2(n380), .ZN(n381) );
  XOR2_X1 U434 ( .A(KEYINPUT116), .B(n381), .Z(n382) );
  AND2_X1 U435 ( .A1(n383), .A2(n382), .ZN(n385) );
  XNOR2_X1 U436 ( .A(n385), .B(n384), .ZN(n536) );
  NAND2_X1 U437 ( .A1(n527), .A2(n536), .ZN(n387) );
  XNOR2_X1 U438 ( .A(KEYINPUT123), .B(KEYINPUT54), .ZN(n386) );
  XNOR2_X1 U439 ( .A(n387), .B(n386), .ZN(n573) );
  XOR2_X1 U440 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n389) );
  XNOR2_X1 U441 ( .A(G218GAT), .B(G106GAT), .ZN(n388) );
  XNOR2_X1 U442 ( .A(n389), .B(n388), .ZN(n404) );
  XNOR2_X1 U443 ( .A(n391), .B(n390), .ZN(n402) );
  XOR2_X1 U444 ( .A(n393), .B(n392), .Z(n395) );
  NAND2_X1 U445 ( .A1(G228GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U446 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U447 ( .A(n396), .B(KEYINPUT88), .Z(n400) );
  XOR2_X1 U448 ( .A(KEYINPUT3), .B(KEYINPUT87), .Z(n398) );
  XNOR2_X1 U449 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n397) );
  XNOR2_X1 U450 ( .A(n398), .B(n397), .ZN(n414) );
  XNOR2_X1 U451 ( .A(n414), .B(KEYINPUT22), .ZN(n399) );
  XNOR2_X1 U452 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U453 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U454 ( .A(n404), .B(n403), .ZN(n462) );
  XOR2_X1 U455 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n406) );
  XNOR2_X1 U456 ( .A(KEYINPUT6), .B(KEYINPUT89), .ZN(n405) );
  XNOR2_X1 U457 ( .A(n406), .B(n405), .ZN(n425) );
  XOR2_X1 U458 ( .A(KEYINPUT1), .B(G57GAT), .Z(n408) );
  XNOR2_X1 U459 ( .A(G155GAT), .B(G148GAT), .ZN(n407) );
  XNOR2_X1 U460 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U461 ( .A(G85GAT), .B(G162GAT), .Z(n410) );
  XNOR2_X1 U462 ( .A(G29GAT), .B(G127GAT), .ZN(n409) );
  XNOR2_X1 U463 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U464 ( .A(n412), .B(n411), .ZN(n423) );
  XOR2_X1 U465 ( .A(n414), .B(n413), .Z(n416) );
  NAND2_X1 U466 ( .A1(G225GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U467 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U468 ( .A(n417), .B(KEYINPUT5), .Z(n421) );
  XOR2_X1 U469 ( .A(G120GAT), .B(KEYINPUT0), .Z(n419) );
  XNOR2_X1 U470 ( .A(G134GAT), .B(KEYINPUT81), .ZN(n418) );
  XNOR2_X1 U471 ( .A(n419), .B(n418), .ZN(n441) );
  XNOR2_X1 U472 ( .A(n441), .B(KEYINPUT4), .ZN(n420) );
  XNOR2_X1 U473 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U474 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U475 ( .A(n425), .B(n424), .ZN(n524) );
  INV_X1 U476 ( .A(n524), .ZN(n572) );
  AND2_X1 U477 ( .A1(n462), .A2(n572), .ZN(n426) );
  NAND2_X1 U478 ( .A1(n573), .A2(n426), .ZN(n427) );
  XNOR2_X1 U479 ( .A(n427), .B(KEYINPUT55), .ZN(n447) );
  XOR2_X1 U480 ( .A(G183GAT), .B(KEYINPUT86), .Z(n429) );
  XNOR2_X1 U481 ( .A(KEYINPUT83), .B(KEYINPUT85), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n429), .B(n428), .ZN(n437) );
  XOR2_X1 U483 ( .A(KEYINPUT82), .B(G71GAT), .Z(n431) );
  XNOR2_X1 U484 ( .A(G190GAT), .B(G99GAT), .ZN(n430) );
  XNOR2_X1 U485 ( .A(n431), .B(n430), .ZN(n433) );
  XOR2_X1 U486 ( .A(n433), .B(n432), .Z(n435) );
  XNOR2_X1 U487 ( .A(G43GAT), .B(G113GAT), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U489 ( .A(n437), .B(n436), .ZN(n446) );
  XOR2_X1 U490 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n439) );
  NAND2_X1 U491 ( .A1(G227GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U493 ( .A(n440), .B(G176GAT), .Z(n444) );
  XNOR2_X1 U494 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U495 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U496 ( .A(n446), .B(n445), .ZN(n538) );
  NAND2_X1 U497 ( .A1(n447), .A2(n538), .ZN(n451) );
  NOR2_X1 U498 ( .A1(n548), .A2(n451), .ZN(n450) );
  XNOR2_X1 U499 ( .A(KEYINPUT127), .B(KEYINPUT58), .ZN(n448) );
  NOR2_X1 U500 ( .A1(n559), .A2(n451), .ZN(n454) );
  INV_X1 U501 ( .A(G183GAT), .ZN(n452) );
  XNOR2_X1 U502 ( .A(n452), .B(KEYINPUT126), .ZN(n453) );
  XNOR2_X1 U503 ( .A(n454), .B(n453), .ZN(G1350GAT) );
  NOR2_X1 U504 ( .A1(n576), .A2(n580), .ZN(n488) );
  NAND2_X1 U505 ( .A1(n583), .A2(n548), .ZN(n457) );
  XNOR2_X1 U506 ( .A(KEYINPUT16), .B(KEYINPUT80), .ZN(n455) );
  XNOR2_X1 U507 ( .A(n455), .B(KEYINPUT79), .ZN(n456) );
  XNOR2_X1 U508 ( .A(n457), .B(n456), .ZN(n469) );
  NAND2_X1 U509 ( .A1(n538), .A2(n527), .ZN(n458) );
  NAND2_X1 U510 ( .A1(n462), .A2(n458), .ZN(n459) );
  XNOR2_X1 U511 ( .A(n459), .B(KEYINPUT25), .ZN(n460) );
  NAND2_X1 U512 ( .A1(n460), .A2(n572), .ZN(n468) );
  INV_X1 U513 ( .A(n538), .ZN(n499) );
  XOR2_X1 U514 ( .A(KEYINPUT28), .B(n462), .Z(n537) );
  INV_X1 U515 ( .A(n537), .ZN(n503) );
  NAND2_X1 U516 ( .A1(n499), .A2(n503), .ZN(n461) );
  NAND2_X1 U517 ( .A1(n461), .A2(n524), .ZN(n466) );
  XOR2_X1 U518 ( .A(n527), .B(KEYINPUT27), .Z(n534) );
  NOR2_X1 U519 ( .A1(n462), .A2(n538), .ZN(n463) );
  XNOR2_X1 U520 ( .A(n463), .B(KEYINPUT26), .ZN(n574) );
  NOR2_X1 U521 ( .A1(n574), .A2(n524), .ZN(n464) );
  NOR2_X1 U522 ( .A1(n534), .A2(n464), .ZN(n465) );
  NAND2_X1 U523 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U524 ( .A1(n468), .A2(n467), .ZN(n484) );
  NAND2_X1 U525 ( .A1(n469), .A2(n484), .ZN(n470) );
  XNOR2_X1 U526 ( .A(KEYINPUT93), .B(n470), .ZN(n507) );
  NAND2_X1 U527 ( .A1(n488), .A2(n507), .ZN(n479) );
  NOR2_X1 U528 ( .A1(n572), .A2(n479), .ZN(n472) );
  XNOR2_X1 U529 ( .A(KEYINPUT94), .B(KEYINPUT34), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U531 ( .A(G1GAT), .B(n473), .Z(G1324GAT) );
  INV_X1 U532 ( .A(n527), .ZN(n496) );
  NOR2_X1 U533 ( .A1(n496), .A2(n479), .ZN(n475) );
  XNOR2_X1 U534 ( .A(KEYINPUT95), .B(KEYINPUT96), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U536 ( .A(G8GAT), .B(n476), .ZN(G1325GAT) );
  NOR2_X1 U537 ( .A1(n499), .A2(n479), .ZN(n478) );
  XNOR2_X1 U538 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n478), .B(n477), .ZN(G1326GAT) );
  NOR2_X1 U540 ( .A1(n503), .A2(n479), .ZN(n481) );
  XNOR2_X1 U541 ( .A(KEYINPUT97), .B(KEYINPUT98), .ZN(n480) );
  XNOR2_X1 U542 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U543 ( .A(G22GAT), .B(n482), .ZN(G1327GAT) );
  NAND2_X1 U544 ( .A1(n559), .A2(n484), .ZN(n485) );
  NOR2_X1 U545 ( .A1(n483), .A2(n485), .ZN(n487) );
  XOR2_X1 U546 ( .A(KEYINPUT100), .B(KEYINPUT37), .Z(n486) );
  XNOR2_X1 U547 ( .A(n487), .B(n486), .ZN(n522) );
  NAND2_X1 U548 ( .A1(n522), .A2(n488), .ZN(n491) );
  XOR2_X1 U549 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n489) );
  XNOR2_X1 U550 ( .A(KEYINPUT38), .B(n489), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(n502) );
  NOR2_X1 U552 ( .A1(n572), .A2(n502), .ZN(n495) );
  XNOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n492), .B(KEYINPUT103), .ZN(n493) );
  XNOR2_X1 U555 ( .A(KEYINPUT99), .B(n493), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(G1328GAT) );
  NOR2_X1 U557 ( .A1(n496), .A2(n502), .ZN(n497) );
  XOR2_X1 U558 ( .A(G36GAT), .B(n497), .Z(n498) );
  XNOR2_X1 U559 ( .A(KEYINPUT104), .B(n498), .ZN(G1329GAT) );
  NOR2_X1 U560 ( .A1(n499), .A2(n502), .ZN(n500) );
  XOR2_X1 U561 ( .A(KEYINPUT40), .B(n500), .Z(n501) );
  XNOR2_X1 U562 ( .A(G43GAT), .B(n501), .ZN(G1330GAT) );
  NOR2_X1 U563 ( .A1(n503), .A2(n502), .ZN(n505) );
  XNOR2_X1 U564 ( .A(G50GAT), .B(KEYINPUT105), .ZN(n504) );
  XNOR2_X1 U565 ( .A(n505), .B(n504), .ZN(G1331GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT42), .B(KEYINPUT107), .Z(n510) );
  INV_X1 U567 ( .A(n576), .ZN(n506) );
  NOR2_X1 U568 ( .A1(n506), .A2(n566), .ZN(n521) );
  NAND2_X1 U569 ( .A1(n507), .A2(n521), .ZN(n508) );
  XOR2_X1 U570 ( .A(KEYINPUT106), .B(n508), .Z(n517) );
  NAND2_X1 U571 ( .A1(n517), .A2(n524), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(n511), .ZN(G1332GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n513) );
  NAND2_X1 U575 ( .A1(n527), .A2(n517), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U577 ( .A(G64GAT), .B(n514), .ZN(G1333GAT) );
  NAND2_X1 U578 ( .A1(n517), .A2(n538), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n515), .B(KEYINPUT110), .ZN(n516) );
  XNOR2_X1 U580 ( .A(G71GAT), .B(n516), .ZN(G1334GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U582 ( .A1(n517), .A2(n537), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U584 ( .A(G78GAT), .B(n520), .Z(G1335GAT) );
  XOR2_X1 U585 ( .A(G85GAT), .B(KEYINPUT113), .Z(n526) );
  NAND2_X1 U586 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U587 ( .A(KEYINPUT112), .B(n523), .Z(n530) );
  NAND2_X1 U588 ( .A1(n530), .A2(n524), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n526), .B(n525), .ZN(G1336GAT) );
  NAND2_X1 U590 ( .A1(n530), .A2(n527), .ZN(n528) );
  XNOR2_X1 U591 ( .A(n528), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U592 ( .A1(n530), .A2(n538), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n529), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT114), .B(KEYINPUT44), .Z(n532) );
  NAND2_X1 U595 ( .A1(n530), .A2(n537), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U597 ( .A(G106GAT), .B(n533), .Z(G1339GAT) );
  NOR2_X1 U598 ( .A1(n572), .A2(n534), .ZN(n535) );
  NAND2_X1 U599 ( .A1(n536), .A2(n535), .ZN(n551) );
  NOR2_X1 U600 ( .A1(n537), .A2(n551), .ZN(n539) );
  NAND2_X1 U601 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U602 ( .A(n540), .B(KEYINPUT118), .ZN(n547) );
  NOR2_X1 U603 ( .A1(n576), .A2(n547), .ZN(n541) );
  XOR2_X1 U604 ( .A(G113GAT), .B(n541), .Z(G1340GAT) );
  NOR2_X1 U605 ( .A1(n547), .A2(n566), .ZN(n543) );
  XNOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n543), .B(n542), .ZN(G1341GAT) );
  NOR2_X1 U608 ( .A1(n547), .A2(n559), .ZN(n545) );
  XNOR2_X1 U609 ( .A(KEYINPUT119), .B(KEYINPUT50), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  XNOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n550) );
  NOR2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  INV_X1 U615 ( .A(n551), .ZN(n552) );
  NAND2_X1 U616 ( .A1(n552), .A2(n574), .ZN(n562) );
  NOR2_X1 U617 ( .A1(n576), .A2(n562), .ZN(n553) );
  XOR2_X1 U618 ( .A(G141GAT), .B(n553), .Z(G1344GAT) );
  NOR2_X1 U619 ( .A1(n566), .A2(n562), .ZN(n558) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT121), .Z(n555) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(KEYINPUT120), .B(n556), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n562), .ZN(n560) );
  XOR2_X1 U626 ( .A(KEYINPUT122), .B(n560), .Z(n561) );
  XNOR2_X1 U627 ( .A(G155GAT), .B(n561), .ZN(G1346GAT) );
  NOR2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U629 ( .A(G162GAT), .B(n564), .Z(G1347GAT) );
  NOR2_X1 U630 ( .A1(n576), .A2(n451), .ZN(n565) );
  XOR2_X1 U631 ( .A(G169GAT), .B(n565), .Z(G1348GAT) );
  NOR2_X1 U632 ( .A1(n566), .A2(n451), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n568) );
  XNOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(KEYINPUT124), .B(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1349GAT) );
  AND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n586) );
  NOR2_X1 U640 ( .A1(n576), .A2(n586), .ZN(n578) );
  XNOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .Z(n582) );
  INV_X1 U645 ( .A(n586), .ZN(n584) );
  NAND2_X1 U646 ( .A1(n584), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NAND2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(n585), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U650 ( .A1(n483), .A2(n586), .ZN(n587) );
  XOR2_X1 U651 ( .A(KEYINPUT62), .B(n587), .Z(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

