

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775;

  OR2_X2 U379 ( .A1(n685), .A2(n688), .ZN(n721) );
  XNOR2_X2 U380 ( .A(KEYINPUT32), .B(n615), .ZN(n775) );
  XNOR2_X1 U381 ( .A(n355), .B(n465), .ZN(n464) );
  NAND2_X1 U382 ( .A1(n626), .A2(n627), .ZN(n355) );
  OR2_X2 U383 ( .A1(n389), .A2(n613), .ZN(n398) );
  XNOR2_X2 U384 ( .A(n440), .B(n439), .ZN(n389) );
  NOR2_X2 U385 ( .A1(n405), .A2(n399), .ZN(n358) );
  AND2_X2 U386 ( .A1(n448), .A2(n445), .ZN(n424) );
  XNOR2_X2 U387 ( .A(n523), .B(n373), .ZN(n667) );
  XNOR2_X2 U388 ( .A(n757), .B(G146), .ZN(n523) );
  NOR2_X2 U389 ( .A1(n427), .A2(n618), .ZN(n671) );
  NOR2_X1 U390 ( .A1(n583), .A2(n716), .ZN(n585) );
  XNOR2_X1 U391 ( .A(KEYINPUT1), .B(n569), .ZN(n706) );
  INV_X2 U392 ( .A(G143), .ZN(n426) );
  NAND2_X1 U393 ( .A1(n706), .A2(n705), .ZN(n619) );
  INV_X1 U394 ( .A(n703), .ZN(n356) );
  XNOR2_X1 U395 ( .A(n363), .B(n481), .ZN(n518) );
  INV_X1 U396 ( .A(KEYINPUT72), .ZN(n484) );
  NOR2_X1 U397 ( .A1(n405), .A2(n399), .ZN(n763) );
  OR2_X1 U398 ( .A1(n629), .A2(KEYINPUT44), .ZN(n630) );
  BUF_X1 U399 ( .A(n771), .Z(n387) );
  XNOR2_X1 U400 ( .A(n372), .B(n586), .ZN(n771) );
  XNOR2_X1 U401 ( .A(n422), .B(KEYINPUT79), .ZN(n571) );
  INV_X2 U402 ( .A(n623), .ZN(n357) );
  XNOR2_X1 U403 ( .A(n412), .B(n479), .ZN(n569) );
  XNOR2_X1 U404 ( .A(n428), .B(n539), .ZN(n703) );
  OR2_X1 U405 ( .A1(n740), .A2(G902), .ZN(n412) );
  XNOR2_X1 U406 ( .A(n432), .B(n374), .ZN(n373) );
  XNOR2_X1 U407 ( .A(n525), .B(n522), .ZN(n432) );
  XNOR2_X1 U408 ( .A(n519), .B(n518), .ZN(n374) );
  XNOR2_X1 U409 ( .A(n381), .B(KEYINPUT77), .ZN(n524) );
  XNOR2_X1 U410 ( .A(n491), .B(n490), .ZN(n548) );
  NOR2_X1 U411 ( .A1(n662), .A2(n634), .ZN(n491) );
  BUF_X1 U412 ( .A(n697), .Z(n359) );
  BUF_X1 U413 ( .A(n662), .Z(n360) );
  BUF_X1 U414 ( .A(n746), .Z(n750) );
  AND2_X1 U415 ( .A1(n580), .A2(n581), .ZN(n473) );
  INV_X1 U416 ( .A(KEYINPUT18), .ZN(n386) );
  XNOR2_X1 U417 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U418 ( .A(n480), .B(G469), .ZN(n479) );
  INV_X1 U419 ( .A(KEYINPUT71), .ZN(n480) );
  NAND2_X1 U420 ( .A1(n705), .A2(n433), .ZN(n621) );
  XOR2_X1 U421 ( .A(KEYINPUT8), .B(KEYINPUT70), .Z(n502) );
  NOR2_X1 U422 ( .A1(n702), .A2(n415), .ZN(n414) );
  OR2_X1 U423 ( .A1(G237), .A2(G902), .ZN(n492) );
  NAND2_X1 U424 ( .A1(n701), .A2(n382), .ZN(n381) );
  INV_X1 U425 ( .A(G237), .ZN(n382) );
  INV_X1 U426 ( .A(G137), .ZN(n420) );
  XNOR2_X1 U427 ( .A(n434), .B(G146), .ZN(n510) );
  INV_X1 U428 ( .A(G125), .ZN(n434) );
  XNOR2_X1 U429 ( .A(n512), .B(n379), .ZN(n513) );
  XNOR2_X1 U430 ( .A(KEYINPUT103), .B(KEYINPUT12), .ZN(n512) );
  XNOR2_X1 U431 ( .A(KEYINPUT11), .B(KEYINPUT102), .ZN(n379) );
  XOR2_X1 U432 ( .A(G122), .B(G104), .Z(n509) );
  XNOR2_X1 U433 ( .A(G143), .B(G113), .ZN(n508) );
  XNOR2_X1 U434 ( .A(n476), .B(G140), .ZN(n511) );
  INV_X1 U435 ( .A(G131), .ZN(n476) );
  INV_X1 U436 ( .A(n510), .ZN(n485) );
  INV_X1 U437 ( .A(n573), .ZN(n589) );
  NOR2_X1 U438 ( .A1(n752), .A2(G902), .ZN(n428) );
  XNOR2_X1 U439 ( .A(KEYINPUT67), .B(G101), .ZN(n477) );
  NAND2_X1 U440 ( .A1(n403), .A2(n400), .ZN(n399) );
  NOR2_X1 U441 ( .A1(n402), .A2(n401), .ZN(n400) );
  XNOR2_X1 U442 ( .A(n518), .B(n442), .ZN(n652) );
  XNOR2_X1 U443 ( .A(n482), .B(G122), .ZN(n442) );
  XOR2_X1 U444 ( .A(KEYINPUT75), .B(KEYINPUT16), .Z(n482) );
  XNOR2_X1 U445 ( .A(G128), .B(G119), .ZN(n459) );
  XNOR2_X1 U446 ( .A(n457), .B(n456), .ZN(n455) );
  XNOR2_X1 U447 ( .A(KEYINPUT24), .B(KEYINPUT97), .ZN(n457) );
  XNOR2_X1 U448 ( .A(G137), .B(KEYINPUT23), .ZN(n456) );
  XNOR2_X1 U449 ( .A(n510), .B(KEYINPUT10), .ZN(n532) );
  INV_X1 U450 ( .A(KEYINPUT91), .ZN(n549) );
  NOR2_X1 U451 ( .A1(n589), .A2(n588), .ZN(n605) );
  XNOR2_X1 U452 ( .A(n561), .B(n436), .ZN(n563) );
  XNOR2_X1 U453 ( .A(n437), .B(KEYINPUT28), .ZN(n436) );
  AND2_X1 U454 ( .A1(n450), .A2(n357), .ZN(n449) );
  NOR2_X1 U455 ( .A1(n621), .A2(KEYINPUT99), .ZN(n450) );
  INV_X1 U456 ( .A(KEYINPUT64), .ZN(n423) );
  XNOR2_X1 U457 ( .A(n529), .B(KEYINPUT20), .ZN(n535) );
  NOR2_X1 U458 ( .A1(n691), .A2(n555), .ZN(n581) );
  AND2_X1 U459 ( .A1(n380), .A2(KEYINPUT84), .ZN(n577) );
  INV_X1 U460 ( .A(KEYINPUT46), .ZN(n472) );
  NAND2_X1 U461 ( .A1(n771), .A2(n773), .ZN(n593) );
  INV_X1 U462 ( .A(KEYINPUT108), .ZN(n391) );
  NAND2_X1 U463 ( .A1(n362), .A2(n411), .ZN(n705) );
  XOR2_X1 U464 ( .A(KEYINPUT25), .B(KEYINPUT80), .Z(n537) );
  INV_X1 U465 ( .A(n693), .ZN(n401) );
  NOR2_X1 U466 ( .A1(n694), .A2(KEYINPUT88), .ZN(n404) );
  XNOR2_X1 U467 ( .A(n493), .B(KEYINPUT94), .ZN(n566) );
  INV_X1 U468 ( .A(KEYINPUT95), .ZN(n462) );
  XNOR2_X1 U469 ( .A(KEYINPUT30), .B(KEYINPUT111), .ZN(n567) );
  INV_X1 U470 ( .A(KEYINPUT113), .ZN(n437) );
  NOR2_X1 U471 ( .A1(n560), .A2(n559), .ZN(n561) );
  BUF_X1 U472 ( .A(n569), .Z(n433) );
  INV_X1 U473 ( .A(KEYINPUT22), .ZN(n439) );
  XNOR2_X1 U474 ( .A(G131), .B(KEYINPUT100), .ZN(n520) );
  XOR2_X1 U475 ( .A(KEYINPUT76), .B(KEYINPUT5), .Z(n521) );
  XNOR2_X1 U476 ( .A(G122), .B(KEYINPUT9), .ZN(n497) );
  XOR2_X1 U477 ( .A(KEYINPUT105), .B(KEYINPUT7), .Z(n498) );
  XNOR2_X1 U478 ( .A(G116), .B(G107), .ZN(n496) );
  XNOR2_X1 U479 ( .A(n435), .B(n755), .ZN(n638) );
  XNOR2_X1 U480 ( .A(n515), .B(n364), .ZN(n435) );
  XNOR2_X1 U481 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U482 ( .A(n495), .B(n475), .ZN(n474) );
  XNOR2_X1 U483 ( .A(n511), .B(KEYINPUT96), .ZN(n475) );
  XNOR2_X1 U484 ( .A(n383), .B(n393), .ZN(n662) );
  XNOR2_X1 U485 ( .A(n652), .B(n394), .ZN(n393) );
  XNOR2_X1 U486 ( .A(n388), .B(n384), .ZN(n383) );
  NAND2_X1 U487 ( .A1(G234), .A2(G237), .ZN(n528) );
  XNOR2_X1 U488 ( .A(n585), .B(n584), .ZN(n595) );
  XNOR2_X1 U489 ( .A(n378), .B(n376), .ZN(n573) );
  XNOR2_X1 U490 ( .A(n516), .B(n377), .ZN(n376) );
  OR2_X1 U491 ( .A1(n638), .A2(G902), .ZN(n378) );
  INV_X1 U492 ( .A(G475), .ZN(n377) );
  BUF_X1 U493 ( .A(n703), .Z(n427) );
  XNOR2_X1 U494 ( .A(n534), .B(n533), .ZN(n752) );
  XNOR2_X1 U495 ( .A(n454), .B(n532), .ZN(n533) );
  NOR2_X1 U496 ( .A1(n478), .A2(n631), .ZN(n635) );
  XOR2_X1 U497 ( .A(KEYINPUT92), .B(n641), .Z(n739) );
  XNOR2_X1 U498 ( .A(n606), .B(KEYINPUT35), .ZN(n467) );
  NOR2_X1 U499 ( .A1(n599), .A2(n587), .ZN(n682) );
  NAND2_X1 U500 ( .A1(n446), .A2(n357), .ZN(n447) );
  INV_X1 U501 ( .A(n694), .ZN(n470) );
  AND2_X1 U502 ( .A1(n570), .A2(n461), .ZN(n361) );
  NAND2_X1 U503 ( .A1(n407), .A2(n415), .ZN(n362) );
  XOR2_X1 U504 ( .A(G113), .B(G116), .Z(n363) );
  XOR2_X1 U505 ( .A(n509), .B(n508), .Z(n364) );
  AND2_X1 U506 ( .A1(n414), .A2(n361), .ZN(n365) );
  AND2_X1 U507 ( .A1(n361), .A2(n415), .ZN(n366) );
  NOR2_X1 U508 ( .A1(n452), .A2(n623), .ZN(n367) );
  NOR2_X1 U509 ( .A1(n608), .A2(n702), .ZN(n368) );
  INV_X1 U510 ( .A(n721), .ZN(n624) );
  INV_X1 U511 ( .A(n733), .ZN(n461) );
  XNOR2_X1 U512 ( .A(KEYINPUT66), .B(KEYINPUT0), .ZN(n369) );
  NAND2_X1 U513 ( .A1(n598), .A2(n461), .ZN(n370) );
  INV_X1 U514 ( .A(n631), .ZN(n634) );
  XOR2_X1 U515 ( .A(KEYINPUT86), .B(KEYINPUT2), .Z(n371) );
  INV_X1 U516 ( .A(KEYINPUT88), .ZN(n417) );
  NAND2_X1 U517 ( .A1(n595), .A2(n685), .ZN(n372) );
  XNOR2_X2 U518 ( .A(n756), .B(n477), .ZN(n519) );
  XNOR2_X2 U519 ( .A(n506), .B(n420), .ZN(n757) );
  XNOR2_X2 U520 ( .A(n494), .B(G134), .ZN(n506) );
  XNOR2_X2 U521 ( .A(n375), .B(n519), .ZN(n388) );
  XNOR2_X2 U522 ( .A(n650), .B(n484), .ZN(n375) );
  NAND2_X1 U523 ( .A1(n682), .A2(n721), .ZN(n380) );
  XNOR2_X1 U524 ( .A(n486), .B(n385), .ZN(n384) );
  XNOR2_X1 U525 ( .A(n494), .B(n386), .ZN(n385) );
  XNOR2_X1 U526 ( .A(n421), .B(n523), .ZN(n740) );
  BUF_X1 U527 ( .A(n548), .Z(n582) );
  XNOR2_X1 U528 ( .A(n460), .B(n459), .ZN(n458) );
  XNOR2_X1 U529 ( .A(n458), .B(n455), .ZN(n454) );
  XNOR2_X1 U530 ( .A(G140), .B(G110), .ZN(n460) );
  XNOR2_X1 U531 ( .A(n418), .B(n594), .ZN(n406) );
  NAND2_X1 U532 ( .A1(n444), .A2(n357), .ZN(n443) );
  NOR2_X1 U533 ( .A1(n406), .A2(n417), .ZN(n405) );
  NAND2_X1 U534 ( .A1(n406), .A2(n404), .ZN(n403) );
  BUF_X1 U535 ( .A(n772), .Z(n390) );
  XNOR2_X1 U536 ( .A(n392), .B(n391), .ZN(n625) );
  NAND2_X1 U537 ( .A1(n429), .A2(n721), .ZN(n392) );
  XNOR2_X1 U538 ( .A(n468), .B(n467), .ZN(n772) );
  XNOR2_X1 U539 ( .A(n425), .B(n620), .ZN(n689) );
  NAND2_X1 U540 ( .A1(n469), .A2(n605), .ZN(n468) );
  XNOR2_X1 U541 ( .A(n604), .B(n603), .ZN(n469) );
  XNOR2_X1 U542 ( .A(n388), .B(n474), .ZN(n421) );
  INV_X1 U543 ( .A(n622), .ZN(n451) );
  XNOR2_X1 U544 ( .A(n485), .B(n487), .ZN(n394) );
  NAND2_X1 U545 ( .A1(n712), .A2(n395), .ZN(n425) );
  AND2_X1 U546 ( .A1(n395), .A2(n368), .ZN(n440) );
  XNOR2_X1 U547 ( .A(n395), .B(n462), .ZN(n602) );
  XNOR2_X2 U548 ( .A(n419), .B(n369), .ZN(n395) );
  OR2_X1 U549 ( .A1(n389), .A2(n396), .ZN(n615) );
  NAND2_X1 U550 ( .A1(n614), .A2(n397), .ZN(n396) );
  INV_X1 U551 ( .A(n613), .ZN(n397) );
  XNOR2_X1 U552 ( .A(n398), .B(KEYINPUT89), .ZN(n431) );
  NOR2_X1 U553 ( .A1(n470), .A2(n417), .ZN(n402) );
  NAND2_X1 U554 ( .A1(n407), .A2(n366), .ZN(n409) );
  NAND2_X1 U555 ( .A1(n356), .A2(n607), .ZN(n407) );
  NAND2_X1 U556 ( .A1(n408), .A2(n569), .ZN(n422) );
  NAND2_X1 U557 ( .A1(n410), .A2(n409), .ZN(n408) );
  NAND2_X1 U558 ( .A1(n365), .A2(n356), .ZN(n410) );
  NAND2_X1 U559 ( .A1(n356), .A2(n414), .ZN(n411) );
  XNOR2_X2 U560 ( .A(n413), .B(n556), .ZN(n599) );
  NOR2_X1 U561 ( .A1(n413), .A2(n551), .ZN(n552) );
  XNOR2_X2 U562 ( .A(n416), .B(n549), .ZN(n413) );
  INV_X1 U563 ( .A(KEYINPUT68), .ZN(n415) );
  NAND2_X1 U564 ( .A1(n548), .A2(n566), .ZN(n416) );
  NAND2_X1 U565 ( .A1(n471), .A2(n473), .ZN(n418) );
  NOR2_X2 U566 ( .A1(n599), .A2(n370), .ZN(n419) );
  XNOR2_X1 U567 ( .A(n430), .B(KEYINPUT78), .ZN(n583) );
  XNOR2_X2 U568 ( .A(n423), .B(G953), .ZN(n767) );
  NAND2_X1 U569 ( .A1(n424), .A2(n443), .ZN(n429) );
  XNOR2_X2 U570 ( .A(n426), .B(G128), .ZN(n494) );
  NOR2_X1 U571 ( .A1(n772), .A2(n677), .ZN(n616) );
  XNOR2_X1 U572 ( .A(n568), .B(n567), .ZN(n572) );
  INV_X1 U573 ( .A(n453), .ZN(n444) );
  NAND2_X1 U574 ( .A1(n571), .A2(n572), .ZN(n430) );
  XNOR2_X1 U575 ( .A(n593), .B(n472), .ZN(n471) );
  NAND2_X1 U576 ( .A1(n431), .A2(n617), .ZN(n618) );
  NOR2_X2 U577 ( .A1(n667), .A2(G902), .ZN(n526) );
  XNOR2_X2 U578 ( .A(KEYINPUT15), .B(G902), .ZN(n631) );
  NAND2_X1 U579 ( .A1(n746), .A2(G210), .ZN(n663) );
  NAND2_X2 U580 ( .A1(n637), .A2(n636), .ZN(n746) );
  NAND2_X1 U581 ( .A1(n438), .A2(n739), .ZN(n670) );
  XNOR2_X1 U582 ( .A(n668), .B(n669), .ZN(n438) );
  XNOR2_X2 U583 ( .A(G104), .B(G110), .ZN(n483) );
  NAND2_X1 U584 ( .A1(n441), .A2(n739), .ZN(n666) );
  XNOR2_X1 U585 ( .A(n663), .B(n664), .ZN(n441) );
  XNOR2_X2 U586 ( .A(n526), .B(n527), .ZN(n558) );
  NAND2_X1 U587 ( .A1(n451), .A2(n449), .ZN(n448) );
  NOR2_X1 U588 ( .A1(n689), .A2(n367), .ZN(n445) );
  NAND2_X1 U589 ( .A1(n453), .A2(n452), .ZN(n446) );
  NAND2_X1 U590 ( .A1(n447), .A2(n448), .ZN(n673) );
  NAND2_X1 U591 ( .A1(n621), .A2(KEYINPUT99), .ZN(n452) );
  NAND2_X1 U592 ( .A1(n622), .A2(KEYINPUT99), .ZN(n453) );
  NOR2_X1 U593 ( .A1(KEYINPUT47), .A2(n577), .ZN(n578) );
  XNOR2_X2 U594 ( .A(n558), .B(n557), .ZN(n609) );
  INV_X1 U595 ( .A(n602), .ZN(n622) );
  NAND2_X1 U596 ( .A1(n466), .A2(n697), .ZN(n695) );
  XNOR2_X2 U597 ( .A(n463), .B(KEYINPUT45), .ZN(n697) );
  NAND2_X1 U598 ( .A1(n464), .A2(n630), .ZN(n463) );
  INV_X1 U599 ( .A(KEYINPUT90), .ZN(n465) );
  XNOR2_X1 U600 ( .A(n763), .B(KEYINPUT86), .ZN(n466) );
  XNOR2_X2 U601 ( .A(n483), .B(G107), .ZN(n650) );
  INV_X1 U602 ( .A(n478), .ZN(n696) );
  NAND2_X1 U603 ( .A1(n358), .A2(n371), .ZN(n478) );
  INV_X1 U604 ( .A(KEYINPUT48), .ZN(n594) );
  INV_X1 U605 ( .A(KEYINPUT87), .ZN(n606) );
  XNOR2_X1 U606 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U607 ( .A(n658), .B(n657), .ZN(G69) );
  XNOR2_X1 U608 ( .A(G119), .B(KEYINPUT3), .ZN(n481) );
  XOR2_X2 U609 ( .A(KEYINPUT4), .B(KEYINPUT69), .Z(n756) );
  NAND2_X1 U610 ( .A1(G224), .A2(n767), .ZN(n486) );
  XNOR2_X1 U611 ( .A(KEYINPUT17), .B(KEYINPUT81), .ZN(n487) );
  NAND2_X1 U612 ( .A1(G210), .A2(n492), .ZN(n489) );
  INV_X1 U613 ( .A(KEYINPUT93), .ZN(n488) );
  NAND2_X1 U614 ( .A1(n492), .A2(G214), .ZN(n493) );
  INV_X1 U615 ( .A(n566), .ZN(n717) );
  NAND2_X1 U616 ( .A1(G227), .A2(n767), .ZN(n495) );
  INV_X1 U617 ( .A(n706), .ZN(n617) );
  XNOR2_X1 U618 ( .A(n496), .B(KEYINPUT106), .ZN(n500) );
  XNOR2_X1 U619 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U620 ( .A(n500), .B(n499), .Z(n504) );
  NAND2_X1 U621 ( .A1(G234), .A2(n767), .ZN(n501) );
  XNOR2_X1 U622 ( .A(n502), .B(n501), .ZN(n531) );
  NAND2_X1 U623 ( .A1(G217), .A2(n531), .ZN(n503) );
  XNOR2_X1 U624 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U625 ( .A(n506), .B(n505), .ZN(n748) );
  NOR2_X1 U626 ( .A1(n748), .A2(G902), .ZN(n507) );
  XNOR2_X1 U627 ( .A(n507), .B(G478), .ZN(n588) );
  XNOR2_X1 U628 ( .A(KEYINPUT13), .B(KEYINPUT104), .ZN(n516) );
  XNOR2_X1 U629 ( .A(n511), .B(n532), .ZN(n755) );
  NAND2_X1 U630 ( .A1(G214), .A2(n524), .ZN(n514) );
  NAND2_X1 U631 ( .A1(n588), .A2(n573), .ZN(n517) );
  XNOR2_X1 U632 ( .A(KEYINPUT107), .B(n517), .ZN(n554) );
  XNOR2_X1 U633 ( .A(G472), .B(KEYINPUT74), .ZN(n527) );
  XNOR2_X1 U634 ( .A(n521), .B(n520), .ZN(n522) );
  AND2_X1 U635 ( .A1(n524), .A2(G210), .ZN(n525) );
  INV_X1 U636 ( .A(n558), .ZN(n623) );
  XNOR2_X1 U637 ( .A(KEYINPUT6), .B(n357), .ZN(n613) );
  NAND2_X1 U638 ( .A1(n554), .A2(n613), .ZN(n544) );
  XOR2_X1 U639 ( .A(KEYINPUT14), .B(n528), .Z(n733) );
  NAND2_X1 U640 ( .A1(n631), .A2(G234), .ZN(n529) );
  NAND2_X1 U641 ( .A1(G221), .A2(n535), .ZN(n530) );
  XOR2_X1 U642 ( .A(KEYINPUT21), .B(n530), .Z(n607) );
  INV_X1 U643 ( .A(n607), .ZN(n702) );
  NAND2_X1 U644 ( .A1(n531), .A2(G221), .ZN(n534) );
  NAND2_X1 U645 ( .A1(G217), .A2(n535), .ZN(n536) );
  XNOR2_X1 U646 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U647 ( .A(KEYINPUT98), .B(n538), .ZN(n539) );
  INV_X2 U648 ( .A(G953), .ZN(n701) );
  NAND2_X1 U649 ( .A1(G952), .A2(n701), .ZN(n596) );
  NOR2_X1 U650 ( .A1(n767), .A2(G900), .ZN(n540) );
  NAND2_X1 U651 ( .A1(G902), .A2(n540), .ZN(n541) );
  NAND2_X1 U652 ( .A1(n596), .A2(n541), .ZN(n570) );
  NAND2_X1 U653 ( .A1(n703), .A2(n570), .ZN(n542) );
  NOR2_X1 U654 ( .A1(n702), .A2(n542), .ZN(n543) );
  NAND2_X1 U655 ( .A1(n461), .A2(n543), .ZN(n559) );
  NOR2_X1 U656 ( .A1(n544), .A2(n559), .ZN(n550) );
  NAND2_X1 U657 ( .A1(n617), .A2(n550), .ZN(n545) );
  NOR2_X1 U658 ( .A1(n717), .A2(n545), .ZN(n546) );
  XNOR2_X1 U659 ( .A(n546), .B(KEYINPUT43), .ZN(n547) );
  NOR2_X1 U660 ( .A1(n582), .A2(n547), .ZN(n694) );
  INV_X1 U661 ( .A(n550), .ZN(n551) );
  XOR2_X1 U662 ( .A(KEYINPUT36), .B(n552), .Z(n553) );
  NOR2_X1 U663 ( .A1(n617), .A2(n553), .ZN(n691) );
  BUF_X1 U664 ( .A(n554), .Z(n685) );
  NOR2_X1 U665 ( .A1(n588), .A2(n573), .ZN(n688) );
  NOR2_X1 U666 ( .A1(n624), .A2(KEYINPUT84), .ZN(n555) );
  NAND2_X1 U667 ( .A1(KEYINPUT84), .A2(n624), .ZN(n564) );
  INV_X1 U668 ( .A(KEYINPUT19), .ZN(n556) );
  INV_X1 U669 ( .A(KEYINPUT110), .ZN(n557) );
  INV_X1 U670 ( .A(n609), .ZN(n560) );
  XNOR2_X1 U671 ( .A(n433), .B(KEYINPUT112), .ZN(n562) );
  NAND2_X1 U672 ( .A1(n563), .A2(n562), .ZN(n587) );
  NAND2_X1 U673 ( .A1(n564), .A2(n682), .ZN(n565) );
  NAND2_X1 U674 ( .A1(n565), .A2(KEYINPUT47), .ZN(n576) );
  NAND2_X1 U675 ( .A1(n609), .A2(n566), .ZN(n568) );
  INV_X1 U676 ( .A(n605), .ZN(n574) );
  NOR2_X1 U677 ( .A1(n583), .A2(n574), .ZN(n575) );
  NAND2_X1 U678 ( .A1(n582), .A2(n575), .ZN(n681) );
  NAND2_X1 U679 ( .A1(n576), .A2(n681), .ZN(n579) );
  NOR2_X1 U680 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U681 ( .A(n582), .B(KEYINPUT38), .ZN(n716) );
  XNOR2_X1 U682 ( .A(KEYINPUT73), .B(KEYINPUT39), .ZN(n584) );
  XNOR2_X1 U683 ( .A(KEYINPUT40), .B(KEYINPUT114), .ZN(n586) );
  INV_X1 U684 ( .A(n587), .ZN(n591) );
  NOR2_X1 U685 ( .A1(n717), .A2(n716), .ZN(n722) );
  NAND2_X1 U686 ( .A1(n589), .A2(n588), .ZN(n608) );
  INV_X1 U687 ( .A(n608), .ZN(n719) );
  NAND2_X1 U688 ( .A1(n722), .A2(n719), .ZN(n590) );
  XNOR2_X1 U689 ( .A(n590), .B(KEYINPUT41), .ZN(n714) );
  NAND2_X1 U690 ( .A1(n591), .A2(n714), .ZN(n592) );
  XNOR2_X1 U691 ( .A(n592), .B(KEYINPUT42), .ZN(n773) );
  NAND2_X1 U692 ( .A1(n688), .A2(n595), .ZN(n693) );
  NOR2_X1 U693 ( .A1(G898), .A2(n701), .ZN(n654) );
  NAND2_X1 U694 ( .A1(n654), .A2(G902), .ZN(n597) );
  NAND2_X1 U695 ( .A1(n597), .A2(n596), .ZN(n598) );
  INV_X1 U696 ( .A(n619), .ZN(n600) );
  NAND2_X1 U697 ( .A1(n613), .A2(n600), .ZN(n601) );
  XNOR2_X1 U698 ( .A(n601), .B(KEYINPUT33), .ZN(n726) );
  NAND2_X1 U699 ( .A1(n602), .A2(n726), .ZN(n604) );
  XOR2_X1 U700 ( .A(KEYINPUT34), .B(KEYINPUT82), .Z(n603) );
  NOR2_X1 U701 ( .A1(n609), .A2(n706), .ZN(n610) );
  NAND2_X1 U702 ( .A1(n427), .A2(n610), .ZN(n611) );
  NOR2_X1 U703 ( .A1(n389), .A2(n611), .ZN(n677) );
  NAND2_X1 U704 ( .A1(n427), .A2(n706), .ZN(n612) );
  XNOR2_X1 U705 ( .A(KEYINPUT109), .B(n612), .ZN(n614) );
  NAND2_X1 U706 ( .A1(n616), .A2(n775), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n629), .A2(KEYINPUT44), .ZN(n627) );
  XOR2_X1 U708 ( .A(KEYINPUT31), .B(KEYINPUT101), .Z(n620) );
  NOR2_X1 U709 ( .A1(n357), .A2(n619), .ZN(n712) );
  NOR2_X1 U710 ( .A1(n671), .A2(n625), .ZN(n626) );
  XNOR2_X1 U711 ( .A(n631), .B(KEYINPUT85), .ZN(n632) );
  AND2_X1 U712 ( .A1(n632), .A2(KEYINPUT2), .ZN(n633) );
  NAND2_X1 U713 ( .A1(n695), .A2(n633), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n697), .A2(n635), .ZN(n636) );
  NAND2_X1 U715 ( .A1(n746), .A2(G475), .ZN(n640) );
  XNOR2_X1 U716 ( .A(n638), .B(KEYINPUT59), .ZN(n639) );
  XNOR2_X1 U717 ( .A(n640), .B(n639), .ZN(n642) );
  NOR2_X1 U718 ( .A1(n767), .A2(G952), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n642), .A2(n739), .ZN(n644) );
  XNOR2_X1 U720 ( .A(KEYINPUT60), .B(KEYINPUT65), .ZN(n643) );
  XNOR2_X1 U721 ( .A(n644), .B(n643), .ZN(G60) );
  NAND2_X1 U722 ( .A1(n701), .A2(n359), .ZN(n648) );
  NAND2_X1 U723 ( .A1(G953), .A2(G224), .ZN(n645) );
  XNOR2_X1 U724 ( .A(KEYINPUT61), .B(n645), .ZN(n646) );
  NAND2_X1 U725 ( .A1(n646), .A2(G898), .ZN(n647) );
  NAND2_X1 U726 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U727 ( .A(n649), .B(KEYINPUT123), .ZN(n658) );
  XOR2_X1 U728 ( .A(n650), .B(G101), .Z(n651) );
  XNOR2_X1 U729 ( .A(n652), .B(n651), .ZN(n653) );
  NOR2_X1 U730 ( .A1(n654), .A2(n653), .ZN(n656) );
  INV_X1 U731 ( .A(KEYINPUT122), .ZN(n655) );
  XOR2_X1 U732 ( .A(KEYINPUT54), .B(KEYINPUT120), .Z(n660) );
  XNOR2_X1 U733 ( .A(KEYINPUT83), .B(KEYINPUT55), .ZN(n659) );
  XNOR2_X1 U734 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U735 ( .A(n360), .B(n661), .ZN(n664) );
  INV_X1 U736 ( .A(KEYINPUT56), .ZN(n665) );
  XNOR2_X1 U737 ( .A(n666), .B(n665), .ZN(G51) );
  XOR2_X1 U738 ( .A(n667), .B(KEYINPUT62), .Z(n669) );
  NAND2_X1 U739 ( .A1(n746), .A2(G472), .ZN(n668) );
  XNOR2_X1 U740 ( .A(n670), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U741 ( .A(G101), .B(n671), .Z(G3) );
  NAND2_X1 U742 ( .A1(n673), .A2(n685), .ZN(n672) );
  XNOR2_X1 U743 ( .A(n672), .B(G104), .ZN(G6) );
  XOR2_X1 U744 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n675) );
  NAND2_X1 U745 ( .A1(n673), .A2(n688), .ZN(n674) );
  XNOR2_X1 U746 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U747 ( .A(G107), .B(n676), .ZN(G9) );
  XOR2_X1 U748 ( .A(G110), .B(n677), .Z(G12) );
  XOR2_X1 U749 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n679) );
  NAND2_X1 U750 ( .A1(n682), .A2(n688), .ZN(n678) );
  XNOR2_X1 U751 ( .A(n679), .B(n678), .ZN(n680) );
  XOR2_X1 U752 ( .A(G128), .B(n680), .Z(G30) );
  XNOR2_X1 U753 ( .A(G143), .B(n681), .ZN(G45) );
  NAND2_X1 U754 ( .A1(n682), .A2(n685), .ZN(n683) );
  XNOR2_X1 U755 ( .A(n683), .B(KEYINPUT116), .ZN(n684) );
  XNOR2_X1 U756 ( .A(G146), .B(n684), .ZN(G48) );
  XOR2_X1 U757 ( .A(G113), .B(KEYINPUT117), .Z(n687) );
  NAND2_X1 U758 ( .A1(n689), .A2(n685), .ZN(n686) );
  XNOR2_X1 U759 ( .A(n687), .B(n686), .ZN(G15) );
  NAND2_X1 U760 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U761 ( .A(n690), .B(G116), .ZN(G18) );
  XNOR2_X1 U762 ( .A(n691), .B(G125), .ZN(n692) );
  XNOR2_X1 U763 ( .A(n692), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U764 ( .A(G134), .B(n693), .ZN(G36) );
  XOR2_X1 U765 ( .A(G140), .B(n694), .Z(G42) );
  AND2_X1 U766 ( .A1(n695), .A2(KEYINPUT2), .ZN(n699) );
  AND2_X1 U767 ( .A1(n359), .A2(n696), .ZN(n698) );
  NOR2_X1 U768 ( .A1(n699), .A2(n698), .ZN(n737) );
  NAND2_X1 U769 ( .A1(n726), .A2(n714), .ZN(n700) );
  NAND2_X1 U770 ( .A1(n701), .A2(n700), .ZN(n735) );
  NAND2_X1 U771 ( .A1(n427), .A2(n702), .ZN(n704) );
  XNOR2_X1 U772 ( .A(n704), .B(KEYINPUT49), .ZN(n710) );
  NOR2_X1 U773 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U774 ( .A(KEYINPUT50), .B(n707), .Z(n708) );
  NAND2_X1 U775 ( .A1(n357), .A2(n708), .ZN(n709) );
  NOR2_X1 U776 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U777 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U778 ( .A(KEYINPUT51), .B(n713), .ZN(n715) );
  NAND2_X1 U779 ( .A1(n715), .A2(n714), .ZN(n729) );
  NAND2_X1 U780 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U781 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U782 ( .A(n720), .B(KEYINPUT118), .ZN(n724) );
  NAND2_X1 U783 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U784 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U785 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U786 ( .A(KEYINPUT119), .B(n727), .Z(n728) );
  NAND2_X1 U787 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U788 ( .A(KEYINPUT52), .B(n730), .ZN(n731) );
  NAND2_X1 U789 ( .A1(n731), .A2(G952), .ZN(n732) );
  NOR2_X1 U790 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U791 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U792 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U793 ( .A(KEYINPUT53), .B(n738), .Z(G75) );
  INV_X1 U794 ( .A(n739), .ZN(n754) );
  XOR2_X1 U795 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n742) );
  XNOR2_X1 U796 ( .A(n740), .B(KEYINPUT121), .ZN(n741) );
  XNOR2_X1 U797 ( .A(n742), .B(n741), .ZN(n744) );
  NAND2_X1 U798 ( .A1(n746), .A2(G469), .ZN(n743) );
  XOR2_X1 U799 ( .A(n744), .B(n743), .Z(n745) );
  NOR2_X1 U800 ( .A1(n754), .A2(n745), .ZN(G54) );
  NAND2_X1 U801 ( .A1(G478), .A2(n750), .ZN(n747) );
  XNOR2_X1 U802 ( .A(n748), .B(n747), .ZN(n749) );
  NOR2_X1 U803 ( .A1(n754), .A2(n749), .ZN(G63) );
  NAND2_X1 U804 ( .A1(G217), .A2(n750), .ZN(n751) );
  XNOR2_X1 U805 ( .A(n752), .B(n751), .ZN(n753) );
  NOR2_X1 U806 ( .A1(n754), .A2(n753), .ZN(G66) );
  XNOR2_X1 U807 ( .A(n756), .B(n755), .ZN(n758) );
  XNOR2_X1 U808 ( .A(n757), .B(n758), .ZN(n764) );
  INV_X1 U809 ( .A(n764), .ZN(n759) );
  XNOR2_X1 U810 ( .A(G227), .B(n759), .ZN(n760) );
  NAND2_X1 U811 ( .A1(n760), .A2(G900), .ZN(n761) );
  XOR2_X1 U812 ( .A(KEYINPUT125), .B(n761), .Z(n762) );
  NAND2_X1 U813 ( .A1(G953), .A2(n762), .ZN(n769) );
  XNOR2_X1 U814 ( .A(KEYINPUT124), .B(n764), .ZN(n765) );
  XNOR2_X1 U815 ( .A(n358), .B(n765), .ZN(n766) );
  NAND2_X1 U816 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U817 ( .A1(n769), .A2(n768), .ZN(G72) );
  XOR2_X1 U818 ( .A(G131), .B(KEYINPUT127), .Z(n770) );
  XNOR2_X1 U819 ( .A(n387), .B(n770), .ZN(G33) );
  XOR2_X1 U820 ( .A(n390), .B(G122), .Z(G24) );
  XNOR2_X1 U821 ( .A(G137), .B(n773), .ZN(n774) );
  XNOR2_X1 U822 ( .A(n774), .B(KEYINPUT126), .ZN(G39) );
  XNOR2_X1 U823 ( .A(G119), .B(n775), .ZN(G21) );
endmodule

