

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588;

  XNOR2_X1 U324 ( .A(n431), .B(n325), .ZN(n326) );
  XNOR2_X1 U325 ( .A(n327), .B(n326), .ZN(n364) );
  XNOR2_X1 U326 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U327 ( .A(n450), .B(n449), .ZN(G1349GAT) );
  XOR2_X1 U328 ( .A(G43GAT), .B(G29GAT), .Z(n293) );
  XNOR2_X1 U329 ( .A(KEYINPUT7), .B(G50GAT), .ZN(n292) );
  XNOR2_X1 U330 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U331 ( .A(n294), .B(KEYINPUT69), .Z(n296) );
  XNOR2_X1 U332 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n295) );
  XNOR2_X1 U333 ( .A(n296), .B(n295), .ZN(n340) );
  XNOR2_X1 U334 ( .A(G99GAT), .B(G85GAT), .ZN(n325) );
  XNOR2_X1 U335 ( .A(n325), .B(G92GAT), .ZN(n298) );
  NAND2_X1 U336 ( .A1(G232GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U337 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U338 ( .A(KEYINPUT65), .B(G106GAT), .Z(n300) );
  XNOR2_X1 U339 ( .A(G190GAT), .B(G162GAT), .ZN(n299) );
  XNOR2_X1 U340 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U341 ( .A(n302), .B(n301), .Z(n307) );
  XOR2_X1 U342 ( .A(G134GAT), .B(KEYINPUT75), .Z(n404) );
  XOR2_X1 U343 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n304) );
  XNOR2_X1 U344 ( .A(G218GAT), .B(KEYINPUT9), .ZN(n303) );
  XNOR2_X1 U345 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U346 ( .A(n404), .B(n305), .ZN(n306) );
  XNOR2_X1 U347 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U348 ( .A(n340), .B(n308), .Z(n565) );
  XNOR2_X1 U349 ( .A(G176GAT), .B(G92GAT), .ZN(n309) );
  XNOR2_X1 U350 ( .A(n309), .B(G64GAT), .ZN(n374) );
  INV_X1 U351 ( .A(KEYINPUT32), .ZN(n310) );
  NAND2_X1 U352 ( .A1(n374), .A2(n310), .ZN(n313) );
  INV_X1 U353 ( .A(n374), .ZN(n311) );
  NAND2_X1 U354 ( .A1(n311), .A2(KEYINPUT32), .ZN(n312) );
  NAND2_X1 U355 ( .A1(n313), .A2(n312), .ZN(n315) );
  NAND2_X1 U356 ( .A1(G230GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U357 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U358 ( .A(KEYINPUT74), .B(KEYINPUT73), .Z(n317) );
  XNOR2_X1 U359 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n316) );
  XNOR2_X1 U360 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U361 ( .A(n319), .B(n318), .Z(n324) );
  XNOR2_X1 U362 ( .A(G57GAT), .B(KEYINPUT72), .ZN(n320) );
  XNOR2_X1 U363 ( .A(n320), .B(KEYINPUT13), .ZN(n355) );
  XOR2_X1 U364 ( .A(G78GAT), .B(G106GAT), .Z(n322) );
  XNOR2_X1 U365 ( .A(G148GAT), .B(G204GAT), .ZN(n321) );
  XNOR2_X1 U366 ( .A(n322), .B(n321), .ZN(n417) );
  XNOR2_X1 U367 ( .A(n355), .B(n417), .ZN(n323) );
  XNOR2_X1 U368 ( .A(n324), .B(n323), .ZN(n327) );
  XOR2_X1 U369 ( .A(G120GAT), .B(G71GAT), .Z(n431) );
  XNOR2_X1 U370 ( .A(KEYINPUT41), .B(n364), .ZN(n446) );
  XOR2_X1 U371 ( .A(G1GAT), .B(G15GAT), .Z(n351) );
  XOR2_X1 U372 ( .A(G141GAT), .B(G22GAT), .Z(n416) );
  XOR2_X1 U373 ( .A(n351), .B(n416), .Z(n329) );
  NAND2_X1 U374 ( .A1(G229GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U375 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U376 ( .A(G169GAT), .B(G8GAT), .Z(n381) );
  XOR2_X1 U377 ( .A(n330), .B(n381), .Z(n338) );
  XOR2_X1 U378 ( .A(KEYINPUT70), .B(KEYINPUT66), .Z(n332) );
  XNOR2_X1 U379 ( .A(G113GAT), .B(G197GAT), .ZN(n331) );
  XNOR2_X1 U380 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U381 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n334) );
  XNOR2_X1 U382 ( .A(KEYINPUT68), .B(KEYINPUT30), .ZN(n333) );
  XNOR2_X1 U383 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U384 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U385 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U386 ( .A(n340), .B(n339), .Z(n571) );
  NOR2_X1 U387 ( .A1(n446), .A2(n571), .ZN(n341) );
  XNOR2_X1 U388 ( .A(n341), .B(KEYINPUT46), .ZN(n360) );
  XOR2_X1 U389 ( .A(G78GAT), .B(G64GAT), .Z(n343) );
  XNOR2_X1 U390 ( .A(G8GAT), .B(G71GAT), .ZN(n342) );
  XNOR2_X1 U391 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U392 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n345) );
  XNOR2_X1 U393 ( .A(G22GAT), .B(KEYINPUT76), .ZN(n344) );
  XNOR2_X1 U394 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U395 ( .A(n347), .B(n346), .ZN(n359) );
  XOR2_X1 U396 ( .A(G211GAT), .B(G155GAT), .Z(n349) );
  XNOR2_X1 U397 ( .A(G183GAT), .B(G127GAT), .ZN(n348) );
  XNOR2_X1 U398 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U399 ( .A(n351), .B(n350), .Z(n353) );
  NAND2_X1 U400 ( .A1(G231GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U401 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U402 ( .A(n354), .B(KEYINPUT15), .Z(n357) );
  XNOR2_X1 U403 ( .A(n355), .B(KEYINPUT77), .ZN(n356) );
  XNOR2_X1 U404 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U405 ( .A(n359), .B(n358), .ZN(n580) );
  NOR2_X1 U406 ( .A1(n360), .A2(n580), .ZN(n361) );
  XNOR2_X1 U407 ( .A(n361), .B(KEYINPUT107), .ZN(n362) );
  NOR2_X1 U408 ( .A1(n565), .A2(n362), .ZN(n363) );
  XNOR2_X1 U409 ( .A(n363), .B(KEYINPUT47), .ZN(n369) );
  INV_X1 U410 ( .A(n565), .ZN(n558) );
  XNOR2_X1 U411 ( .A(KEYINPUT36), .B(n558), .ZN(n585) );
  INV_X1 U412 ( .A(n580), .ZN(n555) );
  NOR2_X1 U413 ( .A1(n585), .A2(n555), .ZN(n365) );
  XOR2_X1 U414 ( .A(KEYINPUT45), .B(n365), .Z(n366) );
  NOR2_X1 U415 ( .A1(n364), .A2(n366), .ZN(n367) );
  XOR2_X1 U416 ( .A(n571), .B(KEYINPUT71), .Z(n533) );
  NAND2_X1 U417 ( .A1(n367), .A2(n533), .ZN(n368) );
  NAND2_X1 U418 ( .A1(n369), .A2(n368), .ZN(n370) );
  XNOR2_X1 U419 ( .A(n370), .B(KEYINPUT48), .ZN(n525) );
  XOR2_X1 U420 ( .A(KEYINPUT18), .B(G190GAT), .Z(n372) );
  XNOR2_X1 U421 ( .A(KEYINPUT19), .B(G183GAT), .ZN(n371) );
  XNOR2_X1 U422 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U423 ( .A(KEYINPUT17), .B(n373), .Z(n441) );
  BUF_X1 U424 ( .A(n374), .Z(n375) );
  XNOR2_X1 U425 ( .A(n441), .B(n375), .ZN(n385) );
  XOR2_X1 U426 ( .A(G211GAT), .B(KEYINPUT21), .Z(n377) );
  XNOR2_X1 U427 ( .A(G197GAT), .B(G218GAT), .ZN(n376) );
  XNOR2_X1 U428 ( .A(n377), .B(n376), .ZN(n421) );
  XOR2_X1 U429 ( .A(n421), .B(G204GAT), .Z(n379) );
  NAND2_X1 U430 ( .A1(G226GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U431 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U432 ( .A(n380), .B(KEYINPUT88), .Z(n383) );
  XNOR2_X1 U433 ( .A(G36GAT), .B(n381), .ZN(n382) );
  XNOR2_X1 U434 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U435 ( .A(n385), .B(n384), .ZN(n490) );
  NAND2_X1 U436 ( .A1(n525), .A2(n490), .ZN(n387) );
  XOR2_X1 U437 ( .A(KEYINPUT118), .B(KEYINPUT54), .Z(n386) );
  XNOR2_X1 U438 ( .A(n387), .B(n386), .ZN(n412) );
  XOR2_X1 U439 ( .A(KEYINPUT83), .B(G162GAT), .Z(n389) );
  XNOR2_X1 U440 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n388) );
  XNOR2_X1 U441 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U442 ( .A(KEYINPUT3), .B(n390), .ZN(n426) );
  XOR2_X1 U443 ( .A(KEYINPUT84), .B(KEYINPUT4), .Z(n392) );
  XNOR2_X1 U444 ( .A(KEYINPUT1), .B(KEYINPUT85), .ZN(n391) );
  XNOR2_X1 U445 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U446 ( .A(G148GAT), .B(KEYINPUT86), .Z(n394) );
  XNOR2_X1 U447 ( .A(G141GAT), .B(KEYINPUT5), .ZN(n393) );
  XNOR2_X1 U448 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U449 ( .A(n396), .B(n395), .Z(n410) );
  XOR2_X1 U450 ( .A(G127GAT), .B(KEYINPUT79), .Z(n398) );
  XNOR2_X1 U451 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n397) );
  XNOR2_X1 U452 ( .A(n398), .B(n397), .ZN(n430) );
  XOR2_X1 U453 ( .A(n430), .B(G1GAT), .Z(n400) );
  NAND2_X1 U454 ( .A1(G225GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U455 ( .A(n400), .B(n399), .ZN(n408) );
  XOR2_X1 U456 ( .A(KEYINPUT87), .B(KEYINPUT6), .Z(n402) );
  XNOR2_X1 U457 ( .A(G120GAT), .B(G57GAT), .ZN(n401) );
  XNOR2_X1 U458 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U459 ( .A(n403), .B(G85GAT), .Z(n406) );
  XNOR2_X1 U460 ( .A(G29GAT), .B(n404), .ZN(n405) );
  XNOR2_X1 U461 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U462 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U463 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U464 ( .A(n426), .B(n411), .ZN(n470) );
  INV_X1 U465 ( .A(n470), .ZN(n513) );
  NAND2_X1 U466 ( .A1(n412), .A2(n513), .ZN(n413) );
  XOR2_X1 U467 ( .A(KEYINPUT64), .B(n413), .Z(n570) );
  XOR2_X1 U468 ( .A(KEYINPUT81), .B(KEYINPUT22), .Z(n415) );
  XNOR2_X1 U469 ( .A(G50GAT), .B(KEYINPUT23), .ZN(n414) );
  XNOR2_X1 U470 ( .A(n415), .B(n414), .ZN(n425) );
  XOR2_X1 U471 ( .A(n417), .B(n416), .Z(n419) );
  NAND2_X1 U472 ( .A1(G228GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U473 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U474 ( .A(n420), .B(KEYINPUT24), .Z(n423) );
  XNOR2_X1 U475 ( .A(n421), .B(KEYINPUT82), .ZN(n422) );
  XNOR2_X1 U476 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U477 ( .A(n425), .B(n424), .ZN(n427) );
  XNOR2_X1 U478 ( .A(n427), .B(n426), .ZN(n458) );
  NAND2_X1 U479 ( .A1(n570), .A2(n458), .ZN(n429) );
  XOR2_X1 U480 ( .A(KEYINPUT119), .B(KEYINPUT55), .Z(n428) );
  XNOR2_X1 U481 ( .A(n429), .B(n428), .ZN(n444) );
  XOR2_X1 U482 ( .A(n431), .B(n430), .Z(n433) );
  NAND2_X1 U483 ( .A1(G227GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U484 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U485 ( .A(KEYINPUT80), .B(KEYINPUT20), .Z(n435) );
  XNOR2_X1 U486 ( .A(G15GAT), .B(G176GAT), .ZN(n434) );
  XNOR2_X1 U487 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U488 ( .A(n437), .B(n436), .Z(n443) );
  XOR2_X1 U489 ( .A(G99GAT), .B(G134GAT), .Z(n439) );
  XNOR2_X1 U490 ( .A(G169GAT), .B(G43GAT), .ZN(n438) );
  XNOR2_X1 U491 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U492 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U493 ( .A(n443), .B(n442), .ZN(n528) );
  AND2_X1 U494 ( .A1(n444), .A2(n528), .ZN(n445) );
  XNOR2_X2 U495 ( .A(KEYINPUT120), .B(n445), .ZN(n566) );
  BUF_X1 U496 ( .A(n446), .Z(n552) );
  INV_X1 U497 ( .A(n552), .ZN(n536) );
  NAND2_X1 U498 ( .A1(n566), .A2(n536), .ZN(n450) );
  XOR2_X1 U499 ( .A(G176GAT), .B(KEYINPUT56), .Z(n448) );
  XNOR2_X1 U500 ( .A(KEYINPUT57), .B(KEYINPUT122), .ZN(n447) );
  XNOR2_X1 U501 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n472) );
  NOR2_X1 U502 ( .A1(n533), .A2(n364), .ZN(n485) );
  XOR2_X1 U503 ( .A(KEYINPUT78), .B(KEYINPUT16), .Z(n452) );
  NAND2_X1 U504 ( .A1(n580), .A2(n558), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n452), .B(n451), .ZN(n468) );
  XOR2_X1 U506 ( .A(n490), .B(KEYINPUT27), .Z(n461) );
  NOR2_X1 U507 ( .A1(n461), .A2(n513), .ZN(n453) );
  XOR2_X1 U508 ( .A(KEYINPUT89), .B(n453), .Z(n526) );
  XOR2_X1 U509 ( .A(KEYINPUT28), .B(n458), .Z(n531) );
  NOR2_X1 U510 ( .A1(n528), .A2(n531), .ZN(n454) );
  NAND2_X1 U511 ( .A1(n526), .A2(n454), .ZN(n455) );
  XOR2_X1 U512 ( .A(KEYINPUT90), .B(n455), .Z(n466) );
  NAND2_X1 U513 ( .A1(n528), .A2(n490), .ZN(n456) );
  NAND2_X1 U514 ( .A1(n458), .A2(n456), .ZN(n457) );
  XNOR2_X1 U515 ( .A(n457), .B(KEYINPUT25), .ZN(n463) );
  NOR2_X1 U516 ( .A1(n458), .A2(n528), .ZN(n459) );
  XNOR2_X1 U517 ( .A(n459), .B(KEYINPUT26), .ZN(n569) );
  INV_X1 U518 ( .A(n569), .ZN(n460) );
  NOR2_X1 U519 ( .A1(n461), .A2(n460), .ZN(n462) );
  NOR2_X1 U520 ( .A1(n463), .A2(n462), .ZN(n464) );
  NOR2_X1 U521 ( .A1(n470), .A2(n464), .ZN(n465) );
  NOR2_X1 U522 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U523 ( .A(KEYINPUT91), .B(n467), .ZN(n481) );
  AND2_X1 U524 ( .A1(n468), .A2(n481), .ZN(n500) );
  NAND2_X1 U525 ( .A1(n485), .A2(n500), .ZN(n469) );
  XOR2_X1 U526 ( .A(KEYINPUT92), .B(n469), .Z(n478) );
  NAND2_X1 U527 ( .A1(n470), .A2(n478), .ZN(n471) );
  XNOR2_X1 U528 ( .A(n472), .B(n471), .ZN(G1324GAT) );
  XOR2_X1 U529 ( .A(G8GAT), .B(KEYINPUT93), .Z(n474) );
  NAND2_X1 U530 ( .A1(n490), .A2(n478), .ZN(n473) );
  XNOR2_X1 U531 ( .A(n474), .B(n473), .ZN(G1325GAT) );
  XOR2_X1 U532 ( .A(KEYINPUT94), .B(KEYINPUT35), .Z(n476) );
  NAND2_X1 U533 ( .A1(n528), .A2(n478), .ZN(n475) );
  XNOR2_X1 U534 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U535 ( .A(G15GAT), .B(n477), .ZN(G1326GAT) );
  NAND2_X1 U536 ( .A1(n478), .A2(n531), .ZN(n479) );
  XNOR2_X1 U537 ( .A(n479), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U538 ( .A(KEYINPUT38), .B(KEYINPUT97), .Z(n487) );
  NOR2_X1 U539 ( .A1(n585), .A2(n580), .ZN(n480) );
  NAND2_X1 U540 ( .A1(n481), .A2(n480), .ZN(n482) );
  XNOR2_X1 U541 ( .A(KEYINPUT96), .B(n482), .ZN(n484) );
  XOR2_X1 U542 ( .A(KEYINPUT37), .B(KEYINPUT95), .Z(n483) );
  XNOR2_X1 U543 ( .A(n484), .B(n483), .ZN(n511) );
  NAND2_X1 U544 ( .A1(n485), .A2(n511), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n487), .B(n486), .ZN(n498) );
  NOR2_X1 U546 ( .A1(n498), .A2(n513), .ZN(n489) );
  XNOR2_X1 U547 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n489), .B(n488), .ZN(G1328GAT) );
  INV_X1 U549 ( .A(n490), .ZN(n515) );
  NOR2_X1 U550 ( .A1(n498), .A2(n515), .ZN(n492) );
  XNOR2_X1 U551 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U553 ( .A(G36GAT), .B(n493), .ZN(G1329GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT101), .B(KEYINPUT40), .Z(n495) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(KEYINPUT100), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(n497) );
  INV_X1 U557 ( .A(n528), .ZN(n517) );
  NOR2_X1 U558 ( .A1(n498), .A2(n517), .ZN(n496) );
  XOR2_X1 U559 ( .A(n497), .B(n496), .Z(G1330GAT) );
  INV_X1 U560 ( .A(n531), .ZN(n521) );
  NOR2_X1 U561 ( .A1(n521), .A2(n498), .ZN(n499) );
  XOR2_X1 U562 ( .A(G50GAT), .B(n499), .Z(G1331GAT) );
  AND2_X1 U563 ( .A1(n536), .A2(n571), .ZN(n512) );
  NAND2_X1 U564 ( .A1(n500), .A2(n512), .ZN(n507) );
  NOR2_X1 U565 ( .A1(n513), .A2(n507), .ZN(n502) );
  XNOR2_X1 U566 ( .A(KEYINPUT102), .B(KEYINPUT42), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U568 ( .A(G57GAT), .B(n503), .Z(G1332GAT) );
  NOR2_X1 U569 ( .A1(n515), .A2(n507), .ZN(n505) );
  XNOR2_X1 U570 ( .A(G64GAT), .B(KEYINPUT103), .ZN(n504) );
  XNOR2_X1 U571 ( .A(n505), .B(n504), .ZN(G1333GAT) );
  NOR2_X1 U572 ( .A1(n517), .A2(n507), .ZN(n506) );
  XOR2_X1 U573 ( .A(G71GAT), .B(n506), .Z(G1334GAT) );
  NOR2_X1 U574 ( .A1(n521), .A2(n507), .ZN(n509) );
  XNOR2_X1 U575 ( .A(KEYINPUT43), .B(KEYINPUT104), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U577 ( .A(G78GAT), .B(n510), .ZN(G1335GAT) );
  NAND2_X1 U578 ( .A1(n512), .A2(n511), .ZN(n520) );
  NOR2_X1 U579 ( .A1(n513), .A2(n520), .ZN(n514) );
  XOR2_X1 U580 ( .A(G85GAT), .B(n514), .Z(G1336GAT) );
  NOR2_X1 U581 ( .A1(n515), .A2(n520), .ZN(n516) );
  XOR2_X1 U582 ( .A(G92GAT), .B(n516), .Z(G1337GAT) );
  NOR2_X1 U583 ( .A1(n517), .A2(n520), .ZN(n519) );
  XNOR2_X1 U584 ( .A(G99GAT), .B(KEYINPUT105), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(G1338GAT) );
  NOR2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n523) );
  XNOR2_X1 U587 ( .A(KEYINPUT44), .B(KEYINPUT106), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U589 ( .A(G106GAT), .B(n524), .Z(G1339GAT) );
  XOR2_X1 U590 ( .A(G113GAT), .B(KEYINPUT111), .Z(n535) );
  NAND2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U592 ( .A(KEYINPUT108), .B(n527), .Z(n547) );
  NAND2_X1 U593 ( .A1(n528), .A2(n547), .ZN(n529) );
  XOR2_X1 U594 ( .A(KEYINPUT109), .B(n529), .Z(n530) );
  NOR2_X1 U595 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U596 ( .A(KEYINPUT110), .B(n532), .ZN(n543) );
  INV_X1 U597 ( .A(n533), .ZN(n561) );
  NAND2_X1 U598 ( .A1(n543), .A2(n561), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT49), .B(KEYINPUT112), .Z(n538) );
  NAND2_X1 U601 ( .A1(n543), .A2(n536), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U603 ( .A(G120GAT), .B(n539), .ZN(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT113), .B(KEYINPUT50), .Z(n541) );
  NAND2_X1 U605 ( .A1(n580), .A2(n543), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT51), .B(KEYINPUT114), .Z(n545) );
  NAND2_X1 U609 ( .A1(n565), .A2(n543), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U611 ( .A(G134GAT), .B(n546), .ZN(G1343GAT) );
  NAND2_X1 U612 ( .A1(n547), .A2(n569), .ZN(n557) );
  NOR2_X1 U613 ( .A1(n571), .A2(n557), .ZN(n549) );
  XNOR2_X1 U614 ( .A(G141GAT), .B(KEYINPUT115), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n551) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(n554) );
  NOR2_X1 U619 ( .A1(n552), .A2(n557), .ZN(n553) );
  XOR2_X1 U620 ( .A(n554), .B(n553), .Z(G1345GAT) );
  NOR2_X1 U621 ( .A1(n555), .A2(n557), .ZN(n556) );
  XOR2_X1 U622 ( .A(G155GAT), .B(n556), .Z(G1346GAT) );
  NOR2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n560) );
  XNOR2_X1 U624 ( .A(G162GAT), .B(KEYINPUT117), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(G1347GAT) );
  XOR2_X1 U626 ( .A(G169GAT), .B(KEYINPUT121), .Z(n563) );
  NAND2_X1 U627 ( .A1(n566), .A2(n561), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(G1348GAT) );
  NAND2_X1 U629 ( .A1(n566), .A2(n580), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n567), .B(KEYINPUT58), .ZN(n568) );
  XNOR2_X1 U633 ( .A(n568), .B(G190GAT), .ZN(G1351GAT) );
  NAND2_X1 U634 ( .A1(n570), .A2(n569), .ZN(n584) );
  NOR2_X1 U635 ( .A1(n571), .A2(n584), .ZN(n576) );
  XOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n573) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(KEYINPUT59), .B(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n578) );
  INV_X1 U642 ( .A(n584), .ZN(n581) );
  NAND2_X1 U643 ( .A1(n581), .A2(n364), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XOR2_X1 U645 ( .A(G204GAT), .B(n579), .Z(G1353GAT) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(KEYINPUT126), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G211GAT), .B(n583), .ZN(G1354GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n587) );
  XNOR2_X1 U650 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

