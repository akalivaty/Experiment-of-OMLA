//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 0 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n187));
  XNOR2_X1  g001(.A(G128), .B(G143), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G122), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G116), .ZN(new_n192));
  INV_X1    g006(.A(G116), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G122), .ZN(new_n194));
  INV_X1    g008(.A(G107), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n192), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n193), .A2(KEYINPUT14), .A3(G122), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n192), .A2(new_n194), .ZN(new_n198));
  OAI211_X1 g012(.A(G107), .B(new_n197), .C1(new_n198), .C2(KEYINPUT14), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n190), .A2(new_n196), .A3(new_n199), .ZN(new_n200));
  XOR2_X1   g014(.A(KEYINPUT9), .B(G234), .Z(new_n201));
  XNOR2_X1  g015(.A(new_n201), .B(KEYINPUT79), .ZN(new_n202));
  INV_X1    g016(.A(G953), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(G217), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT87), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n188), .A2(KEYINPUT13), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  NOR3_X1   g022(.A1(new_n208), .A2(KEYINPUT13), .A3(G143), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(new_n189), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n207), .A2(new_n210), .B1(new_n189), .B2(new_n188), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n192), .A2(new_n194), .A3(new_n195), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n195), .B1(new_n192), .B2(new_n194), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT86), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n198), .A2(G107), .ZN(new_n216));
  AOI21_X1  g030(.A(KEYINPUT86), .B1(new_n216), .B2(new_n196), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n206), .B(new_n211), .C1(new_n215), .C2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n214), .B1(new_n212), .B2(new_n213), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n216), .A2(KEYINPUT86), .A3(new_n196), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n206), .B1(new_n222), .B2(new_n211), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n200), .B(new_n205), .C1(new_n219), .C2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT88), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n222), .A2(new_n211), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT87), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(new_n218), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n229), .A2(KEYINPUT88), .A3(new_n200), .A4(new_n205), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n200), .B1(new_n219), .B2(new_n223), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(new_n204), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n226), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G902), .ZN(new_n234));
  INV_X1    g048(.A(G478), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n235), .A2(KEYINPUT15), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n233), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n237), .B1(new_n233), .B2(new_n234), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n187), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n233), .A2(new_n234), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n236), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n233), .A2(new_n234), .A3(new_n237), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n242), .A2(KEYINPUT89), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(G113), .B(G122), .ZN(new_n246));
  INV_X1    g060(.A(G104), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n246), .B(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G140), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G125), .ZN(new_n250));
  INV_X1    g064(.A(G125), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G140), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n250), .A2(new_n252), .A3(KEYINPUT16), .ZN(new_n253));
  OR3_X1    g067(.A1(new_n251), .A2(KEYINPUT16), .A3(G140), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(G146), .ZN(new_n255));
  NOR2_X1   g069(.A1(G237), .A2(G953), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(G143), .A3(G214), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(G143), .B1(new_n256), .B2(G214), .ZN(new_n259));
  OAI21_X1  g073(.A(G131), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n259), .ZN(new_n261));
  INV_X1    g075(.A(G131), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(new_n262), .A3(new_n257), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(G125), .B(G140), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n265), .B(KEYINPUT19), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n255), .B(new_n264), .C1(new_n267), .C2(G146), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n261), .A2(new_n257), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(KEYINPUT18), .A3(G131), .ZN(new_n270));
  NAND2_X1  g084(.A1(KEYINPUT18), .A2(G131), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n261), .A2(new_n257), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G146), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n265), .B(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n270), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n248), .B1(new_n268), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n275), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT17), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n260), .A2(new_n263), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n269), .A2(KEYINPUT17), .A3(G131), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n255), .A2(KEYINPUT76), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n251), .A2(KEYINPUT16), .A3(G140), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n283), .B1(new_n265), .B2(KEYINPUT16), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT76), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n285), .A3(G146), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT77), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n253), .A2(new_n254), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n287), .B1(new_n288), .B2(new_n273), .ZN(new_n289));
  AOI211_X1 g103(.A(KEYINPUT77), .B(G146), .C1(new_n253), .C2(new_n254), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n282), .B(new_n286), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n281), .B1(new_n291), .B2(KEYINPUT85), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT77), .B1(new_n284), .B2(G146), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n288), .A2(new_n287), .A3(new_n273), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT85), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n295), .A2(new_n296), .A3(new_n282), .A4(new_n286), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n277), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n276), .B1(new_n298), .B2(new_n248), .ZN(new_n299));
  NOR2_X1   g113(.A1(G475), .A2(G902), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT20), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n291), .A2(KEYINPUT85), .ZN(new_n303));
  INV_X1    g117(.A(new_n281), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n297), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(new_n248), .A3(new_n275), .ZN(new_n306));
  INV_X1    g120(.A(new_n276), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT20), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n309), .A3(new_n300), .ZN(new_n310));
  INV_X1    g124(.A(new_n248), .ZN(new_n311));
  AOI211_X1 g125(.A(new_n311), .B(new_n277), .C1(new_n292), .C2(new_n297), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n248), .B1(new_n305), .B2(new_n275), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n234), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n302), .A2(new_n310), .B1(new_n314), .B2(G475), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n203), .A2(G952), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n316), .B1(G234), .B2(G237), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT21), .B(G898), .ZN(new_n318));
  XOR2_X1   g132(.A(new_n318), .B(KEYINPUT90), .Z(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  AOI211_X1 g134(.A(new_n234), .B(new_n203), .C1(G234), .C2(G237), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n317), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n315), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT91), .B1(new_n245), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n302), .A2(new_n310), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n314), .A2(G475), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n326), .A2(new_n323), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT91), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n328), .A2(new_n329), .A3(new_n244), .A4(new_n240), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G217), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n332), .B1(G234), .B2(new_n234), .ZN(new_n333));
  AND2_X1   g147(.A1(KEYINPUT66), .A2(G119), .ZN(new_n334));
  NOR2_X1   g148(.A1(KEYINPUT66), .A2(G119), .ZN(new_n335));
  OAI21_X1  g149(.A(G128), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G119), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n208), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT24), .B(G110), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n339), .A2(KEYINPUT75), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(KEYINPUT75), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n336), .B(new_n338), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT23), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n334), .A2(new_n335), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n343), .B1(new_n344), .B2(G128), .ZN(new_n345));
  INV_X1    g159(.A(G110), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n336), .A2(new_n338), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n345), .B(new_n346), .C1(new_n347), .C2(new_n343), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n342), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n342), .A2(new_n348), .A3(KEYINPUT78), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n265), .A2(new_n273), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n255), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n351), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n345), .B1(new_n347), .B2(new_n343), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n340), .A2(new_n341), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n356), .A2(G110), .B1(new_n357), .B2(new_n347), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n291), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT22), .B(G137), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n203), .A2(G221), .A3(G234), .ZN(new_n361));
  XOR2_X1   g175(.A(new_n360), .B(new_n361), .Z(new_n362));
  AND3_X1   g176(.A1(new_n355), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n362), .B1(new_n355), .B2(new_n359), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT25), .B1(new_n365), .B2(new_n234), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT25), .ZN(new_n367));
  NOR4_X1   g181(.A1(new_n363), .A2(new_n364), .A3(new_n367), .A4(G902), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n333), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n364), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n355), .A2(new_n359), .A3(new_n362), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n333), .A2(G902), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n369), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n256), .A2(G210), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(KEYINPUT27), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT26), .B(G101), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n377), .B(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT28), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n273), .A2(G143), .ZN(new_n382));
  INV_X1    g196(.A(G143), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G146), .ZN(new_n384));
  AND2_X1   g198(.A1(KEYINPUT0), .A2(G128), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n382), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(G143), .B(G146), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT0), .B(G128), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT11), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n391), .B1(new_n189), .B2(G137), .ZN(new_n392));
  INV_X1    g206(.A(G137), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(KEYINPUT11), .A3(G134), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n189), .A2(G137), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n392), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G131), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n392), .A2(new_n394), .A3(new_n262), .A4(new_n395), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n397), .A2(KEYINPUT70), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT70), .B1(new_n397), .B2(new_n398), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n390), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT67), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n402), .B1(new_n337), .B2(G116), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n193), .A2(KEYINPUT67), .A3(G119), .ZN(new_n404));
  AOI22_X1  g218(.A1(new_n344), .A2(G116), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G113), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT2), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT2), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G113), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT68), .B1(new_n405), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n403), .A2(new_n404), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT66), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n337), .ZN(new_n414));
  NAND2_X1  g228(.A1(KEYINPUT66), .A2(G119), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(G116), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT68), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n417), .A2(new_n418), .A3(new_n407), .A4(new_n409), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n412), .A2(new_n416), .A3(new_n410), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT69), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n412), .A2(new_n416), .A3(KEYINPUT69), .A4(new_n410), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n411), .A2(new_n419), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT1), .ZN(new_n425));
  AND4_X1   g239(.A1(new_n425), .A2(new_n382), .A3(new_n384), .A4(G128), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT1), .B1(new_n383), .B2(G146), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n427), .A2(G128), .B1(new_n382), .B2(new_n384), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n189), .A2(G137), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n393), .A2(G134), .ZN(new_n431));
  OAI21_X1  g245(.A(G131), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n398), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(KEYINPUT71), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n427), .A2(G128), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n382), .A2(new_n384), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n387), .A2(G128), .A3(new_n427), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT71), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n439), .A2(new_n440), .A3(new_n398), .A4(new_n432), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n401), .A2(new_n424), .A3(new_n434), .A4(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT65), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n433), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n398), .A2(new_n432), .A3(KEYINPUT65), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n439), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n389), .A2(KEYINPUT64), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n397), .A2(new_n398), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT64), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n386), .B(new_n449), .C1(new_n387), .C2(new_n388), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n447), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n411), .A2(new_n419), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n422), .A2(new_n423), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n381), .B1(new_n442), .B2(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n429), .A2(new_n433), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(KEYINPUT28), .B1(new_n459), .B2(new_n401), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n380), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n379), .A2(KEYINPUT72), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT30), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n446), .A2(new_n465), .A3(new_n451), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n401), .A2(new_n434), .A3(new_n441), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n466), .B1(new_n467), .B2(KEYINPUT30), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n442), .B(new_n464), .C1(new_n468), .C2(new_n424), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT31), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT70), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n448), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n397), .A2(KEYINPUT70), .A3(new_n398), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n389), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n434), .A2(new_n441), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT30), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n446), .A2(new_n451), .A3(new_n465), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n455), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n480), .A2(KEYINPUT31), .A3(new_n442), .A4(new_n464), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n462), .B1(new_n471), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(G472), .A2(G902), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT32), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n442), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n486), .B1(new_n479), .B2(new_n455), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT31), .B1(new_n487), .B2(new_n464), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n424), .B1(new_n477), .B2(new_n478), .ZN(new_n489));
  NOR4_X1   g303(.A1(new_n489), .A2(new_n486), .A3(new_n470), .A4(new_n463), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n461), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT32), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(new_n492), .A3(new_n483), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n485), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n379), .B1(new_n457), .B2(new_n460), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n442), .B(new_n380), .C1(new_n468), .C2(new_n424), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT29), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n434), .A2(new_n441), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT73), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n500), .A2(new_n501), .A3(new_n401), .A4(new_n424), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n475), .A2(new_n476), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n502), .B1(new_n424), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n442), .A2(KEYINPUT73), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT28), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n460), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n380), .A2(new_n498), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n507), .A2(KEYINPUT74), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n499), .A2(new_n234), .A3(new_n510), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n505), .B(new_n502), .C1(new_n424), .C2(new_n503), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n460), .B1(new_n512), .B2(KEYINPUT28), .ZN(new_n513));
  AOI21_X1  g327(.A(KEYINPUT74), .B1(new_n513), .B2(new_n509), .ZN(new_n514));
  OAI21_X1  g328(.A(G472), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n375), .B1(new_n494), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(G214), .B1(G237), .B2(G902), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT3), .B1(new_n247), .B2(G107), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT3), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n195), .A3(G104), .ZN(new_n521));
  INV_X1    g335(.A(G101), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n247), .A2(G107), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n519), .A2(new_n521), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n247), .A2(G107), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n195), .A2(G104), .ZN(new_n526));
  OAI21_X1  g340(.A(G101), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT5), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n344), .A2(new_n529), .A3(G116), .ZN(new_n530));
  OAI211_X1 g344(.A(G113), .B(new_n530), .C1(new_n417), .C2(new_n529), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n454), .A2(new_n528), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n519), .A2(new_n521), .A3(new_n523), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G101), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(KEYINPUT4), .A3(new_n524), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT4), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n533), .A2(new_n536), .A3(G101), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n532), .B1(new_n424), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(G110), .B(G122), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n532), .B(new_n540), .C1(new_n424), .C2(new_n538), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(KEYINPUT6), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT6), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n539), .A2(new_n545), .A3(new_n541), .ZN(new_n546));
  AOI21_X1  g360(.A(G125), .B1(new_n437), .B2(new_n438), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n386), .B(G125), .C1(new_n387), .C2(new_n388), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n203), .A2(G224), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n550), .B(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n544), .A2(new_n546), .A3(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n540), .B(KEYINPUT8), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n454), .A2(new_n528), .A3(new_n531), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n528), .B1(new_n454), .B2(new_n531), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT82), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT82), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n559), .B(new_n554), .C1(new_n555), .C2(new_n556), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n551), .A2(KEYINPUT83), .A3(KEYINPUT7), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n551), .A2(KEYINPUT7), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT83), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n548), .A2(new_n549), .A3(new_n561), .A4(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n549), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n563), .B(new_n562), .C1(new_n547), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n558), .A2(new_n543), .A3(new_n560), .A4(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n553), .A2(new_n234), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(G210), .B1(G237), .B2(G902), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n553), .A2(new_n234), .A3(new_n569), .A4(new_n571), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n518), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n575), .A2(KEYINPUT84), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT84), .ZN(new_n577));
  AOI211_X1 g391(.A(new_n577), .B(new_n518), .C1(new_n573), .C2(new_n574), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(G221), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n580), .B1(new_n202), .B2(new_n234), .ZN(new_n581));
  INV_X1    g395(.A(G469), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n524), .A2(new_n527), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n429), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n524), .B(new_n527), .C1(new_n426), .C2(new_n428), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n448), .A2(KEYINPUT12), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n474), .A2(new_n473), .B1(new_n584), .B2(new_n585), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n588), .B1(new_n589), .B2(KEYINPUT12), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT80), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n585), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT10), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT80), .B1(new_n528), .B2(new_n439), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT10), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n399), .A2(new_n400), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n535), .A2(new_n390), .A3(new_n537), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n593), .A2(new_n596), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(G110), .B(G140), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n203), .A2(G227), .ZN(new_n601));
  XOR2_X1   g415(.A(new_n600), .B(new_n601), .Z(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n590), .A2(new_n599), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n597), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n598), .B1(new_n594), .B2(new_n595), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n592), .A2(KEYINPUT10), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n603), .B1(new_n608), .B2(new_n599), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n582), .B(new_n234), .C1(new_n604), .C2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT81), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n608), .A2(new_n599), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n602), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n590), .A2(new_n599), .A3(new_n603), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT81), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n615), .A2(new_n616), .A3(new_n582), .A4(new_n234), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n603), .B1(new_n590), .B2(new_n599), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n599), .A2(new_n603), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n619), .B1(new_n620), .B2(new_n608), .ZN(new_n621));
  OAI21_X1  g435(.A(G469), .B1(new_n621), .B2(G902), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n581), .B1(new_n618), .B2(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n331), .A2(new_n516), .A3(new_n579), .A4(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G101), .ZN(G3));
  INV_X1    g439(.A(KEYINPUT92), .ZN(new_n626));
  INV_X1    g440(.A(new_n375), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n623), .ZN(new_n628));
  OAI21_X1  g442(.A(G472), .B1(new_n482), .B2(G902), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n491), .A2(new_n483), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n626), .B1(new_n628), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n631), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n633), .A2(KEYINPUT92), .A3(new_n627), .A4(new_n623), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n241), .A2(new_n235), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n233), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n232), .A2(KEYINPUT33), .A3(new_n224), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n234), .A2(G478), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n636), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n299), .A2(KEYINPUT20), .A3(new_n301), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n309), .B1(new_n308), .B2(new_n300), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n327), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n573), .A2(new_n574), .ZN(new_n647));
  AOI21_X1  g461(.A(KEYINPUT93), .B1(new_n647), .B2(new_n517), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT93), .ZN(new_n649));
  AOI211_X1 g463(.A(new_n649), .B(new_n518), .C1(new_n573), .C2(new_n574), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n323), .B(new_n646), .C1(new_n648), .C2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n635), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT34), .B(G104), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G6));
  AOI21_X1  g469(.A(new_n645), .B1(new_n244), .B2(new_n240), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n323), .B(new_n656), .C1(new_n648), .C2(new_n650), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(KEYINPUT94), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n657), .A2(KEYINPUT94), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n635), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT35), .B(G107), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  INV_X1    g476(.A(new_n333), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n367), .B1(new_n372), .B2(G902), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n365), .A2(KEYINPUT25), .A3(new_n234), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n355), .A2(new_n359), .ZN(new_n667));
  INV_X1    g481(.A(new_n362), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n668), .A2(KEYINPUT36), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n667), .B(new_n669), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n670), .A2(new_n373), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n631), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n331), .A2(new_n579), .A3(new_n673), .A4(new_n623), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT37), .B(G110), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G12));
  NAND2_X1  g490(.A1(new_n543), .A2(new_n568), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(KEYINPUT82), .B2(new_n557), .ZN(new_n678));
  AOI21_X1  g492(.A(G902), .B1(new_n678), .B2(new_n560), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n571), .B1(new_n679), .B2(new_n553), .ZN(new_n680));
  INV_X1    g494(.A(new_n574), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n517), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n649), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n575), .A2(KEYINPUT93), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n672), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(G900), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n317), .B1(new_n321), .B2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n656), .A2(new_n688), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n618), .A2(new_n622), .ZN(new_n691));
  INV_X1    g505(.A(new_n581), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n515), .B2(new_n494), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G128), .ZN(G30));
  NOR2_X1   g510(.A1(new_n487), .A2(new_n380), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n698), .B(new_n234), .C1(new_n512), .C2(new_n379), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(G472), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n494), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  XOR2_X1   g516(.A(new_n647), .B(KEYINPUT38), .Z(new_n703));
  AOI21_X1  g517(.A(new_n315), .B1(new_n240), .B2(new_n244), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n672), .A3(new_n517), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n687), .B(KEYINPUT39), .Z(new_n707));
  AND2_X1   g521(.A1(new_n623), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n709), .A2(KEYINPUT40), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(KEYINPUT40), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n706), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G143), .ZN(G45));
  NAND2_X1  g527(.A1(new_n494), .A2(new_n515), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n623), .ZN(new_n715));
  INV_X1    g529(.A(new_n672), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n642), .A2(new_n645), .A3(new_n688), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n716), .B(new_n717), .C1(new_n648), .C2(new_n650), .ZN(new_n718));
  OAI21_X1  g532(.A(KEYINPUT95), .B1(new_n715), .B2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT95), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n694), .A2(new_n685), .A3(new_n720), .A4(new_n717), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G146), .ZN(G48));
  OAI21_X1  g537(.A(new_n234), .B1(new_n604), .B2(new_n609), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(KEYINPUT96), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT96), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n726), .B(new_n234), .C1(new_n604), .C2(new_n609), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n725), .A2(G469), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n618), .A2(new_n728), .A3(new_n692), .ZN(new_n729));
  AOI211_X1 g543(.A(new_n375), .B(new_n729), .C1(new_n494), .C2(new_n515), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT97), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n652), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n729), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n714), .A2(new_n627), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(KEYINPUT97), .B1(new_n734), .B2(new_n651), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT41), .B(G113), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(KEYINPUT98), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n736), .B(new_n738), .ZN(G15));
  NAND2_X1  g553(.A1(new_n657), .A2(KEYINPUT94), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n683), .A2(new_n684), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT94), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n741), .A2(new_n742), .A3(new_n323), .A4(new_n656), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n734), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n193), .ZN(G18));
  INV_X1    g559(.A(KEYINPUT99), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n331), .A2(new_n714), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n733), .B(new_n716), .C1(new_n648), .C2(new_n650), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AOI22_X1  g563(.A1(new_n325), .A2(new_n330), .B1(new_n494), .B2(new_n515), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n750), .A2(KEYINPUT99), .A3(new_n685), .A4(new_n733), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G119), .ZN(G21));
  OAI22_X1  g567(.A1(new_n488), .A2(new_n490), .B1(new_n513), .B2(new_n379), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n483), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n629), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n375), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n729), .A2(new_n322), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n757), .A2(new_n741), .A3(new_n704), .A4(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G122), .ZN(G24));
  NAND3_X1  g574(.A1(new_n717), .A2(new_n629), .A3(new_n755), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n748), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(new_n251), .ZN(G27));
  NAND2_X1  g577(.A1(G469), .A2(G902), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(KEYINPUT100), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n765), .B1(new_n621), .B2(G469), .ZN(new_n766));
  AOI21_X1  g580(.A(G902), .B1(new_n613), .B2(new_n614), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n616), .B1(new_n767), .B2(new_n582), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n610), .A2(KEYINPUT81), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n766), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n692), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT101), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n581), .B1(new_n618), .B2(new_n766), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT101), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n573), .A2(new_n517), .A3(new_n574), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n773), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n778), .A2(KEYINPUT42), .A3(new_n516), .A4(new_n717), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n776), .B1(new_n771), .B2(new_n772), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n516), .A2(new_n780), .A3(new_n717), .A4(new_n775), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT42), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(new_n262), .ZN(G33));
  NAND4_X1  g599(.A1(new_n516), .A2(new_n780), .A3(new_n689), .A4(new_n775), .ZN(new_n786));
  XOR2_X1   g600(.A(KEYINPUT102), .B(G134), .Z(new_n787));
  XNOR2_X1  g601(.A(new_n786), .B(new_n787), .ZN(G36));
  AOI21_X1  g602(.A(KEYINPUT103), .B1(new_n642), .B2(new_n315), .ZN(new_n789));
  XOR2_X1   g603(.A(new_n789), .B(KEYINPUT43), .Z(new_n790));
  NAND3_X1  g604(.A1(new_n790), .A2(new_n631), .A3(new_n716), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT44), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n621), .A2(KEYINPUT45), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n621), .A2(KEYINPUT45), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(G469), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n765), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT46), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n798), .B1(new_n617), .B2(new_n611), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n796), .A2(KEYINPUT46), .A3(new_n797), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n581), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n707), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n793), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n791), .A2(new_n792), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n776), .B(KEYINPUT104), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G137), .ZN(G39));
  XNOR2_X1  g621(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n801), .B(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n717), .A2(new_n375), .A3(new_n777), .ZN(new_n810));
  OR3_X1    g624(.A1(new_n809), .A2(new_n714), .A3(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G140), .ZN(G42));
  NOR2_X1   g626(.A1(new_n756), .A2(new_n672), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n780), .A2(new_n813), .A3(new_n717), .A4(new_n775), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n238), .A2(new_n239), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n315), .A2(new_n815), .A3(new_n688), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n672), .A2(new_n816), .A3(new_n776), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n694), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n786), .A2(new_n814), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n783), .B2(new_n779), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n645), .A2(new_n815), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n579), .A2(KEYINPUT107), .A3(new_n323), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n682), .A2(new_n577), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n575), .A2(KEYINPUT84), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n823), .A2(new_n323), .A3(new_n824), .A4(new_n821), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT107), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n642), .A2(new_n645), .A3(KEYINPUT106), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT106), .B1(new_n642), .B2(new_n645), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n579), .A2(new_n830), .A3(new_n323), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n822), .A2(new_n827), .A3(new_n831), .ZN(new_n832));
  AOI22_X1  g646(.A1(new_n635), .A2(new_n832), .B1(new_n732), .B2(new_n735), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n624), .A2(new_n674), .A3(new_n759), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(new_n744), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n820), .A2(new_n833), .A3(new_n752), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT108), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n624), .A2(new_n674), .A3(new_n759), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n730), .B1(new_n659), .B2(new_n658), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n752), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT108), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n840), .A2(new_n841), .A3(new_n833), .A4(new_n820), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n762), .B1(new_n690), .B2(new_n694), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n774), .A2(new_n672), .A3(new_n688), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT109), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n844), .B(new_n845), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n741), .A2(new_n704), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n701), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n843), .A2(new_n848), .A3(new_n722), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n843), .A2(new_n848), .A3(new_n722), .A4(KEYINPUT52), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n837), .A2(new_n842), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT110), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n854), .A2(KEYINPUT110), .A3(new_n855), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n840), .A2(new_n833), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(new_n853), .A3(KEYINPUT53), .A4(new_n820), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n858), .A2(new_n859), .A3(new_n860), .A4(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n856), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n854), .A2(new_n855), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT54), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(KEYINPUT111), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT111), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n863), .A2(new_n869), .A3(new_n866), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n790), .A2(new_n317), .ZN(new_n871));
  INV_X1    g685(.A(new_n757), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n733), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n874), .B1(new_n683), .B2(new_n684), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n729), .A2(new_n776), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n702), .A2(new_n627), .A3(new_n317), .A4(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  AOI211_X1 g692(.A(new_n316), .B(new_n875), .C1(new_n646), .C2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n790), .A2(new_n317), .A3(new_n876), .ZN(new_n880));
  INV_X1    g694(.A(new_n516), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT48), .Z(new_n883));
  INV_X1    g697(.A(KEYINPUT112), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n703), .A2(new_n518), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n884), .B(KEYINPUT50), .C1(new_n874), .C2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT50), .ZN(new_n887));
  NOR4_X1   g701(.A1(new_n871), .A2(new_n729), .A3(new_n872), .A4(new_n885), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n887), .B1(new_n888), .B2(KEYINPUT112), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n618), .A2(new_n728), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n809), .B1(new_n692), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n892), .A2(new_n805), .A3(new_n873), .ZN(new_n893));
  INV_X1    g707(.A(new_n813), .ZN(new_n894));
  OR2_X1    g708(.A1(new_n642), .A2(new_n645), .ZN(new_n895));
  OAI22_X1  g709(.A1(new_n880), .A2(new_n894), .B1(new_n877), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n893), .A2(KEYINPUT51), .A3(new_n897), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n879), .B(new_n883), .C1(new_n890), .C2(new_n898), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n886), .A2(KEYINPUT113), .A3(new_n889), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT113), .B1(new_n886), .B2(new_n889), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n897), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(KEYINPUT114), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT114), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n904), .B(new_n897), .C1(new_n900), .C2(new_n901), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n903), .A2(new_n905), .A3(new_n893), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT51), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n899), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n868), .A2(new_n870), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT115), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT115), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n868), .A2(new_n911), .A3(new_n870), .A4(new_n908), .ZN(new_n912));
  OR2_X1    g726(.A1(G952), .A2(G953), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n910), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n891), .B(KEYINPUT49), .Z(new_n915));
  NAND2_X1  g729(.A1(new_n642), .A2(new_n315), .ZN(new_n916));
  NOR4_X1   g730(.A1(new_n375), .A2(new_n916), .A3(new_n581), .A4(new_n518), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n915), .A2(new_n702), .A3(new_n703), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n914), .A2(new_n918), .ZN(G75));
  NAND3_X1  g733(.A1(new_n858), .A2(new_n860), .A3(new_n862), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n920), .A2(G210), .A3(G902), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n921), .A2(KEYINPUT118), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(KEYINPUT118), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n544), .A2(new_n546), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT116), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT117), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT55), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(new_n552), .ZN(new_n928));
  XNOR2_X1  g742(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n922), .A2(new_n923), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n203), .A2(G952), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT56), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n921), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n932), .B1(new_n934), .B2(new_n928), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n931), .A2(new_n935), .ZN(G51));
  XNOR2_X1  g750(.A(new_n765), .B(KEYINPUT57), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n920), .A2(KEYINPUT54), .ZN(new_n938));
  INV_X1    g752(.A(new_n863), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n615), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n920), .A2(G902), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n942), .A2(new_n796), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n932), .B1(new_n941), .B2(new_n943), .ZN(G54));
  NAND2_X1  g758(.A1(KEYINPUT58), .A2(G475), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n299), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n932), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n942), .A2(new_n299), .A3(new_n945), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(G60));
  INV_X1    g764(.A(new_n640), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n868), .A2(new_n870), .ZN(new_n952));
  NAND2_X1  g766(.A1(G478), .A2(G902), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT59), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n951), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n951), .B(new_n954), .C1(new_n938), .C2(new_n939), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n947), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n955), .A2(new_n957), .ZN(G63));
  XNOR2_X1  g772(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n332), .A2(new_n234), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n920), .A2(new_n670), .A3(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n920), .A2(new_n961), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n947), .B(new_n962), .C1(new_n963), .C2(new_n365), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g779(.A(new_n203), .B1(new_n319), .B2(G224), .ZN(new_n966));
  INV_X1    g780(.A(new_n861), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n966), .B1(new_n967), .B2(new_n203), .ZN(new_n968));
  INV_X1    g782(.A(G898), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n925), .B1(new_n969), .B2(G953), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n968), .B(new_n970), .ZN(G69));
  NOR2_X1   g785(.A1(new_n709), .A2(new_n776), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n972), .B(new_n516), .C1(new_n821), .C2(new_n830), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT122), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n974), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n806), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT123), .Z(new_n978));
  AND2_X1   g792(.A1(new_n843), .A2(new_n722), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n712), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(KEYINPUT121), .B2(KEYINPUT62), .ZN(new_n981));
  XNOR2_X1  g795(.A(KEYINPUT121), .B(KEYINPUT62), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n979), .A2(new_n712), .A3(new_n982), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n978), .A2(new_n811), .A3(new_n981), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n203), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n479), .B(new_n267), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n986), .B1(G900), .B2(G953), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n801), .A2(new_n516), .A3(new_n707), .A4(new_n847), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n811), .A2(new_n806), .A3(new_n786), .A4(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n979), .ZN(new_n991));
  OR3_X1    g805(.A1(new_n990), .A2(new_n991), .A3(new_n784), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n988), .B1(new_n992), .B2(G953), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n987), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n203), .B1(G227), .B2(G900), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n995), .B1(new_n993), .B2(KEYINPUT124), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n994), .B(new_n996), .Z(G72));
  NAND2_X1  g811(.A1(G472), .A2(G902), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT63), .Z(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT125), .Z(new_n1000));
  OAI21_X1  g814(.A(new_n1000), .B1(new_n984), .B2(new_n967), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n932), .B1(new_n1001), .B2(new_n697), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n864), .A2(new_n865), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n496), .A2(new_n999), .ZN(new_n1004));
  OR3_X1    g818(.A1(new_n1003), .A2(new_n697), .A3(new_n1004), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1000), .B1(new_n992), .B2(new_n967), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n496), .B1(new_n1006), .B2(KEYINPUT126), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1007), .B1(KEYINPUT126), .B2(new_n1006), .ZN(new_n1008));
  AND3_X1   g822(.A1(new_n1002), .A2(new_n1005), .A3(new_n1008), .ZN(G57));
endmodule


