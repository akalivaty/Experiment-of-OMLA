//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 0 0 0 1 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1229, new_n1230,
    new_n1231, new_n1233, new_n1234, new_n1235, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  NOR2_X1   g0004(.A1(G58), .A2(G68), .ZN(new_n205));
  OR2_X1    g0005(.A1(new_n205), .A2(KEYINPUT65), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(KEYINPUT65), .ZN(new_n207));
  NAND3_X1  g0007(.A1(new_n206), .A2(G50), .A3(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G1), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n211), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT66), .Z(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n220));
  AND3_X1   g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n215), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT1), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n213), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G13), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n215), .A2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT64), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT0), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n224), .B(new_n230), .C1(new_n223), .C2(new_n222), .ZN(G361));
  XOR2_X1   g0031(.A(G250), .B(G257), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT67), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n235), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  XNOR2_X1  g0049(.A(KEYINPUT3), .B(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n250), .A2(G222), .A3(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G77), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n250), .A2(G1698), .ZN(new_n254));
  INV_X1    g0054(.A(G223), .ZN(new_n255));
  OAI221_X1 g0055(.A(new_n252), .B1(new_n253), .B2(new_n250), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  AND2_X1   g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(new_n210), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G274), .ZN(new_n260));
  AND2_X1   g0060(.A1(G1), .A2(G13), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G41), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT69), .B(G45), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n263), .B(new_n214), .C1(new_n264), .C2(G41), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT70), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G41), .A2(G45), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n266), .B1(new_n267), .B2(G1), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n214), .B(KEYINPUT70), .C1(G41), .C2(G45), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n258), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G226), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n259), .A2(new_n265), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G190), .ZN(new_n274));
  XOR2_X1   g0074(.A(new_n274), .B(KEYINPUT71), .Z(new_n275));
  NAND3_X1  g0075(.A1(new_n214), .A2(G13), .A3(G20), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G50), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n276), .A2(new_n210), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n214), .A2(G20), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G50), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n211), .B1(new_n205), .B2(new_n278), .ZN(new_n284));
  INV_X1    g0084(.A(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n211), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G150), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n211), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G58), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT8), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT8), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G58), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  AOI211_X1 g0095(.A(new_n284), .B(new_n288), .C1(new_n290), .C2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n280), .A2(new_n210), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  OAI221_X1 g0098(.A(new_n279), .B1(new_n281), .B2(new_n283), .C1(new_n296), .C2(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT9), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n272), .A2(G200), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT72), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n275), .A2(new_n303), .A3(new_n304), .A4(KEYINPUT10), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT10), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n306), .A2(KEYINPUT72), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(KEYINPUT72), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n274), .B(KEYINPUT71), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n308), .B(new_n309), .C1(new_n310), .C2(new_n302), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n272), .A2(new_n312), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n313), .B(new_n299), .C1(G179), .C2(new_n272), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n305), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n295), .A2(new_n282), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n317), .A2(new_n281), .B1(new_n276), .B2(new_n295), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT77), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n318), .B(new_n319), .ZN(new_n320));
  AND2_X1   g0120(.A1(KEYINPUT3), .A2(G33), .ZN(new_n321));
  NOR2_X1   g0121(.A1(KEYINPUT3), .A2(G33), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT7), .B1(new_n323), .B2(new_n211), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT7), .ZN(new_n325));
  NOR4_X1   g0125(.A1(new_n321), .A2(new_n322), .A3(new_n325), .A4(G20), .ZN(new_n326));
  OAI21_X1  g0126(.A(G68), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G68), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n291), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(G20), .B1(new_n329), .B2(new_n205), .ZN(new_n330));
  INV_X1    g0130(.A(new_n286), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G159), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n327), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT16), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n298), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n327), .A2(KEYINPUT16), .A3(new_n334), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n320), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G200), .ZN(new_n340));
  NOR2_X1   g0140(.A1(G223), .A2(G1698), .ZN(new_n341));
  INV_X1    g0141(.A(G226), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n341), .B1(new_n342), .B2(G1698), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n343), .A2(new_n250), .B1(G33), .B2(G87), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n261), .A2(new_n262), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n265), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G41), .ZN(new_n347));
  INV_X1    g0147(.A(G45), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(KEYINPUT70), .B1(new_n349), .B2(new_n214), .ZN(new_n350));
  NOR3_X1   g0150(.A1(new_n267), .A2(new_n266), .A3(G1), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n345), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(new_n237), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n340), .B1(new_n346), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n342), .A2(G1698), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(G223), .B2(G1698), .ZN(new_n356));
  INV_X1    g0156(.A(G87), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n356), .A2(new_n323), .B1(new_n285), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n258), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n270), .A2(G232), .ZN(new_n360));
  INV_X1    g0160(.A(G190), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n359), .A2(new_n360), .A3(new_n361), .A4(new_n265), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n354), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT78), .B1(new_n339), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n325), .B1(new_n250), .B2(G20), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n323), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n328), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n336), .B1(new_n367), .B2(new_n333), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n368), .A2(new_n338), .A3(new_n297), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n318), .B(KEYINPUT77), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n363), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT78), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT17), .B1(new_n364), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(G169), .B1(new_n346), .B2(new_n353), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n359), .A2(new_n360), .A3(G179), .A4(new_n265), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n369), .A2(new_n370), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g0177(.A(new_n377), .B(KEYINPUT18), .ZN(new_n378));
  AND3_X1   g0178(.A1(new_n363), .A2(new_n369), .A3(new_n370), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(KEYINPUT17), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n374), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n250), .A2(G232), .A3(new_n251), .ZN(new_n383));
  INV_X1    g0183(.A(G107), .ZN(new_n384));
  INV_X1    g0184(.A(G238), .ZN(new_n385));
  OAI221_X1 g0185(.A(new_n383), .B1(new_n384), .B2(new_n250), .C1(new_n254), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n258), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n270), .A2(G244), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n387), .A2(new_n265), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n312), .ZN(new_n390));
  INV_X1    g0190(.A(new_n295), .ZN(new_n391));
  OAI22_X1  g0191(.A1(new_n391), .A2(new_n286), .B1(new_n211), .B2(new_n253), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n357), .A2(KEYINPUT15), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT15), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G87), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n397), .A2(new_n289), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n297), .B1(new_n392), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n282), .A2(G77), .ZN(new_n400));
  OAI221_X1 g0200(.A(new_n399), .B1(G77), .B2(new_n276), .C1(new_n281), .C2(new_n400), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n390), .A2(new_n401), .ZN(new_n402));
  OR2_X1    g0202(.A1(new_n389), .A2(G179), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n401), .B1(G200), .B2(new_n389), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n361), .B2(new_n389), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n316), .A2(new_n382), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n277), .A2(new_n328), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n409), .B(KEYINPUT12), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n331), .A2(G50), .B1(G20), .B2(new_n328), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(new_n253), .B2(new_n289), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n412), .A2(KEYINPUT11), .A3(new_n297), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n282), .A2(G68), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n410), .B(new_n413), .C1(new_n281), .C2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT11), .B1(new_n412), .B2(new_n297), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n342), .A2(new_n251), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n237), .A2(G1698), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n419), .B(new_n420), .C1(new_n321), .C2(new_n322), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G33), .A2(G97), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AND2_X1   g0223(.A1(KEYINPUT69), .A2(G45), .ZN(new_n424));
  NOR2_X1   g0224(.A1(KEYINPUT69), .A2(G45), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(G1), .B1(new_n426), .B2(new_n347), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n258), .A2(new_n423), .B1(new_n427), .B2(new_n263), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT13), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT73), .ZN(new_n430));
  OAI21_X1  g0230(.A(G238), .B1(new_n270), .B2(new_n430), .ZN(new_n431));
  AOI211_X1 g0231(.A(KEYINPUT73), .B(new_n258), .C1(new_n268), .C2(new_n269), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n428), .B(new_n429), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n352), .A2(KEYINPUT73), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n270), .A2(new_n430), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(G238), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n429), .B1(new_n437), .B2(new_n428), .ZN(new_n438));
  OAI21_X1  g0238(.A(G169), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT14), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n428), .B1(new_n431), .B2(new_n432), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT13), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n433), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n444), .A2(KEYINPUT14), .A3(G169), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n429), .B1(new_n442), .B2(KEYINPUT74), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT74), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n437), .A2(new_n448), .A3(new_n428), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(G179), .A3(new_n433), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT76), .B1(new_n446), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT76), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n433), .A2(G179), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n454), .B1(new_n447), .B2(new_n449), .ZN(new_n455));
  AOI211_X1 g0255(.A(new_n453), .B(new_n455), .C1(new_n441), .C2(new_n445), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n418), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n444), .A2(G200), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n417), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n434), .A2(new_n361), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n450), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT75), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n450), .A2(new_n460), .A3(KEYINPUT75), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n459), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n457), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n408), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(G244), .B(new_n251), .C1(new_n321), .C2(new_n322), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT4), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n250), .A2(KEYINPUT4), .A3(G244), .A4(new_n251), .ZN(new_n472));
  NAND2_X1  g0272(.A1(G33), .A2(G283), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n250), .A2(G250), .A3(G1698), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n471), .A2(new_n472), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n258), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT79), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n348), .A2(G1), .ZN(new_n478));
  NAND2_X1  g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(KEYINPUT5), .A2(G41), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(G274), .B1(new_n257), .B2(new_n210), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n477), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n214), .A2(G45), .ZN(new_n485));
  OR2_X1    g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n485), .B1(new_n486), .B2(new_n479), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(KEYINPUT79), .A3(new_n263), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n487), .A2(new_n258), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n484), .A2(new_n488), .B1(new_n489), .B2(G257), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n476), .A2(new_n490), .A3(G190), .ZN(new_n491));
  INV_X1    g0291(.A(G97), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n277), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n285), .A2(G1), .ZN(new_n494));
  OR2_X1    g0294(.A1(new_n281), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n493), .B1(new_n495), .B2(new_n492), .ZN(new_n496));
  OAI21_X1  g0296(.A(G107), .B1(new_n324), .B2(new_n326), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT6), .ZN(new_n498));
  AND2_X1   g0298(.A1(G97), .A2(G107), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n498), .B1(new_n499), .B2(new_n202), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n384), .A2(KEYINPUT6), .A3(G97), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n502), .A2(G20), .B1(G77), .B2(new_n331), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n497), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n496), .B1(new_n504), .B2(new_n297), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n484), .A2(new_n488), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n489), .A2(G257), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT80), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n490), .A2(KEYINPUT80), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n510), .A2(new_n511), .B1(new_n258), .B2(new_n475), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n491), .B(new_n505), .C1(new_n512), .C2(new_n340), .ZN(new_n513));
  OAI211_X1 g0313(.A(G257), .B(G1698), .C1(new_n321), .C2(new_n322), .ZN(new_n514));
  OAI211_X1 g0314(.A(G250), .B(new_n251), .C1(new_n321), .C2(new_n322), .ZN(new_n515));
  INV_X1    g0315(.A(G294), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n514), .B(new_n515), .C1(new_n285), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n258), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n489), .A2(G264), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(new_n506), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(G179), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n520), .A2(new_n312), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n211), .B(G87), .C1(new_n321), .C2(new_n322), .ZN(new_n525));
  XNOR2_X1  g0325(.A(new_n525), .B(KEYINPUT22), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G116), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n527), .A2(G20), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT23), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n211), .B2(G107), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n384), .A2(KEYINPUT23), .A3(G20), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n526), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT24), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT24), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n526), .A2(new_n535), .A3(new_n532), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n298), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n495), .A2(new_n384), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n276), .A2(G107), .ZN(new_n539));
  XNOR2_X1  g0339(.A(KEYINPUT84), .B(KEYINPUT25), .ZN(new_n540));
  XNOR2_X1  g0340(.A(new_n539), .B(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n523), .B(new_n524), .C1(new_n537), .C2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n476), .A2(new_n490), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n505), .B1(new_n312), .B2(new_n545), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT80), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT80), .B1(new_n506), .B2(new_n507), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n522), .B(new_n476), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n513), .A2(new_n544), .A3(new_n550), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n526), .A2(new_n535), .A3(new_n532), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n535), .B1(new_n526), .B2(new_n532), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n297), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n520), .A2(G190), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n517), .A2(new_n258), .B1(new_n489), .B2(G264), .ZN(new_n556));
  AOI21_X1  g0356(.A(G200), .B1(new_n556), .B2(new_n506), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n554), .B(new_n542), .C1(new_n555), .C2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT81), .ZN(new_n559));
  OAI21_X1  g0359(.A(G250), .B1(new_n348), .B2(G1), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n559), .B1(new_n258), .B2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n345), .A2(KEYINPUT81), .A3(G250), .A4(new_n485), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n561), .A2(new_n562), .B1(new_n263), .B2(new_n478), .ZN(new_n563));
  OAI211_X1 g0363(.A(G244), .B(G1698), .C1(new_n321), .C2(new_n322), .ZN(new_n564));
  OAI211_X1 g0364(.A(G238), .B(new_n251), .C1(new_n321), .C2(new_n322), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n565), .A3(new_n527), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n258), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n522), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n396), .A2(new_n276), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n250), .A2(new_n211), .A3(G68), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT19), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n211), .B1(new_n422), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(G87), .B2(new_n203), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n572), .B1(new_n289), .B2(new_n492), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n571), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n570), .B1(new_n576), .B2(new_n297), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n397), .B2(new_n495), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n563), .A2(new_n567), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n312), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n569), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT82), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n579), .B2(new_n361), .ZN(new_n583));
  OR2_X1    g0383(.A1(new_n495), .A2(new_n357), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n577), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n563), .A2(new_n567), .A3(KEYINPUT82), .A4(G190), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n579), .A2(G200), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n583), .A2(new_n585), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n558), .A2(new_n581), .A3(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(G264), .B(G1698), .C1(new_n321), .C2(new_n322), .ZN(new_n590));
  OAI211_X1 g0390(.A(G257), .B(new_n251), .C1(new_n321), .C2(new_n322), .ZN(new_n591));
  INV_X1    g0391(.A(G303), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n590), .B(new_n591), .C1(new_n592), .C2(new_n250), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n258), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n489), .A2(G270), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n506), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G200), .ZN(new_n597));
  INV_X1    g0397(.A(G116), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n280), .A2(new_n210), .B1(G20), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(G20), .B1(G33), .B2(G283), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n285), .A2(G97), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT83), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT83), .B1(new_n600), .B2(new_n601), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n599), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT20), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(KEYINPUT20), .B(new_n599), .C1(new_n604), .C2(new_n605), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n495), .A2(G116), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n276), .A2(new_n598), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n608), .A2(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n597), .B(new_n612), .C1(new_n361), .C2(new_n596), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT21), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n596), .A2(G169), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n614), .B1(new_n615), .B2(new_n612), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n610), .A2(new_n611), .ZN(new_n617));
  XNOR2_X1  g0417(.A(new_n602), .B(new_n603), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT20), .B1(new_n618), .B2(new_n599), .ZN(new_n619));
  INV_X1    g0419(.A(new_n609), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n621), .A2(KEYINPUT21), .A3(G169), .A4(new_n596), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n594), .A2(new_n506), .A3(G179), .A4(new_n595), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n613), .A2(new_n616), .A3(new_n622), .A4(new_n625), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n551), .A2(new_n589), .A3(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n468), .A2(new_n627), .ZN(G372));
  OAI21_X1  g0428(.A(new_n457), .B1(new_n465), .B2(new_n404), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n339), .A2(KEYINPUT78), .A3(new_n363), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n371), .A2(new_n372), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n380), .B1(new_n632), .B2(KEYINPUT17), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n378), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n311), .B(new_n305), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n636), .A2(new_n314), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT85), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n588), .A2(new_n581), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n524), .B1(G179), .B2(new_n520), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n640), .B1(new_n554), .B2(new_n542), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n616), .A2(new_n622), .A3(new_n625), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n639), .B(new_n558), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n513), .A2(new_n550), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n638), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n644), .ZN(new_n646));
  INV_X1    g0446(.A(new_n589), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n544), .A2(new_n616), .A3(new_n625), .A4(new_n622), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n646), .A2(new_n647), .A3(KEYINPUT85), .A4(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n581), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n546), .A2(new_n549), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n651), .A2(new_n639), .A3(KEYINPUT26), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT26), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n588), .A2(new_n581), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n653), .B1(new_n550), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n650), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n645), .A2(new_n649), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n468), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n637), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n659), .B(KEYINPUT86), .ZN(G369));
  NAND3_X1  g0460(.A1(new_n214), .A2(new_n211), .A3(G13), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G213), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n537), .B2(new_n543), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n641), .B1(new_n558), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n544), .A2(new_n666), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n666), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n642), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(new_n669), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n612), .A2(new_n671), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n642), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n626), .B2(new_n677), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(G330), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n670), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n676), .A2(new_n682), .ZN(G399));
  NAND2_X1  g0483(.A1(new_n644), .A2(KEYINPUT90), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT90), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n513), .A2(new_n550), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n656), .B1(new_n687), .B2(new_n643), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n688), .A2(KEYINPUT29), .A3(new_n671), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT29), .B1(new_n657), .B2(new_n671), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n666), .A2(KEYINPUT31), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT88), .B1(new_n512), .B2(new_n521), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n476), .B1(new_n547), .B2(new_n548), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT88), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(new_n696), .A3(new_n520), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n596), .A2(new_n522), .A3(new_n579), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n694), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n568), .A2(new_n556), .A3(new_n476), .A4(new_n490), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n701), .B1(new_n702), .B2(new_n623), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n556), .A2(new_n567), .A3(new_n563), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n476), .A2(new_n490), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n704), .A2(new_n705), .A3(new_n624), .A4(KEYINPUT30), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n693), .B1(new_n700), .B2(new_n707), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n708), .A2(KEYINPUT89), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n627), .A2(new_n671), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT31), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n703), .A2(new_n706), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n695), .A2(new_n520), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n698), .B1(new_n713), .B2(KEYINPUT88), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n712), .B1(new_n714), .B2(new_n697), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n711), .B1(new_n715), .B2(new_n671), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n708), .A2(KEYINPUT89), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n709), .A2(new_n710), .A3(new_n716), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G330), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n692), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n214), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n226), .A2(G41), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(G1), .A3(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(new_n208), .B2(new_n723), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT87), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT28), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n721), .A2(new_n728), .ZN(G364));
  NOR2_X1   g0529(.A1(new_n225), .A2(G20), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n214), .B1(new_n730), .B2(G45), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OR3_X1    g0532(.A1(new_n722), .A2(new_n732), .A3(KEYINPUT91), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT91), .B1(new_n722), .B2(new_n732), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n681), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(G330), .B2(new_n679), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n226), .A2(new_n323), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G355), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(G116), .B2(new_n227), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n226), .A2(new_n250), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n743), .B1(new_n209), .B2(new_n426), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n248), .A2(G45), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n741), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G13), .A2(G33), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n210), .B1(G20), .B2(new_n312), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n736), .B1(new_n746), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n340), .A2(G179), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n754), .A2(G20), .A3(G190), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n357), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G179), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G190), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n323), .B(new_n756), .C1(G97), .C2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n757), .A2(G20), .A3(new_n361), .ZN(new_n761));
  INV_X1    g0561(.A(G159), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT32), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n754), .A2(G20), .A3(new_n361), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n765), .A2(KEYINPUT93), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(KEYINPUT93), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n760), .B(new_n764), .C1(new_n384), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(G20), .A2(G179), .ZN(new_n770));
  XOR2_X1   g0570(.A(new_n770), .B(KEYINPUT92), .Z(new_n771));
  NAND3_X1  g0571(.A1(new_n771), .A2(new_n361), .A3(G200), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AND3_X1   g0573(.A1(new_n771), .A2(G190), .A3(new_n340), .ZN(new_n774));
  AOI22_X1  g0574(.A1(G68), .A2(new_n773), .B1(new_n774), .B2(G58), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n771), .A2(G190), .A3(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n771), .A2(new_n361), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(G200), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n775), .B1(new_n278), .B2(new_n776), .C1(new_n253), .C2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n776), .ZN(new_n781));
  AOI22_X1  g0581(.A1(G326), .A2(new_n781), .B1(new_n774), .B2(G322), .ZN(new_n782));
  INV_X1    g0582(.A(G311), .ZN(new_n783));
  XOR2_X1   g0583(.A(KEYINPUT33), .B(G317), .Z(new_n784));
  OAI221_X1 g0584(.A(new_n782), .B1(new_n783), .B2(new_n779), .C1(new_n772), .C2(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n323), .B1(new_n755), .B2(new_n592), .ZN(new_n786));
  INV_X1    g0586(.A(new_n761), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n786), .B1(G329), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n759), .ZN(new_n789));
  INV_X1    g0589(.A(G283), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n788), .B1(new_n516), .B2(new_n789), .C1(new_n790), .C2(new_n768), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n769), .A2(new_n780), .B1(new_n785), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n753), .B1(new_n792), .B2(new_n750), .ZN(new_n793));
  INV_X1    g0593(.A(new_n749), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n793), .B1(new_n679), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n738), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(G396));
  NOR2_X1   g0597(.A1(new_n750), .A2(new_n747), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n735), .B1(new_n253), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n750), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n778), .A2(G159), .B1(new_n774), .B2(G143), .ZN(new_n801));
  INV_X1    g0601(.A(G137), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n801), .B1(new_n802), .B2(new_n776), .C1(new_n287), .C2(new_n772), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT34), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n789), .A2(new_n291), .ZN(new_n805));
  INV_X1    g0605(.A(G132), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n250), .B1(new_n761), .B2(new_n806), .C1(new_n755), .C2(new_n278), .ZN(new_n807));
  INV_X1    g0607(.A(new_n768), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n805), .B(new_n807), .C1(new_n808), .C2(G68), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G283), .A2(new_n773), .B1(new_n781), .B2(G303), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n598), .B2(new_n779), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT94), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n808), .A2(G87), .ZN(new_n813));
  AOI22_X1  g0613(.A1(G311), .A2(new_n787), .B1(new_n759), .B2(G97), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n323), .B1(new_n755), .B2(new_n384), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT95), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(G294), .B2(new_n774), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n804), .A2(new_n809), .B1(new_n812), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n401), .A2(new_n666), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n407), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(KEYINPUT96), .B1(new_n404), .B2(new_n671), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT96), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n402), .A2(new_n823), .A3(new_n403), .A4(new_n666), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n799), .B1(new_n800), .B2(new_n819), .C1(new_n826), .C2(new_n748), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n657), .A2(new_n671), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(new_n826), .ZN(new_n830));
  INV_X1    g0630(.A(new_n719), .ZN(new_n831));
  AND3_X1   g0631(.A1(new_n830), .A2(KEYINPUT97), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(KEYINPUT97), .B1(new_n830), .B2(new_n831), .ZN(new_n833));
  OR3_X1    g0633(.A1(new_n832), .A2(new_n833), .A3(new_n736), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n834), .A2(KEYINPUT98), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n830), .A2(new_n831), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n834), .B2(KEYINPUT98), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n828), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(G384));
  NAND2_X1  g0639(.A1(new_n468), .A2(new_n691), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n637), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n657), .A2(new_n671), .A3(new_n826), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n404), .A2(new_n666), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n418), .A2(new_n666), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n457), .A2(new_n466), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT14), .B1(new_n444), .B2(G169), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n440), .B(new_n312), .C1(new_n443), .C2(new_n433), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n451), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n453), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n446), .A2(KEYINPUT76), .A3(new_n451), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n418), .B(new_n666), .C1(new_n853), .C2(new_n465), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n847), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n845), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT38), .ZN(new_n857));
  INV_X1    g0657(.A(new_n318), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n369), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n664), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(new_n633), .B2(new_n378), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n364), .A2(new_n373), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n664), .B1(new_n369), .B2(new_n370), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n377), .A2(new_n864), .A3(KEYINPUT37), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n375), .A2(new_n376), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n859), .B1(new_n866), .B2(new_n860), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n630), .A2(new_n631), .A3(new_n867), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n863), .A2(new_n865), .B1(new_n868), .B2(KEYINPUT37), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n857), .B1(new_n862), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(KEYINPUT37), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n865), .A2(new_n631), .A3(new_n630), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g0673(.A(KEYINPUT38), .B(new_n873), .C1(new_n382), .C2(new_n861), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  OAI22_X1  g0676(.A1(new_n856), .A2(new_n876), .B1(new_n378), .B2(new_n860), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n457), .A2(new_n666), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT100), .ZN(new_n881));
  INV_X1    g0681(.A(new_n377), .ZN(new_n882));
  INV_X1    g0682(.A(new_n864), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n882), .A2(new_n883), .A3(new_n371), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT37), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT99), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n885), .A2(new_n886), .B1(new_n863), .B2(new_n865), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n884), .A2(KEYINPUT99), .A3(KEYINPUT37), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n374), .A2(new_n378), .A3(new_n381), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n887), .A2(new_n888), .B1(new_n889), .B2(new_n864), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n881), .B1(new_n890), .B2(KEYINPUT38), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(new_n864), .ZN(new_n892));
  NOR3_X1   g0692(.A1(new_n379), .A2(new_n377), .A3(new_n864), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT37), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n886), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(new_n872), .A3(new_n888), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(KEYINPUT100), .A3(new_n857), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n891), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT39), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n874), .A2(new_n900), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n899), .A2(new_n901), .B1(KEYINPUT39), .B2(new_n875), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n878), .B1(new_n880), .B2(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n841), .B(new_n903), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n407), .A2(new_n820), .B1(new_n822), .B2(new_n824), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT101), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n715), .B2(new_n671), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n700), .A2(new_n707), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(KEYINPUT101), .A3(new_n666), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n907), .A2(new_n711), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n708), .B1(new_n627), .B2(new_n671), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n905), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n855), .A2(KEYINPUT40), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT100), .B1(new_n897), .B2(new_n857), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n881), .B(KEYINPUT38), .C1(new_n892), .C2(new_n896), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n874), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n855), .A2(new_n875), .A3(new_n912), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT40), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n913), .A2(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n910), .A2(new_n911), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n468), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(G330), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n920), .B2(new_n922), .ZN(new_n924));
  OAI22_X1  g0724(.A1(new_n904), .A2(new_n924), .B1(new_n214), .B2(new_n730), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n904), .B2(new_n924), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n502), .A2(KEYINPUT35), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n502), .A2(KEYINPUT35), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n927), .A2(G116), .A3(new_n212), .A4(new_n928), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT36), .Z(new_n930));
  OR3_X1    g0730(.A1(new_n208), .A2(new_n253), .A3(new_n329), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n278), .A2(G68), .ZN(new_n932));
  AOI211_X1 g0732(.A(new_n214), .B(G13), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  OR3_X1    g0733(.A1(new_n926), .A2(new_n930), .A3(new_n933), .ZN(G367));
  INV_X1    g0734(.A(KEYINPUT42), .ZN(new_n935));
  INV_X1    g0735(.A(new_n687), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n505), .A2(new_n671), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n651), .A2(new_n666), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n935), .B1(new_n940), .B2(new_n675), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n936), .A2(new_n641), .A3(new_n937), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n666), .B1(new_n942), .B2(new_n550), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(KEYINPUT104), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT104), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n941), .B2(new_n943), .ZN(new_n947));
  INV_X1    g0747(.A(new_n940), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n948), .A2(new_n674), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n935), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n945), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n585), .A2(new_n671), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT102), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n639), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n954), .B(KEYINPUT103), .C1(new_n581), .C2(new_n953), .ZN(new_n955));
  OR3_X1    g0755(.A1(new_n953), .A2(KEYINPUT103), .A3(new_n581), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT43), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n955), .A2(KEYINPUT43), .A3(new_n956), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n951), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n944), .A2(KEYINPUT104), .B1(new_n935), .B2(new_n949), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n962), .A2(new_n958), .A3(new_n957), .A4(new_n947), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n948), .A2(new_n682), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n961), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(KEYINPUT106), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT106), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n961), .A2(new_n963), .A3(new_n967), .A4(new_n964), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n964), .B1(new_n961), .B2(new_n963), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n969), .B1(KEYINPUT105), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n970), .A2(KEYINPUT105), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n972), .A2(new_n966), .A3(new_n968), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n722), .B(KEYINPUT41), .Z(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n676), .A2(new_n940), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT45), .Z(new_n977));
  INV_X1    g0777(.A(new_n682), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(KEYINPUT108), .ZN(new_n979));
  NOR2_X1   g0779(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n980));
  OR3_X1    g0780(.A1(new_n676), .A2(new_n940), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n980), .B1(new_n676), .B2(new_n940), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AND3_X1   g0784(.A1(new_n977), .A2(new_n979), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n979), .B1(new_n977), .B2(new_n984), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n670), .B(new_n673), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n680), .A2(KEYINPUT109), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n987), .B(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n692), .A2(new_n989), .A3(new_n719), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n985), .A2(new_n986), .A3(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n975), .B1(new_n991), .B2(new_n720), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n731), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n971), .A2(new_n973), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n957), .A2(new_n749), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n235), .A2(new_n743), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n752), .B1(new_n226), .B2(new_n396), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n735), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n755), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(G116), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT46), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT110), .Z(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G311), .B2(new_n781), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n774), .A2(G303), .ZN(new_n1005));
  INV_X1    g0805(.A(G317), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n323), .B1(new_n1006), .B2(new_n761), .C1(new_n789), .C2(new_n384), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n768), .A2(new_n492), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1007), .B(new_n1008), .C1(new_n1001), .C2(new_n1000), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(G283), .A2(new_n778), .B1(new_n773), .B2(G294), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1004), .A2(new_n1005), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n774), .ZN(new_n1012));
  INV_X1    g0812(.A(G143), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n1012), .A2(new_n287), .B1(new_n1013), .B2(new_n776), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(G159), .B2(new_n773), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n323), .B1(new_n808), .B2(G77), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1016), .A2(KEYINPUT111), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(KEYINPUT111), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n999), .A2(G58), .B1(new_n787), .B2(G137), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n328), .B2(new_n789), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G50), .B2(new_n778), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1015), .A2(new_n1017), .A3(new_n1018), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1011), .A2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n995), .B(new_n998), .C1(new_n800), .C2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n994), .A2(new_n1026), .ZN(G387));
  NAND2_X1  g0827(.A1(new_n989), .A2(new_n732), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G68), .A2(new_n778), .B1(new_n781), .B2(G159), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n295), .A2(new_n773), .B1(new_n774), .B2(G50), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1008), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n250), .B1(new_n761), .B2(new_n287), .C1(new_n755), .C2(new_n253), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(new_n396), .B2(new_n759), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n250), .B1(new_n787), .B2(G326), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n789), .A2(new_n790), .B1(new_n755), .B2(new_n516), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n778), .A2(G303), .B1(new_n774), .B2(G317), .ZN(new_n1037));
  INV_X1    g0837(.A(G322), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1037), .B1(new_n783), .B2(new_n772), .C1(new_n1038), .C2(new_n776), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT48), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1036), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n1040), .B2(new_n1039), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT49), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1035), .B1(new_n598), .B2(new_n768), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1034), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n800), .B1(new_n1046), .B2(KEYINPUT113), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(KEYINPUT113), .B2(new_n1046), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n240), .A2(new_n426), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n724), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1049), .A2(new_n742), .B1(new_n1050), .B2(new_n739), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n724), .B(new_n348), .C1(new_n328), .C2(new_n253), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT50), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n391), .B2(G50), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n295), .A2(KEYINPUT50), .A3(new_n278), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1052), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n1051), .A2(new_n1056), .B1(G107), .B2(new_n227), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n735), .B1(new_n1057), .B2(new_n751), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1048), .B(new_n1058), .C1(new_n670), .C2(new_n794), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n990), .A2(new_n722), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n989), .B1(new_n692), .B2(new_n719), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1028), .B(new_n1059), .C1(new_n1060), .C2(new_n1061), .ZN(G393));
  NOR2_X1   g0862(.A1(new_n991), .A2(new_n723), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n990), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n977), .A2(new_n984), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(new_n682), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1063), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n732), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n245), .A2(new_n743), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n751), .B1(new_n492), .B2(new_n227), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n773), .A2(G303), .B1(G116), .B2(new_n759), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(KEYINPUT116), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n755), .A2(new_n790), .B1(new_n1038), .B2(new_n761), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT115), .Z(new_n1075));
  OAI211_X1 g0875(.A(new_n1075), .B(new_n323), .C1(new_n384), .C2(new_n768), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1071), .A2(KEYINPUT116), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n779), .A2(new_n516), .ZN(new_n1078));
  NOR4_X1   g0878(.A1(new_n1073), .A2(new_n1076), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n1012), .A2(new_n783), .B1(new_n1006), .B2(new_n776), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT52), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n1012), .A2(new_n762), .B1(new_n287), .B2(new_n776), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT51), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n295), .A2(new_n778), .B1(new_n773), .B2(G50), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n323), .B1(new_n759), .B2(G77), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n755), .A2(new_n328), .B1(new_n1013), .B2(new_n761), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT114), .Z(new_n1087));
  AND4_X1   g0887(.A1(new_n813), .A2(new_n1084), .A3(new_n1085), .A4(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1079), .A2(new_n1081), .B1(new_n1083), .B2(new_n1088), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n736), .B1(new_n1069), .B2(new_n1070), .C1(new_n1089), .C2(new_n800), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT117), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n794), .B2(new_n940), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1067), .A2(new_n1068), .A3(new_n1092), .ZN(G390));
  AND3_X1   g0893(.A1(new_n718), .A2(G330), .A3(new_n826), .ZN(new_n1094));
  OAI21_X1  g0894(.A(KEYINPUT118), .B1(new_n1094), .B2(new_n855), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n855), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT118), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1096), .B(new_n1097), .C1(new_n719), .C2(new_n905), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n855), .A2(new_n912), .A3(G330), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1095), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n845), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n688), .A2(new_n826), .A3(new_n671), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n844), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n1094), .B2(new_n855), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n912), .A2(G330), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n1096), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1101), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n468), .A2(G330), .A3(new_n921), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n637), .A2(new_n840), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n879), .B1(new_n1103), .B2(new_n855), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n916), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1094), .A2(new_n855), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n901), .B1(new_n914), .B2(new_n915), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n875), .A2(KEYINPUT39), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n879), .B1(new_n845), .B2(new_n855), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1113), .B(new_n1114), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n856), .A2(new_n880), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n902), .A2(new_n1120), .B1(new_n916), .B2(new_n1112), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1119), .B1(new_n1121), .B2(new_n1099), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n1111), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n723), .B1(new_n1111), .B2(new_n1122), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  OR2_X1    g0925(.A1(new_n1122), .A2(new_n731), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n250), .B(new_n756), .C1(G294), .C2(new_n787), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n1127), .B1(new_n328), .B2(new_n768), .C1(new_n253), .C2(new_n789), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(G107), .A2(new_n773), .B1(new_n774), .B2(G116), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n492), .B2(new_n779), .C1(new_n790), .C2(new_n776), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(G128), .A2(new_n781), .B1(new_n774), .B2(G132), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT54), .B(G143), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n1131), .B1(new_n802), .B2(new_n772), .C1(new_n779), .C2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n789), .A2(new_n762), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n323), .B(new_n1134), .C1(G125), .C2(new_n787), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n755), .A2(new_n287), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT53), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1135), .B(new_n1137), .C1(new_n278), .C2(new_n768), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n1128), .A2(new_n1130), .B1(new_n1133), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n750), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n735), .B1(new_n391), .B2(new_n798), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1140), .B(new_n1141), .C1(new_n1117), .C2(new_n748), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1125), .A2(new_n1126), .A3(new_n1142), .ZN(G378));
  NAND2_X1  g0943(.A1(new_n913), .A2(new_n916), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n315), .A2(new_n299), .A3(new_n860), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n299), .A2(new_n860), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n305), .A2(new_n311), .A3(new_n314), .A4(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1145), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n917), .A2(new_n918), .ZN(new_n1154));
  AND4_X1   g0954(.A1(G330), .A2(new_n1144), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1153), .B1(new_n919), .B2(G330), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n903), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1144), .A2(G330), .A3(new_n1154), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1153), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n877), .B1(new_n879), .B2(new_n1117), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n919), .A2(G330), .A3(new_n1153), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1157), .A2(new_n1163), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1100), .A2(new_n845), .B1(new_n1106), .B2(new_n1104), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1110), .B1(new_n1122), .B2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1164), .A2(new_n1166), .A3(KEYINPUT57), .ZN(new_n1167));
  AOI21_X1  g0967(.A(KEYINPUT57), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n722), .B(new_n1167), .C1(new_n1168), .C2(KEYINPUT119), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT119), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1170), .B(KEYINPUT57), .C1(new_n1164), .C2(new_n1166), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1153), .A2(new_n748), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n735), .B1(new_n278), .B2(new_n798), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n789), .A2(new_n287), .B1(new_n1132), .B2(new_n755), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(G125), .A2(new_n781), .B1(new_n774), .B2(G128), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n802), .B2(new_n779), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1175), .B(new_n1177), .C1(G132), .C2(new_n773), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT59), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n808), .A2(G159), .ZN(new_n1182));
  AOI211_X1 g0982(.A(G33), .B(G41), .C1(new_n787), .C2(G124), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n779), .A2(new_n397), .B1(new_n492), .B2(new_n772), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n1012), .A2(new_n384), .B1(new_n598), .B2(new_n776), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n768), .A2(new_n291), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n323), .A2(new_n347), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n999), .B2(G77), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(new_n328), .B2(new_n789), .C1(new_n790), .C2(new_n761), .ZN(new_n1190));
  NOR4_X1   g0990(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .A4(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(KEYINPUT58), .ZN(new_n1192));
  OR2_X1    g0992(.A1(new_n1191), .A2(KEYINPUT58), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1188), .B(new_n278), .C1(G33), .C2(G41), .ZN(new_n1194));
  AND4_X1   g0994(.A1(new_n1184), .A2(new_n1192), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1174), .B1(new_n1195), .B2(new_n800), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1173), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n1164), .B2(new_n732), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1172), .A2(new_n1198), .ZN(G375));
  INV_X1    g0999(.A(new_n1110), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n1165), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1201), .A2(new_n975), .A3(new_n1111), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT120), .B1(new_n1096), .B2(new_n747), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1096), .A2(KEYINPUT120), .A3(new_n747), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n806), .A2(new_n776), .B1(new_n772), .B2(new_n1132), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G137), .B2(new_n774), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT122), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n250), .B1(new_n755), .B2(new_n762), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G128), .B2(new_n787), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n278), .B2(new_n789), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1187), .B(new_n1210), .C1(G150), .C2(new_n778), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1207), .A2(new_n1211), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n779), .A2(new_n384), .B1(new_n598), .B2(new_n772), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G283), .B2(new_n774), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n999), .A2(G97), .B1(new_n787), .B2(G303), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n397), .B2(new_n789), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G294), .B2(new_n781), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n808), .A2(G77), .ZN(new_n1218));
  AOI21_X1  g1018(.A(KEYINPUT121), .B1(new_n1218), .B2(new_n323), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1218), .A2(KEYINPUT121), .A3(new_n323), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1214), .B(new_n1217), .C1(new_n1219), .C2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n800), .B1(new_n1212), .B2(new_n1221), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n735), .B(new_n1222), .C1(new_n328), .C2(new_n798), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1223), .B(KEYINPUT123), .Z(new_n1224));
  NAND2_X1  g1024(.A1(new_n1204), .A2(new_n1224), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n1165), .A2(new_n731), .B1(new_n1203), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1202), .A2(new_n1227), .ZN(G381));
  OR2_X1    g1028(.A1(G393), .A2(G396), .ZN(new_n1229));
  OR2_X1    g1029(.A1(G390), .A2(new_n1229), .ZN(new_n1230));
  OR4_X1    g1030(.A1(G384), .A2(new_n1230), .A3(G378), .A4(G381), .ZN(new_n1231));
  OR3_X1    g1031(.A1(new_n1231), .A2(G387), .A3(G375), .ZN(G407));
  NAND2_X1  g1032(.A1(new_n665), .A2(G213), .ZN(new_n1233));
  XOR2_X1   g1033(.A(new_n1233), .B(KEYINPUT124), .Z(new_n1234));
  OR3_X1    g1034(.A1(G375), .A2(G378), .A3(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(G407), .A2(G213), .A3(new_n1235), .ZN(G409));
  INV_X1    g1036(.A(G390), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(G387), .A2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n994), .A2(G390), .A3(new_n1026), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(G393), .B(new_n796), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT125), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1238), .A2(new_n1239), .A3(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1240), .A2(KEYINPUT125), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(G378), .B(new_n1198), .C1(new_n1169), .C2(new_n1171), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1126), .A2(new_n1142), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1164), .A2(new_n975), .A3(new_n1166), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1198), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1248), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1246), .A2(new_n1251), .B1(G213), .B2(new_n665), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1111), .A2(KEYINPUT60), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1201), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1200), .A2(KEYINPUT60), .A3(new_n1165), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1255), .A2(new_n722), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1226), .B(new_n838), .C1(new_n1254), .C2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1254), .ZN(new_n1258));
  AOI21_X1  g1058(.A(G384), .B1(new_n1258), .B2(new_n1227), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT62), .B1(new_n1252), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1246), .A2(new_n1251), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1234), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT126), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1262), .A2(KEYINPUT126), .A3(new_n1234), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1260), .A2(KEYINPUT62), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1261), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(G2897), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1233), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1260), .A2(new_n1271), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n1257), .A2(new_n1259), .B1(new_n1270), .B2(new_n1234), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1265), .A2(new_n1266), .A3(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT61), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1245), .B1(new_n1269), .B2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1252), .B1(new_n1273), .B2(new_n1272), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1245), .A2(new_n1279), .A3(KEYINPUT61), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1267), .A2(KEYINPUT63), .A3(new_n1260), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1252), .A2(new_n1260), .ZN(new_n1282));
  OR2_X1    g1082(.A1(new_n1282), .A2(KEYINPUT63), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1280), .A2(new_n1281), .A3(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1278), .A2(new_n1284), .ZN(G405));
  NOR2_X1   g1085(.A1(new_n1260), .A2(KEYINPUT127), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(G375), .A2(new_n1248), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1286), .B1(new_n1246), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1260), .A2(KEYINPUT127), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1287), .A2(new_n1260), .A3(KEYINPUT127), .A4(new_n1246), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  OR2_X1    g1092(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1290), .A2(new_n1245), .A3(new_n1291), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(G402));
endmodule


