//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 1 0 1 1 1 1 1 1 1 0 1 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n774, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963;
  AND2_X1   g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT41), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G134gat), .ZN(new_n204));
  INV_X1    g003(.A(G162gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G190gat), .B(G218gat), .Z(new_n207));
  XNOR2_X1  g006(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT89), .B(KEYINPUT17), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n211));
  NOR3_X1   g010(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n212), .A2(KEYINPUT88), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT88), .ZN(new_n214));
  NOR4_X1   g013(.A1(new_n214), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n211), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G29gat), .A2(G36gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(G43gat), .B(G50gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT15), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n218), .A2(KEYINPUT15), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n216), .A2(new_n217), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n219), .ZN(new_n222));
  INV_X1    g021(.A(new_n211), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n217), .B1(new_n223), .B2(new_n212), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n210), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n221), .A2(new_n225), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n226), .B1(KEYINPUT17), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G85gat), .A2(G92gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT7), .ZN(new_n230));
  NAND2_X1  g029(.A1(G99gat), .A2(G106gat), .ZN(new_n231));
  INV_X1    g030(.A(G85gat), .ZN(new_n232));
  INV_X1    g031(.A(G92gat), .ZN(new_n233));
  AOI22_X1  g032(.A1(KEYINPUT8), .A2(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  XOR2_X1   g034(.A(G99gat), .B(G106gat), .Z(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n228), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n227), .ZN(new_n239));
  INV_X1    g038(.A(new_n237), .ZN(new_n240));
  AOI22_X1  g039(.A1(new_n239), .A2(new_n240), .B1(KEYINPUT41), .B2(new_n202), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n209), .B1(new_n238), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n206), .B1(new_n242), .B2(KEYINPUT104), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(KEYINPUT105), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n238), .A2(new_n209), .A3(new_n241), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n244), .B1(new_n242), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G183gat), .B(G211gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(KEYINPUT101), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT99), .ZN(new_n250));
  XOR2_X1   g049(.A(G57gat), .B(G64gat), .Z(new_n251));
  NAND2_X1  g050(.A1(G71gat), .A2(G78gat), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT9), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT98), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT98), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n252), .A2(new_n256), .A3(new_n253), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n251), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n252), .ZN(new_n259));
  NOR2_X1   g058(.A1(G71gat), .A2(G78gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(KEYINPUT97), .B1(G71gat), .B2(G78gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n258), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n262), .B1(new_n258), .B2(new_n263), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n250), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n258), .A2(new_n263), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n261), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n269), .A2(KEYINPUT99), .A3(new_n264), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT21), .ZN(new_n273));
  NAND2_X1  g072(.A1(G231gat), .A2(G233gat), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  OAI211_X1 g074(.A(G231gat), .B(G233gat), .C1(new_n271), .C2(KEYINPUT21), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G127gat), .B(G155gat), .ZN(new_n278));
  XOR2_X1   g077(.A(new_n278), .B(KEYINPUT20), .Z(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n279), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n275), .A2(new_n281), .A3(new_n276), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n249), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n280), .A2(new_n249), .A3(new_n282), .ZN(new_n285));
  XNOR2_X1  g084(.A(G15gat), .B(G22gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT16), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n286), .B1(new_n287), .B2(G1gat), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n288), .B1(G1gat), .B2(new_n286), .ZN(new_n289));
  INV_X1    g088(.A(G8gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT90), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n291), .B1(new_n286), .B2(G1gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n289), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  OAI221_X1 g092(.A(new_n288), .B1(new_n291), .B2(G8gat), .C1(G1gat), .C2(new_n286), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(new_n272), .B2(new_n273), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n296), .B(new_n297), .Z(new_n298));
  NAND3_X1  g097(.A1(new_n284), .A2(new_n285), .A3(new_n298), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n243), .A2(KEYINPUT105), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n245), .A2(new_n242), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n243), .A2(KEYINPUT105), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n298), .ZN(new_n304));
  INV_X1    g103(.A(new_n285), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n304), .B1(new_n305), .B2(new_n283), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n246), .A2(new_n299), .A3(new_n303), .A4(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G230gat), .ZN(new_n308));
  INV_X1    g107(.A(G233gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT106), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n235), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n312), .B(new_n236), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(new_n266), .B2(new_n265), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT10), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n267), .A2(new_n270), .A3(new_n237), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n271), .A2(KEYINPUT10), .A3(new_n240), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n310), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n314), .A2(new_n316), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n310), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G120gat), .B(G148gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(G176gat), .B(G204gat), .ZN(new_n325));
  XOR2_X1   g124(.A(new_n324), .B(new_n325), .Z(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n320), .A2(new_n322), .A3(new_n326), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(KEYINPUT107), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT107), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n323), .A2(new_n331), .A3(new_n327), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  OR3_X1    g133(.A1(new_n307), .A2(KEYINPUT108), .A3(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT108), .B1(new_n307), .B2(new_n334), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT96), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n339));
  NAND2_X1  g138(.A1(KEYINPUT69), .A2(G183gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT27), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT27), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(KEYINPUT69), .A3(G183gat), .ZN(new_n343));
  INV_X1    g142(.A(G190gat), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT28), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT27), .B(G183gat), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(KEYINPUT28), .A3(new_n344), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G169gat), .A2(G176gat), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT26), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(G169gat), .A2(G176gat), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AND2_X1   g154(.A1(G183gat), .A2(G190gat), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n356), .B1(KEYINPUT26), .B2(new_n354), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n350), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT23), .B1(new_n354), .B2(KEYINPUT65), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT65), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT23), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n360), .B(new_n361), .C1(G169gat), .C2(G176gat), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n359), .A2(KEYINPUT25), .A3(new_n362), .A4(new_n351), .ZN(new_n363));
  NOR2_X1   g162(.A1(G183gat), .A2(G190gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(G183gat), .A2(G190gat), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT66), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n366), .A2(KEYINPUT24), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT24), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n368), .A2(KEYINPUT66), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n365), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT67), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n364), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n368), .A2(KEYINPUT66), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n366), .A2(KEYINPUT24), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n356), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT68), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g177(.A1(KEYINPUT68), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n375), .A2(KEYINPUT67), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n363), .B1(new_n372), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n359), .A2(new_n362), .A3(new_n351), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  OR2_X1    g182(.A1(new_n376), .A2(KEYINPUT64), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n365), .B1(new_n364), .B2(new_n368), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n376), .A2(KEYINPUT64), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT25), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n358), .B1(new_n381), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(G134gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n390), .A2(G127gat), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT70), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT1), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n394), .B1(G113gat), .B2(G120gat), .ZN(new_n395));
  AND2_X1   g194(.A1(G113gat), .A2(G120gat), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n393), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(G127gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n398), .A2(G134gat), .ZN(new_n399));
  NOR3_X1   g198(.A1(new_n399), .A2(new_n391), .A3(new_n392), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT72), .B1(new_n399), .B2(new_n391), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n390), .A2(G127gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n398), .A2(G134gat), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT72), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT73), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT71), .B(G120gat), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n395), .B1(new_n410), .B2(G113gat), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n409), .B1(new_n408), .B2(new_n411), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n402), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n339), .B1(new_n389), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n357), .B1(new_n354), .B2(new_n353), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n416), .B1(new_n347), .B2(new_n349), .ZN(new_n417));
  INV_X1    g216(.A(new_n363), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n378), .A2(new_n379), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n419), .B1(new_n370), .B2(new_n371), .ZN(new_n420));
  OAI22_X1  g219(.A1(new_n375), .A2(KEYINPUT67), .B1(G183gat), .B2(G190gat), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n418), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT25), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n423), .B1(new_n424), .B2(new_n382), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n417), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n407), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n406), .B1(new_n404), .B2(new_n405), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n411), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT73), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n401), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n426), .A2(new_n432), .A3(KEYINPUT74), .ZN(new_n433));
  NAND2_X1  g232(.A1(G227gat), .A2(G233gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n389), .A2(new_n414), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n415), .A2(new_n433), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(KEYINPUT34), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT32), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n415), .A2(new_n433), .A3(new_n435), .ZN(new_n439));
  INV_X1    g238(.A(new_n434), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(KEYINPUT75), .B(KEYINPUT33), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n442), .B1(new_n439), .B2(new_n440), .ZN(new_n443));
  XOR2_X1   g242(.A(G15gat), .B(G43gat), .Z(new_n444));
  XNOR2_X1  g243(.A(G71gat), .B(G99gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n441), .A2(new_n443), .A3(new_n447), .ZN(new_n448));
  AOI221_X4 g247(.A(new_n438), .B1(new_n442), .B2(new_n446), .C1(new_n439), .C2(new_n440), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n437), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n443), .A2(new_n447), .ZN(new_n451));
  INV_X1    g250(.A(new_n441), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n437), .ZN(new_n454));
  INV_X1    g253(.A(new_n449), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n450), .A2(new_n456), .A3(KEYINPUT77), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT36), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT77), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n459), .B(new_n437), .C1(new_n448), .C2(new_n449), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n457), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT76), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n450), .A2(new_n462), .ZN(new_n463));
  OAI211_X1 g262(.A(KEYINPUT76), .B(new_n437), .C1(new_n448), .C2(new_n449), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n463), .A2(KEYINPUT36), .A3(new_n464), .A4(new_n456), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT86), .ZN(new_n467));
  INV_X1    g266(.A(G155gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n205), .ZN(new_n469));
  NAND2_X1  g268(.A1(G155gat), .A2(G162gat), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(KEYINPUT2), .ZN(new_n472));
  XNOR2_X1  g271(.A(G141gat), .B(G148gat), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n472), .B1(new_n473), .B2(KEYINPUT79), .ZN(new_n474));
  INV_X1    g273(.A(G141gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(G148gat), .ZN(new_n476));
  INV_X1    g275(.A(G148gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(G141gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT79), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n471), .B1(new_n474), .B2(new_n481), .ZN(new_n482));
  OR2_X1    g281(.A1(new_n478), .A2(KEYINPUT80), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n478), .A2(KEYINPUT80), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n484), .A3(new_n476), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n470), .B1(new_n469), .B2(KEYINPUT2), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n414), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(G225gat), .A2(G233gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n479), .A2(new_n480), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n473), .A2(KEYINPUT79), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n492), .A3(new_n472), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n493), .A2(new_n471), .B1(new_n485), .B2(new_n486), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n494), .B(new_n402), .C1(new_n412), .C2(new_n413), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n489), .A2(new_n490), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT39), .ZN(new_n497));
  INV_X1    g296(.A(new_n490), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n432), .A2(KEYINPUT4), .A3(new_n494), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n488), .A2(KEYINPUT3), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT3), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n482), .A2(new_n487), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n414), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n500), .A2(new_n501), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n497), .B1(new_n498), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT39), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n508), .A3(new_n498), .ZN(new_n509));
  XOR2_X1   g308(.A(G1gat), .B(G29gat), .Z(new_n510));
  XNOR2_X1  g309(.A(G57gat), .B(G85gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT85), .ZN(new_n516));
  OAI22_X1  g315(.A1(new_n507), .A2(new_n515), .B1(new_n516), .B2(KEYINPUT40), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n506), .A2(new_n498), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n518), .A2(KEYINPUT39), .A3(new_n496), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n516), .A2(KEYINPUT40), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n519), .A2(new_n514), .A3(new_n520), .A4(new_n509), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n500), .A2(new_n501), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n523), .A2(KEYINPUT5), .A3(new_n490), .A4(new_n505), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n490), .B1(new_n489), .B2(new_n495), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT5), .ZN(new_n526));
  OAI22_X1  g325(.A1(new_n506), .A2(new_n498), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n514), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n524), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT78), .ZN(new_n530));
  NAND2_X1  g329(.A1(G226gat), .A2(G233gat), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT29), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n532), .B1(new_n389), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n426), .A2(new_n531), .ZN(new_n535));
  XNOR2_X1  g334(.A(G197gat), .B(G204gat), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT22), .ZN(new_n537));
  INV_X1    g336(.A(G211gat), .ZN(new_n538));
  INV_X1    g337(.A(G218gat), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  XOR2_X1   g340(.A(G211gat), .B(G218gat), .Z(new_n542));
  OR2_X1    g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n542), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NOR3_X1   g345(.A1(new_n534), .A2(new_n535), .A3(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n531), .B1(new_n426), .B2(KEYINPUT29), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n389), .A2(new_n532), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n545), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n530), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G8gat), .B(G36gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(G64gat), .B(G92gat), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n552), .B(new_n553), .Z(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n546), .B1(new_n534), .B2(new_n535), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n548), .A2(new_n545), .A3(new_n549), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT78), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n551), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n556), .A2(new_n557), .A3(new_n554), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT30), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT30), .A4(new_n554), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n529), .B1(new_n559), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n467), .B1(new_n522), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n551), .A2(KEYINPUT37), .A3(new_n558), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n547), .A2(new_n550), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT37), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n554), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT38), .ZN(new_n572));
  XOR2_X1   g371(.A(KEYINPUT82), .B(KEYINPUT6), .Z(new_n573));
  NAND2_X1  g372(.A1(new_n524), .A2(new_n527), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n573), .B1(new_n574), .B2(new_n514), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n529), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n524), .A2(new_n527), .A3(new_n528), .A4(new_n573), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n556), .A2(new_n557), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT38), .B1(new_n578), .B2(KEYINPUT37), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n570), .A2(new_n579), .B1(new_n554), .B2(new_n568), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n572), .A2(new_n576), .A3(new_n577), .A4(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT31), .B(G50gat), .ZN(new_n582));
  INV_X1    g381(.A(G228gat), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n583), .A2(new_n309), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n504), .A2(new_n533), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT84), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n504), .A2(KEYINPUT84), .A3(new_n533), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n588), .A2(new_n546), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT3), .B1(new_n545), .B2(new_n533), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n591), .A2(new_n494), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n585), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT29), .B1(new_n494), .B2(new_n503), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n595), .A2(new_n545), .ZN(new_n596));
  NOR3_X1   g395(.A1(new_n596), .A2(new_n592), .A3(new_n584), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n582), .B1(new_n594), .B2(new_n597), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n593), .B(new_n585), .C1(new_n545), .C2(new_n595), .ZN(new_n599));
  INV_X1    g398(.A(new_n582), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n545), .B1(new_n595), .B2(KEYINPUT84), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n592), .B1(new_n601), .B2(new_n588), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n599), .B(new_n600), .C1(new_n602), .C2(new_n585), .ZN(new_n603));
  XNOR2_X1  g402(.A(G78gat), .B(G106gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(G22gat), .ZN(new_n605));
  AND3_X1   g404(.A1(new_n598), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n605), .B1(new_n598), .B2(new_n603), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n517), .A2(new_n521), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n551), .A2(new_n555), .A3(new_n558), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n610), .A2(new_n562), .A3(new_n563), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n609), .A2(KEYINPUT86), .A3(new_n611), .A4(new_n529), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n566), .A2(new_n581), .A3(new_n608), .A4(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n607), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n598), .A2(new_n603), .A3(new_n605), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT83), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n529), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n524), .A2(new_n527), .A3(KEYINPUT83), .A4(new_n528), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n575), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n620), .A2(new_n577), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n616), .B1(new_n621), .B2(new_n611), .ZN(new_n622));
  AND3_X1   g421(.A1(new_n466), .A2(new_n613), .A3(new_n622), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n463), .A2(new_n464), .A3(new_n456), .A4(new_n608), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT87), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n621), .A2(new_n611), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n456), .A2(new_n615), .A3(new_n614), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT87), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n627), .A2(new_n628), .A3(new_n463), .A4(new_n464), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n625), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT35), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n576), .A2(new_n577), .ZN(new_n632));
  NOR4_X1   g431(.A1(new_n632), .A2(KEYINPUT35), .A3(new_n616), .A4(new_n611), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n457), .A2(new_n460), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n623), .B1(new_n631), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT91), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n293), .A2(new_n637), .A3(new_n294), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n637), .B1(new_n293), .B2(new_n294), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n221), .A2(KEYINPUT17), .A3(new_n225), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n641), .B1(new_n227), .B2(new_n210), .ZN(new_n642));
  OAI21_X1  g441(.A(KEYINPUT92), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n295), .A2(KEYINPUT91), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n293), .A2(new_n637), .A3(new_n294), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT92), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n646), .A2(new_n228), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G229gat), .A2(G233gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT93), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n227), .A2(new_n295), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n643), .A2(new_n648), .A3(new_n651), .A4(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT18), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n227), .B(new_n295), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT94), .B(KEYINPUT13), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n650), .B(new_n657), .ZN(new_n658));
  AOI22_X1  g457(.A1(new_n654), .A2(new_n655), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n640), .A2(new_n642), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n652), .B1(new_n660), .B2(new_n647), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n661), .A2(KEYINPUT18), .A3(new_n651), .A4(new_n643), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G113gat), .B(G141gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(G197gat), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT11), .B(G169gat), .Z(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT12), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT95), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n655), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n658), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n662), .A2(new_n672), .A3(new_n668), .A4(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n670), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  AOI211_X1 g474(.A(new_n671), .B(new_n668), .C1(new_n659), .C2(new_n662), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n338), .B1(new_n636), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n674), .A2(new_n671), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n668), .B1(new_n659), .B2(new_n662), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(new_n676), .ZN(new_n683));
  AOI22_X1  g482(.A1(new_n630), .A2(KEYINPUT35), .B1(new_n634), .B2(new_n633), .ZN(new_n684));
  OAI211_X1 g483(.A(KEYINPUT96), .B(new_n683), .C1(new_n684), .C2(new_n623), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n337), .B1(new_n679), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n621), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G1gat), .ZN(G1324gat));
  INV_X1    g487(.A(new_n686), .ZN(new_n689));
  INV_X1    g488(.A(new_n611), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT16), .B(G8gat), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n290), .B1(new_n686), .B2(new_n611), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT42), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(KEYINPUT42), .B2(new_n692), .ZN(G1325gat));
  INV_X1    g494(.A(new_n634), .ZN(new_n696));
  OR3_X1    g495(.A1(new_n689), .A2(G15gat), .A3(new_n696), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n466), .A2(KEYINPUT109), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n466), .A2(KEYINPUT109), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G15gat), .B1(new_n689), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n697), .A2(new_n701), .ZN(G1326gat));
  NAND2_X1  g501(.A1(new_n679), .A2(new_n685), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n703), .A2(new_n616), .A3(new_n336), .A4(new_n335), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT43), .B(G22gat), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1327gat));
  NAND2_X1  g505(.A1(new_n246), .A2(new_n303), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n306), .A2(new_n299), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n333), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n712), .B1(new_n679), .B2(new_n685), .ZN(new_n713));
  INV_X1    g512(.A(G29gat), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n713), .A2(new_n714), .A3(new_n621), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT45), .ZN(new_n716));
  OAI21_X1  g515(.A(KEYINPUT44), .B1(new_n636), .B2(new_n708), .ZN(new_n717));
  XNOR2_X1  g516(.A(KEYINPUT112), .B(KEYINPUT44), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n707), .B(new_n718), .C1(new_n684), .C2(new_n623), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(new_n682), .B2(new_n676), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n675), .A2(new_n677), .A3(KEYINPUT110), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n333), .B(KEYINPUT111), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n725), .A2(new_n709), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n720), .A2(new_n621), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n714), .B1(new_n730), .B2(KEYINPUT113), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(KEYINPUT113), .B2(new_n730), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n732), .ZN(G1328gat));
  INV_X1    g532(.A(G36gat), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n713), .A2(new_n734), .A3(new_n611), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT46), .Z(new_n736));
  NAND3_X1  g535(.A1(new_n720), .A2(new_n611), .A3(new_n729), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n734), .B1(new_n737), .B2(KEYINPUT114), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(KEYINPUT114), .B2(new_n737), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n736), .A2(new_n739), .ZN(G1329gat));
  NOR2_X1   g539(.A1(new_n696), .A2(G43gat), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n713), .A2(new_n741), .ZN(new_n742));
  AOI211_X1 g541(.A(new_n466), .B(new_n728), .C1(new_n717), .C2(new_n719), .ZN(new_n743));
  INV_X1    g542(.A(G43gat), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n742), .B(KEYINPUT47), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n720), .A2(new_n699), .A3(new_n698), .A4(new_n729), .ZN(new_n746));
  AOI22_X1  g545(.A1(new_n746), .A2(G43gat), .B1(new_n713), .B2(new_n741), .ZN(new_n747));
  XOR2_X1   g546(.A(KEYINPUT115), .B(KEYINPUT47), .Z(new_n748));
  OAI21_X1  g547(.A(new_n745), .B1(new_n747), .B2(new_n748), .ZN(G1330gat));
  NOR2_X1   g548(.A1(new_n712), .A2(G50gat), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n703), .A2(new_n616), .A3(new_n750), .ZN(new_n751));
  AOI211_X1 g550(.A(new_n608), .B(new_n728), .C1(new_n717), .C2(new_n719), .ZN(new_n752));
  INV_X1    g551(.A(G50gat), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT116), .B1(new_n752), .B2(new_n753), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n754), .A2(new_n755), .A3(KEYINPUT48), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT48), .ZN(new_n757));
  OAI221_X1 g556(.A(new_n751), .B1(KEYINPUT116), .B2(new_n757), .C1(new_n752), .C2(new_n753), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n756), .A2(new_n758), .ZN(G1331gat));
  INV_X1    g558(.A(new_n636), .ZN(new_n760));
  INV_X1    g559(.A(new_n307), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n760), .A2(new_n761), .A3(new_n724), .A4(new_n726), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n620), .A2(new_n577), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XOR2_X1   g563(.A(KEYINPUT117), .B(G57gat), .Z(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(G1332gat));
  AOI211_X1 g565(.A(new_n690), .B(new_n762), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n767));
  NOR2_X1   g566(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n767), .B(new_n768), .ZN(G1333gat));
  OAI21_X1  g568(.A(G71gat), .B1(new_n762), .B2(new_n700), .ZN(new_n770));
  OR2_X1    g569(.A1(new_n696), .A2(G71gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n762), .B2(new_n771), .ZN(new_n772));
  XOR2_X1   g571(.A(new_n772), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g572(.A1(new_n762), .A2(new_n608), .ZN(new_n774));
  XOR2_X1   g573(.A(new_n774), .B(G78gat), .Z(G1335gat));
  NAND3_X1  g574(.A1(new_n724), .A2(new_n709), .A3(new_n334), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n776), .B1(new_n717), .B2(new_n719), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(G85gat), .B1(new_n778), .B2(new_n763), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n760), .A2(KEYINPUT51), .A3(new_n724), .A4(new_n711), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n724), .B(new_n711), .C1(new_n684), .C2(new_n623), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n334), .A2(new_n232), .A3(new_n621), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n779), .B1(new_n785), .B2(new_n786), .ZN(G1336gat));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n788));
  AOI211_X1 g587(.A(new_n690), .B(new_n776), .C1(new_n717), .C2(new_n719), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n726), .A2(new_n233), .A3(new_n611), .ZN(new_n790));
  OAI221_X1 g589(.A(new_n788), .B1(new_n789), .B2(new_n233), .C1(new_n785), .C2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n776), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n720), .A2(new_n611), .A3(new_n792), .ZN(new_n793));
  XOR2_X1   g592(.A(new_n790), .B(KEYINPUT118), .Z(new_n794));
  AOI22_X1  g593(.A1(new_n793), .A2(G92gat), .B1(new_n784), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT119), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n795), .A2(new_n796), .A3(new_n788), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n781), .A2(new_n782), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n794), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n800), .B1(new_n789), .B2(new_n233), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT119), .B1(new_n801), .B2(KEYINPUT52), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n791), .B1(new_n797), .B2(new_n802), .ZN(G1337gat));
  OAI21_X1  g602(.A(G99gat), .B1(new_n778), .B2(new_n700), .ZN(new_n804));
  OR3_X1    g603(.A1(new_n696), .A2(G99gat), .A3(new_n333), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n785), .B2(new_n805), .ZN(G1338gat));
  INV_X1    g605(.A(G106gat), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n616), .A2(new_n807), .ZN(new_n808));
  AOI211_X1 g607(.A(new_n727), .B(new_n808), .C1(new_n780), .C2(new_n783), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n807), .B1(new_n777), .B2(new_n616), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g610(.A(KEYINPUT120), .B(KEYINPUT53), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n811), .B(new_n812), .ZN(G1339gat));
  NAND3_X1  g612(.A1(new_n317), .A2(new_n310), .A3(new_n318), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n320), .A2(KEYINPUT54), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n326), .B1(new_n319), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(KEYINPUT55), .A3(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n818), .A2(new_n329), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n815), .A2(new_n817), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n722), .A2(new_n723), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n651), .B1(new_n661), .B2(new_n643), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n656), .A2(new_n658), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n667), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n827), .A2(new_n674), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n334), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n707), .B1(new_n824), .B2(new_n829), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n823), .A2(new_n707), .A3(new_n828), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n709), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n724), .A2(new_n761), .A3(new_n333), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n616), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n763), .A2(new_n611), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n634), .A3(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(G113gat), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n836), .A2(new_n837), .A3(new_n678), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n763), .B1(new_n832), .B2(new_n833), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n625), .A2(new_n629), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(new_n690), .A3(new_n725), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n838), .B1(new_n843), .B2(new_n837), .ZN(G1340gat));
  OAI21_X1  g643(.A(G120gat), .B1(new_n836), .B2(new_n727), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n842), .A2(new_n690), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n333), .A2(new_n410), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(G1341gat));
  OAI21_X1  g647(.A(G127gat), .B1(new_n836), .B2(new_n709), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n710), .A2(new_n398), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n849), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT121), .ZN(G1342gat));
  NOR2_X1   g651(.A1(new_n708), .A2(new_n611), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n842), .A2(new_n390), .A3(new_n853), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n854), .A2(KEYINPUT56), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(KEYINPUT56), .ZN(new_n856));
  OAI21_X1  g655(.A(G134gat), .B1(new_n836), .B2(new_n708), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(G1343gat));
  AOI21_X1  g657(.A(new_n608), .B1(new_n832), .B2(new_n833), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n466), .A2(new_n835), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n675), .A2(new_n677), .A3(new_n822), .A4(new_n819), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n707), .B1(new_n863), .B2(new_n829), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n709), .B1(new_n864), .B2(new_n831), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n833), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n616), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n862), .B1(new_n867), .B2(KEYINPUT57), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n861), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n725), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n608), .B1(new_n698), .B2(new_n699), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n839), .A2(new_n871), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n872), .A2(new_n690), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n678), .A2(G141gat), .ZN(new_n874));
  AOI22_X1  g673(.A1(new_n870), .A2(G141gat), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT58), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n475), .B1(new_n869), .B2(new_n683), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n872), .A2(new_n690), .A3(new_n874), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n876), .ZN(new_n879));
  OAI22_X1  g678(.A1(new_n875), .A2(new_n876), .B1(new_n877), .B2(new_n879), .ZN(G1344gat));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n865), .B1(new_n337), .B2(new_n683), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n860), .A3(new_n616), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n862), .A2(new_n333), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n883), .B(new_n884), .C1(new_n859), .C2(new_n860), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(G148gat), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n861), .A2(new_n868), .A3(new_n334), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n477), .A2(KEYINPUT59), .ZN(new_n888));
  AOI22_X1  g687(.A1(new_n886), .A2(KEYINPUT59), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n333), .A2(G148gat), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n872), .A2(new_n690), .A3(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n881), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n887), .A2(new_n888), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n895), .B1(new_n885), .B2(G148gat), .ZN(new_n896));
  OAI211_X1 g695(.A(KEYINPUT122), .B(new_n891), .C1(new_n894), .C2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n893), .A2(new_n897), .ZN(G1345gat));
  INV_X1    g697(.A(new_n869), .ZN(new_n899));
  OAI21_X1  g698(.A(G155gat), .B1(new_n899), .B2(new_n709), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n873), .A2(new_n468), .A3(new_n710), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(G1346gat));
  OAI21_X1  g701(.A(G162gat), .B1(new_n899), .B2(new_n708), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n872), .A2(new_n205), .A3(new_n853), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1347gat));
  AOI21_X1  g704(.A(new_n621), .B1(new_n832), .B2(new_n833), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n840), .A2(new_n611), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(G169gat), .B1(new_n909), .B2(new_n725), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n763), .A2(new_n611), .ZN(new_n911));
  XOR2_X1   g710(.A(new_n911), .B(KEYINPUT123), .Z(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n634), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n913), .B(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n834), .ZN(new_n916));
  INV_X1    g715(.A(G169gat), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n916), .A2(new_n917), .A3(new_n678), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n910), .A2(new_n918), .ZN(G1348gat));
  OAI21_X1  g718(.A(G176gat), .B1(new_n916), .B2(new_n727), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n333), .A2(G176gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n908), .B2(new_n921), .ZN(G1349gat));
  OAI21_X1  g721(.A(G183gat), .B1(new_n916), .B2(new_n709), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n710), .A2(new_n348), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n908), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g725(.A1(new_n909), .A2(new_n344), .A3(new_n707), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n915), .A2(new_n834), .A3(new_n707), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(G190gat), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(KEYINPUT125), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT61), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n928), .A2(new_n932), .A3(G190gat), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n931), .B1(new_n930), .B2(new_n933), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n927), .B1(new_n934), .B2(new_n935), .ZN(G1351gat));
  AND2_X1   g735(.A1(new_n700), .A2(new_n912), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n883), .B(new_n937), .C1(new_n859), .C2(new_n860), .ZN(new_n938));
  INV_X1    g737(.A(G197gat), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n938), .A2(new_n939), .A3(new_n678), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n871), .A2(new_n611), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n906), .A2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n944), .A2(KEYINPUT126), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(KEYINPUT126), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n945), .A2(new_n725), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n940), .B1(new_n947), .B2(new_n939), .ZN(G1352gat));
  NOR3_X1   g747(.A1(new_n943), .A2(G204gat), .A3(new_n333), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT62), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n950), .ZN(new_n952));
  OAI21_X1  g751(.A(G204gat), .B1(new_n938), .B2(new_n727), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(G1353gat));
  OR2_X1    g753(.A1(new_n938), .A2(new_n709), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT63), .B1(new_n955), .B2(G211gat), .ZN(new_n956));
  OAI211_X1 g755(.A(KEYINPUT63), .B(G211gat), .C1(new_n938), .C2(new_n709), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n945), .A2(new_n946), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n710), .A2(new_n538), .ZN(new_n960));
  OAI22_X1  g759(.A1(new_n956), .A2(new_n958), .B1(new_n959), .B2(new_n960), .ZN(G1354gat));
  OAI21_X1  g760(.A(G218gat), .B1(new_n938), .B2(new_n708), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n707), .A2(new_n539), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n959), .B2(new_n963), .ZN(G1355gat));
endmodule


