//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 0 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(KEYINPUT23), .A3(G119), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT73), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G128), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT74), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  OAI22_X1  g010(.A1(new_n193), .A2(new_n194), .B1(new_n192), .B2(G128), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n190), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(G119), .B(G128), .ZN(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT24), .B(G110), .ZN(new_n200));
  XNOR2_X1  g014(.A(new_n200), .B(KEYINPUT72), .ZN(new_n201));
  OAI22_X1  g015(.A1(new_n198), .A2(G110), .B1(new_n199), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G125), .ZN(new_n204));
  NOR3_X1   g018(.A1(new_n204), .A2(KEYINPUT75), .A3(KEYINPUT16), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(G125), .B(G140), .ZN(new_n207));
  AOI21_X1  g021(.A(KEYINPUT75), .B1(new_n207), .B2(KEYINPUT16), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n204), .A2(KEYINPUT16), .ZN(new_n209));
  OAI211_X1 g023(.A(G146), .B(new_n206), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G125), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G140), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT64), .A2(G146), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n213), .A2(new_n204), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n202), .A2(new_n210), .A3(new_n217), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n198), .A2(G110), .B1(new_n201), .B2(new_n199), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n204), .A2(new_n215), .A3(KEYINPUT16), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT75), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n209), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n212), .B1(new_n222), .B2(new_n205), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n210), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n218), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT22), .B(G137), .ZN(new_n227));
  INV_X1    g041(.A(G953), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(G221), .A3(G234), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n227), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n230), .B(KEYINPUT76), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G902), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n218), .A2(new_n225), .A3(new_n230), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT25), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n232), .A2(KEYINPUT25), .A3(new_n233), .A4(new_n234), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  XOR2_X1   g053(.A(KEYINPUT71), .B(G217), .Z(new_n240));
  AOI21_X1  g054(.A(new_n240), .B1(G234), .B2(new_n233), .ZN(new_n241));
  AOI21_X1  g055(.A(KEYINPUT77), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT77), .ZN(new_n243));
  INV_X1    g057(.A(new_n241), .ZN(new_n244));
  AOI211_X1 g058(.A(new_n243), .B(new_n244), .C1(new_n237), .C2(new_n238), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n232), .A2(new_n234), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n241), .A2(G902), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(G237), .A2(G953), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G210), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n253), .B(KEYINPUT68), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT26), .B(G101), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n257));
  XOR2_X1   g071(.A(new_n256), .B(new_n257), .Z(new_n258));
  NAND2_X1  g072(.A1(new_n192), .A2(G116), .ZN(new_n259));
  INV_X1    g073(.A(G116), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G119), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT2), .B(G113), .ZN(new_n263));
  OR2_X1    g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n263), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n213), .A2(G143), .A3(new_n216), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n212), .A2(G143), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n187), .A2(KEYINPUT1), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n187), .B1(new_n267), .B2(KEYINPUT1), .ZN(new_n272));
  INV_X1    g086(.A(G143), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(G146), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n213), .A2(new_n216), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n274), .B1(new_n275), .B2(new_n273), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n271), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT66), .ZN(new_n278));
  INV_X1    g092(.A(G137), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n278), .B1(new_n279), .B2(G134), .ZN(new_n280));
  INV_X1    g094(.A(G134), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(KEYINPUT66), .A3(G137), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n280), .A2(new_n282), .B1(G134), .B2(new_n279), .ZN(new_n283));
  INV_X1    g097(.A(G131), .ZN(new_n284));
  OR2_X1    g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT11), .B1(new_n281), .B2(G137), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT11), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(new_n279), .A3(G134), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n286), .A2(new_n288), .B1(new_n281), .B2(G137), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n284), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n277), .A2(new_n285), .A3(new_n290), .ZN(new_n291));
  AND2_X1   g105(.A1(KEYINPUT64), .A2(G146), .ZN(new_n292));
  NOR2_X1   g106(.A1(KEYINPUT64), .A2(G146), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n268), .B1(new_n294), .B2(G143), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(KEYINPUT0), .A3(G128), .ZN(new_n296));
  INV_X1    g110(.A(new_n274), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n297), .B1(new_n294), .B2(G143), .ZN(new_n298));
  XOR2_X1   g112(.A(KEYINPUT0), .B(G128), .Z(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n284), .A2(KEYINPUT65), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n289), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n289), .A2(new_n302), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n296), .B(new_n300), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT30), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n291), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n306), .B1(new_n291), .B2(new_n305), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n266), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n266), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n291), .A2(new_n305), .A3(new_n310), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n258), .A2(new_n309), .A3(KEYINPUT31), .A4(new_n311), .ZN(new_n312));
  AND2_X1   g126(.A1(new_n312), .A2(new_n233), .ZN(new_n313));
  INV_X1    g127(.A(G472), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n256), .B(new_n257), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT28), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n291), .A2(new_n305), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n266), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n316), .B1(new_n318), .B2(new_n311), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n311), .A2(new_n316), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n315), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n258), .A2(new_n309), .A3(new_n311), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT31), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  AND3_X1   g139(.A1(new_n313), .A2(new_n314), .A3(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n308), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n291), .A2(new_n305), .A3(new_n306), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n310), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n311), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n315), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT29), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n310), .B1(new_n291), .B2(new_n305), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT28), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(new_n258), .A3(new_n320), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n331), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n334), .A2(new_n258), .A3(KEYINPUT29), .A4(new_n320), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n233), .A3(new_n337), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n326), .A2(KEYINPUT32), .B1(new_n338), .B2(G472), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n313), .A2(new_n325), .A3(new_n314), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT32), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT69), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT69), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n340), .A2(new_n344), .A3(new_n341), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n339), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT70), .ZN(new_n347));
  AND3_X1   g161(.A1(new_n340), .A2(new_n344), .A3(new_n341), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n344), .B1(new_n340), .B2(new_n341), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT70), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n351), .A3(new_n339), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n251), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(G214), .B1(G237), .B2(G902), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n296), .A2(new_n300), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G125), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n356), .B1(G125), .B2(new_n277), .ZN(new_n357));
  INV_X1    g171(.A(G224), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n358), .A2(G953), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n359), .B(KEYINPUT85), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n357), .B(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G101), .ZN(new_n363));
  INV_X1    g177(.A(G107), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G104), .ZN(new_n365));
  INV_X1    g179(.A(G104), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G107), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n363), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT3), .B1(new_n366), .B2(G107), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT3), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(new_n364), .A3(G104), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n370), .A2(new_n372), .A3(new_n363), .A4(new_n367), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT78), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n373), .A2(new_n374), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n369), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT81), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n372), .A2(new_n367), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n379), .A2(KEYINPUT78), .A3(new_n363), .A4(new_n370), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n373), .A2(new_n374), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n368), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT81), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n259), .A2(new_n261), .A3(KEYINPUT5), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n385), .B(G113), .C1(KEYINPUT5), .C2(new_n259), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n386), .A2(new_n264), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n378), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n370), .A2(new_n372), .A3(new_n367), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT4), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n389), .A2(new_n390), .A3(G101), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n380), .A2(new_n381), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n390), .B1(new_n389), .B2(G101), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n266), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n388), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(G110), .B(G122), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT83), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n396), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n401), .B1(new_n396), .B2(new_n398), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT84), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n406), .B1(new_n396), .B2(new_n398), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n388), .A2(KEYINPUT84), .A3(new_n395), .A4(new_n397), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(KEYINPUT6), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n362), .B1(new_n405), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT7), .B1(new_n358), .B2(G953), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n357), .B(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n377), .B(new_n387), .ZN(new_n413));
  XOR2_X1   g227(.A(new_n397), .B(KEYINPUT8), .Z(new_n414));
  NOR2_X1   g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n407), .A2(new_n408), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n233), .ZN(new_n419));
  OAI21_X1  g233(.A(G210), .B1(G237), .B2(G902), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NOR3_X1   g235(.A1(new_n410), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n407), .A2(KEYINPUT6), .A3(new_n408), .ZN(new_n423));
  INV_X1    g237(.A(new_n404), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n402), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n361), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(G902), .B1(new_n416), .B2(new_n417), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n420), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n354), .B1(new_n422), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G469), .ZN(new_n430));
  XNOR2_X1  g244(.A(G110), .B(G140), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n228), .A2(G227), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n431), .B(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n277), .A2(KEYINPUT10), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n378), .A2(new_n384), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n394), .A2(new_n296), .A3(new_n300), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT80), .ZN(new_n438));
  XOR2_X1   g252(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n439));
  AOI21_X1  g253(.A(new_n187), .B1(new_n297), .B2(KEYINPUT1), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n271), .B1(new_n295), .B2(new_n440), .ZN(new_n441));
  AOI211_X1 g255(.A(new_n438), .B(new_n439), .C1(new_n382), .C2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n392), .A2(new_n369), .A3(new_n441), .ZN(new_n443));
  INV_X1    g257(.A(new_n439), .ZN(new_n444));
  AOI21_X1  g258(.A(KEYINPUT80), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n436), .B(new_n437), .C1(new_n442), .C2(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n303), .A2(new_n304), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(KEYINPUT82), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n434), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n443), .B1(new_n277), .B2(new_n382), .ZN(new_n451));
  INV_X1    g265(.A(new_n447), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(KEYINPUT12), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n452), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT12), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n450), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n436), .A2(new_n437), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n443), .A2(new_n444), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n438), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n443), .A2(KEYINPUT80), .A3(new_n444), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n458), .A2(new_n462), .A3(new_n448), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n446), .A2(new_n452), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n434), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n430), .B(new_n233), .C1(new_n457), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(G469), .A2(G902), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n451), .A2(KEYINPUT12), .A3(new_n452), .ZN(new_n468));
  AOI21_X1  g282(.A(KEYINPUT12), .B1(new_n451), .B2(new_n452), .ZN(new_n469));
  OAI22_X1  g283(.A1(new_n446), .A2(new_n449), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n433), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n463), .A2(new_n464), .A3(new_n434), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(new_n472), .A3(G469), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n466), .A2(new_n467), .A3(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT9), .B(G234), .ZN(new_n475));
  OAI21_X1  g289(.A(G221), .B1(new_n475), .B2(G902), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT87), .ZN(new_n478));
  INV_X1    g292(.A(G237), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(new_n228), .A3(G214), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n273), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n252), .A2(G143), .A3(G214), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n478), .B1(new_n483), .B2(G131), .ZN(new_n484));
  AOI211_X1 g298(.A(KEYINPUT87), .B(new_n284), .C1(new_n481), .C2(new_n482), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT17), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT89), .ZN(new_n487));
  INV_X1    g301(.A(new_n224), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT89), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n489), .B(KEYINPUT17), .C1(new_n484), .C2(new_n485), .ZN(new_n490));
  AND4_X1   g304(.A1(G143), .A2(new_n479), .A3(new_n228), .A4(G214), .ZN(new_n491));
  AOI21_X1  g305(.A(G143), .B1(new_n252), .B2(G214), .ZN(new_n492));
  OAI21_X1  g306(.A(G131), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT87), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n483), .A2(new_n478), .A3(G131), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT17), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n481), .A2(new_n284), .A3(new_n482), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n494), .A2(new_n495), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n487), .A2(new_n488), .A3(new_n490), .A4(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n214), .A2(G140), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n203), .A2(G125), .ZN(new_n501));
  OAI21_X1  g315(.A(G146), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n217), .ZN(new_n503));
  NAND2_X1  g317(.A1(KEYINPUT18), .A2(G131), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n505), .B1(new_n491), .B2(new_n492), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n481), .A2(new_n482), .A3(new_n504), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n503), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT86), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT86), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n503), .A2(new_n506), .A3(new_n510), .A4(new_n507), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n499), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(G113), .B(G122), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(new_n366), .ZN(new_n515));
  OR2_X1    g329(.A1(new_n515), .A2(KEYINPUT90), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n233), .B1(new_n513), .B2(new_n516), .ZN(new_n518));
  OAI21_X1  g332(.A(G475), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(G475), .A2(G902), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT88), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n207), .A2(KEYINPUT19), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT19), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n524), .B1(new_n500), .B2(new_n501), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n275), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n222), .A2(new_n205), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n526), .B1(new_n527), .B2(G146), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n528), .A2(new_n529), .B1(new_n509), .B2(new_n511), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n522), .B1(new_n530), .B2(new_n515), .ZN(new_n531));
  INV_X1    g345(.A(new_n526), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n529), .A2(new_n210), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n512), .ZN(new_n534));
  INV_X1    g348(.A(new_n515), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(KEYINPUT88), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n499), .A2(new_n515), .A3(new_n512), .ZN(new_n538));
  AOI211_X1 g352(.A(KEYINPUT20), .B(new_n521), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT20), .ZN(new_n540));
  AOI21_X1  g354(.A(KEYINPUT88), .B1(new_n534), .B2(new_n535), .ZN(new_n541));
  AOI211_X1 g355(.A(new_n522), .B(new_n515), .C1(new_n533), .C2(new_n512), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n538), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n540), .B1(new_n543), .B2(new_n520), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n519), .B1(new_n539), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT91), .ZN(new_n546));
  NAND2_X1  g360(.A1(G234), .A2(G237), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n547), .A2(G952), .A3(new_n228), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n547), .A2(G902), .A3(G953), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT21), .B(G898), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT91), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n553), .B(new_n519), .C1(new_n539), .C2(new_n544), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT93), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n260), .A2(G122), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n260), .A2(G122), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n555), .B(new_n556), .C1(new_n557), .C2(KEYINPUT14), .ZN(new_n558));
  INV_X1    g372(.A(G122), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(G116), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT14), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(G116), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(KEYINPUT93), .B1(new_n556), .B2(KEYINPUT14), .ZN(new_n564));
  OAI211_X1 g378(.A(G107), .B(new_n558), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n562), .A2(new_n556), .A3(new_n364), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT92), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(new_n273), .B2(G128), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n187), .A2(KEYINPUT92), .A3(G143), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n273), .A2(G128), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n281), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n281), .B1(new_n570), .B2(new_n571), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n565), .B(new_n566), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT13), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n273), .A2(KEYINPUT13), .A3(G128), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n570), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(G107), .B1(new_n557), .B2(new_n560), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n579), .A2(G134), .B1(new_n580), .B2(new_n566), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n572), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n575), .A2(new_n582), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n240), .A2(G953), .A3(new_n475), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT94), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n575), .A2(new_n582), .A3(new_n584), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n583), .A2(KEYINPUT94), .A3(new_n585), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(new_n233), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(G478), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(KEYINPUT15), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n591), .A2(new_n593), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n546), .A2(new_n552), .A3(new_n554), .A4(new_n597), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n429), .A2(new_n477), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n353), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(G101), .ZN(G3));
  NAND2_X1  g415(.A1(new_n313), .A2(new_n325), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G472), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n246), .A2(new_n340), .A3(new_n250), .A4(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n604), .A2(new_n477), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(KEYINPUT95), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n354), .B(new_n552), .C1(new_n422), .C2(new_n428), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n546), .A2(new_n554), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n592), .A2(G902), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n610));
  INV_X1    g424(.A(new_n588), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n584), .B1(new_n575), .B2(new_n582), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n611), .B1(KEYINPUT96), .B2(new_n612), .ZN(new_n613));
  OR2_X1    g427(.A1(new_n612), .A2(KEYINPUT96), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n610), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(KEYINPUT33), .B1(new_n589), .B2(new_n590), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n609), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n591), .A2(new_n592), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n608), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n607), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n606), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT34), .B(G104), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  INV_X1    g438(.A(KEYINPUT98), .ZN(new_n625));
  INV_X1    g439(.A(new_n512), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n496), .B1(new_n494), .B2(new_n495), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT89), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n488), .A2(new_n498), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n626), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n630), .A2(new_n515), .B1(new_n531), .B2(new_n536), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT20), .B1(new_n631), .B2(new_n521), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT97), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n543), .A2(new_n540), .A3(new_n520), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n539), .A2(KEYINPUT97), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n596), .A2(new_n519), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n625), .B1(new_n607), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n354), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n421), .B1(new_n410), .B2(new_n419), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n426), .A2(new_n420), .A3(new_n427), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n638), .A2(new_n636), .A3(new_n635), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n644), .A2(new_n645), .A3(KEYINPUT98), .A4(new_n552), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n606), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT99), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT35), .B(G107), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G9));
  NAND2_X1  g465(.A1(new_n239), .A2(new_n241), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n243), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n226), .B(KEYINPUT100), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n231), .A2(KEYINPUT36), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n654), .A2(KEYINPUT36), .A3(new_n231), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n249), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n239), .A2(KEYINPUT77), .A3(new_n241), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n653), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(new_n474), .A3(new_n476), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n603), .A2(new_n340), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n598), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n664), .A2(new_n644), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT37), .B(G110), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  INV_X1    g482(.A(G900), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n548), .B1(new_n549), .B2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n639), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n662), .A2(new_n429), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n351), .B1(new_n350), .B2(new_n339), .ZN(new_n673));
  AND4_X1   g487(.A1(new_n351), .A2(new_n339), .A3(new_n343), .A4(new_n345), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n671), .B(new_n672), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G128), .ZN(G30));
  INV_X1    g490(.A(KEYINPUT40), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n670), .B(KEYINPUT39), .Z(new_n678));
  NAND4_X1  g492(.A1(new_n474), .A2(new_n677), .A3(new_n476), .A4(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n642), .A2(new_n643), .A3(KEYINPUT38), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT38), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n681), .B1(new_n422), .B2(new_n428), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n679), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n661), .A2(new_n641), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n313), .A2(new_n325), .A3(KEYINPUT32), .A4(new_n314), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n315), .B1(new_n330), .B2(new_n333), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n323), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g501(.A(G472), .B1(new_n687), .B2(G902), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n343), .A2(new_n689), .A3(new_n345), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n597), .B1(new_n546), .B2(new_n554), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n684), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n678), .ZN(new_n693));
  OAI21_X1  g507(.A(KEYINPUT40), .B1(new_n477), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n683), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G143), .ZN(G45));
  NAND2_X1  g510(.A1(new_n347), .A2(new_n352), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT101), .ZN(new_n698));
  INV_X1    g512(.A(new_n670), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n608), .A2(new_n698), .A3(new_n619), .A4(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n608), .A2(new_n619), .A3(new_n699), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT101), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n697), .A2(new_n672), .A3(new_n700), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  OAI21_X1  g518(.A(new_n233), .B1(new_n457), .B2(new_n465), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(G469), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n476), .A3(new_n466), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n353), .A2(new_n621), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT41), .B(G113), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G15));
  NAND3_X1  g525(.A1(new_n353), .A2(new_n647), .A3(new_n708), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G116), .ZN(G18));
  INV_X1    g527(.A(new_n661), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n429), .A2(new_n714), .A3(new_n707), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n697), .A2(new_n665), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  XNOR2_X1  g531(.A(new_n691), .B(KEYINPUT103), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n429), .A2(new_n707), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n720), .B1(new_n603), .B2(new_n340), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT102), .B1(new_n602), .B2(G472), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n251), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n718), .A2(new_n552), .A3(new_n719), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G122), .ZN(G24));
  NOR2_X1   g539(.A1(new_n721), .A2(new_n722), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n715), .A2(new_n702), .A3(new_n700), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G125), .ZN(G27));
  INV_X1    g542(.A(KEYINPUT42), .ZN(new_n729));
  INV_X1    g543(.A(new_n251), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n642), .A2(new_n643), .A3(new_n354), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n477), .A2(new_n731), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n730), .B(new_n732), .C1(new_n673), .C2(new_n674), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n702), .A2(new_n700), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n729), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n734), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT104), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n339), .A2(new_n342), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n730), .A2(KEYINPUT42), .A3(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n736), .A2(new_n737), .A3(new_n732), .A4(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n739), .A2(new_n700), .A3(new_n702), .A4(new_n732), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT104), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n735), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(KEYINPUT105), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT105), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n735), .A2(new_n740), .A3(new_n745), .A4(new_n742), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n284), .ZN(G33));
  INV_X1    g562(.A(new_n671), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n733), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(new_n281), .ZN(G36));
  INV_X1    g565(.A(KEYINPUT106), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT45), .B1(new_n471), .B2(new_n472), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n752), .B1(new_n753), .B2(new_n430), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n447), .B1(new_n458), .B2(new_n462), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n450), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n456), .A2(new_n453), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n434), .B1(new_n463), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n755), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(KEYINPUT106), .A3(G469), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT45), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n754), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(KEYINPUT46), .A3(new_n467), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT46), .B1(new_n763), .B2(new_n467), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT107), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n466), .B(new_n764), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  AOI211_X1 g581(.A(KEYINPUT107), .B(KEYINPUT46), .C1(new_n763), .C2(new_n467), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n476), .B(new_n678), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n661), .A2(new_n663), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT109), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n632), .A2(new_n634), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n553), .B1(new_n774), .B2(new_n519), .ZN(new_n775));
  INV_X1    g589(.A(new_n554), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n773), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n546), .A2(KEYINPUT109), .A3(new_n554), .ZN(new_n778));
  INV_X1    g592(.A(new_n619), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT43), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n777), .A2(new_n778), .A3(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT108), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n619), .A2(KEYINPUT108), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n784), .A2(new_n546), .A3(new_n554), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n780), .ZN(new_n787));
  AOI211_X1 g601(.A(new_n771), .B(new_n772), .C1(new_n782), .C2(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT110), .B1(new_n788), .B2(new_n731), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT110), .ZN(new_n790));
  INV_X1    g604(.A(new_n731), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n782), .A2(new_n787), .ZN(new_n792));
  INV_X1    g606(.A(new_n772), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n790), .B(new_n791), .C1(new_n794), .C2(new_n771), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n771), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n770), .A2(new_n789), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G137), .ZN(G39));
  OAI21_X1  g612(.A(new_n476), .B1(new_n767), .B2(new_n768), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT47), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI211_X1 g615(.A(KEYINPUT47), .B(new_n476), .C1(new_n767), .C2(new_n768), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT111), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n730), .A2(new_n731), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n347), .A3(new_n352), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n804), .B1(new_n807), .B2(new_n736), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n806), .A2(new_n734), .A3(KEYINPUT111), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n803), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G140), .ZN(G42));
  NAND2_X1  g626(.A1(new_n706), .A2(new_n466), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n813), .A2(KEYINPUT49), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(KEYINPUT49), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n619), .A2(new_n476), .A3(new_n354), .ZN(new_n816));
  NOR4_X1   g630(.A1(new_n814), .A2(new_n815), .A3(new_n251), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n682), .A2(new_n680), .ZN(new_n818));
  AND4_X1   g632(.A1(new_n350), .A2(new_n777), .A3(new_n689), .A4(new_n778), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n712), .A2(new_n709), .A3(new_n716), .A4(new_n724), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT112), .ZN(new_n823));
  INV_X1    g637(.A(new_n607), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n546), .A2(new_n554), .A3(new_n597), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n608), .A2(new_n779), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n605), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n600), .A2(new_n823), .A3(new_n666), .A4(new_n827), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n697), .A2(new_n730), .A3(new_n599), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n827), .A2(new_n666), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT112), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n822), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n637), .A2(new_n519), .A3(new_n597), .A4(new_n699), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n833), .A2(new_n662), .A3(new_n731), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n697), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n835), .B1(new_n733), .B2(new_n749), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n714), .A2(new_n721), .A3(new_n722), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n702), .A2(new_n837), .A3(new_n700), .A4(new_n732), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT113), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n836), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n832), .A2(new_n744), .A3(new_n746), .A4(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n246), .A2(new_n659), .A3(new_n699), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT114), .B1(new_n477), .B2(new_n844), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n653), .A2(new_n659), .A3(new_n660), .A4(new_n699), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT114), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n846), .A2(new_n847), .A3(new_n476), .A4(new_n474), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(new_n718), .A3(new_n644), .A4(new_n690), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n850), .A2(new_n703), .A3(new_n675), .A4(new_n727), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT52), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n727), .A2(new_n675), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT52), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n853), .A2(new_n854), .A3(new_n703), .A4(new_n850), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n821), .B1(new_n843), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n831), .A2(new_n828), .ZN(new_n858));
  INV_X1    g672(.A(new_n822), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n858), .A2(new_n842), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n856), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n727), .A2(new_n675), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n821), .B1(new_n862), .B2(KEYINPUT52), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n860), .A2(new_n861), .A3(new_n743), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n857), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT115), .B1(new_n865), .B2(KEYINPUT54), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n858), .A2(new_n842), .A3(new_n859), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n747), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT53), .B1(new_n868), .B2(new_n861), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT53), .B1(new_n862), .B2(KEYINPUT52), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n843), .A2(new_n856), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT54), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT115), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n857), .A2(new_n864), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(G952), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n708), .A2(new_n791), .ZN(new_n877));
  INV_X1    g691(.A(new_n548), .ZN(new_n878));
  NOR4_X1   g692(.A1(new_n877), .A2(new_n251), .A3(new_n878), .A4(new_n690), .ZN(new_n879));
  INV_X1    g693(.A(new_n620), .ZN(new_n880));
  AOI211_X1 g694(.A(new_n876), .B(G953), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n878), .B1(new_n782), .B2(new_n787), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n723), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n719), .ZN(new_n885));
  AOI211_X1 g699(.A(new_n878), .B(new_n877), .C1(new_n787), .C2(new_n782), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n251), .B1(new_n339), .B2(new_n342), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT48), .ZN(new_n889));
  OR2_X1    g703(.A1(new_n889), .A2(KEYINPUT118), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n881), .B(new_n885), .C1(new_n888), .C2(new_n890), .ZN(new_n891));
  XNOR2_X1  g705(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n891), .B1(new_n888), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n813), .A2(new_n476), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n803), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n884), .A2(new_n791), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n707), .A2(new_n354), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n882), .A2(new_n818), .A3(new_n723), .A4(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT116), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT50), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n608), .A2(new_n619), .ZN(new_n904));
  AOI22_X1  g718(.A1(new_n886), .A2(new_n837), .B1(new_n879), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n899), .A2(new_n900), .A3(KEYINPUT50), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n903), .A2(new_n905), .A3(KEYINPUT51), .A4(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n893), .B1(new_n897), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n903), .A2(new_n906), .A3(new_n905), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT117), .ZN(new_n910));
  OR2_X1    g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n911), .B(new_n912), .C1(new_n895), .C2(new_n896), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT51), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n908), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AND4_X1   g729(.A1(new_n866), .A2(new_n872), .A3(new_n875), .A4(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(G952), .A2(G953), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n820), .B1(new_n916), .B2(new_n917), .ZN(G75));
  NOR2_X1   g732(.A1(new_n423), .A2(new_n425), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(new_n361), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT55), .Z(new_n921));
  NAND2_X1  g735(.A1(new_n743), .A2(new_n863), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n867), .A2(new_n856), .A3(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n860), .A2(new_n861), .A3(new_n744), .A4(new_n746), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n923), .B1(new_n924), .B2(new_n821), .ZN(new_n925));
  INV_X1    g739(.A(G210), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n925), .A2(new_n926), .A3(new_n233), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n921), .B1(new_n927), .B2(KEYINPUT56), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT56), .ZN(new_n929));
  INV_X1    g743(.A(new_n921), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n865), .A2(G902), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n929), .B(new_n930), .C1(new_n931), .C2(new_n926), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n228), .A2(G952), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n928), .A2(new_n932), .A3(new_n934), .ZN(G51));
  XOR2_X1   g749(.A(new_n467), .B(KEYINPUT57), .Z(new_n936));
  AND3_X1   g750(.A1(new_n857), .A2(new_n874), .A3(new_n864), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n874), .B1(new_n857), .B2(new_n864), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n457), .A2(new_n465), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n931), .A2(new_n763), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n933), .B1(new_n941), .B2(new_n942), .ZN(G54));
  AND2_X1   g757(.A1(KEYINPUT58), .A2(G475), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n865), .A2(G902), .A3(new_n543), .A4(new_n944), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n945), .A2(KEYINPUT119), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n865), .A2(G902), .A3(new_n944), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n933), .B1(new_n947), .B2(new_n631), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n945), .A2(KEYINPUT119), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(G60));
  NOR2_X1   g764(.A1(new_n615), .A2(new_n616), .ZN(new_n951));
  NAND2_X1  g765(.A1(G478), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT59), .Z(new_n953));
  NOR2_X1   g767(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(new_n937), .B2(new_n938), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n934), .ZN(new_n956));
  INV_X1    g770(.A(new_n953), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n872), .A2(new_n875), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n873), .B1(new_n925), .B2(new_n874), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n956), .B1(new_n951), .B2(new_n960), .ZN(G63));
  XNOR2_X1  g775(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n962));
  NAND2_X1  g776(.A1(G217), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n962), .B(new_n963), .Z(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n965), .B1(new_n857), .B2(new_n864), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n934), .B1(new_n966), .B2(new_n248), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n966), .B1(new_n658), .B2(new_n657), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n968), .A2(KEYINPUT61), .A3(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT61), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n865), .A2(new_n964), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n657), .A2(new_n658), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n971), .B1(new_n974), .B2(new_n967), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n970), .A2(new_n975), .ZN(G66));
  OAI21_X1  g790(.A(G953), .B1(new_n550), .B2(new_n358), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n977), .B1(new_n832), .B2(G953), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n919), .B1(G898), .B2(new_n228), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n978), .B(new_n979), .ZN(G69));
  INV_X1    g794(.A(KEYINPUT123), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n703), .A2(new_n695), .A3(new_n675), .A4(new_n727), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT62), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n853), .A2(KEYINPUT62), .A3(new_n695), .A4(new_n703), .ZN(new_n985));
  AOI22_X1  g799(.A1(new_n984), .A2(new_n985), .B1(new_n803), .B2(new_n810), .ZN(new_n986));
  NOR3_X1   g800(.A1(new_n477), .A2(new_n731), .A3(new_n693), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n353), .A2(new_n825), .A3(new_n826), .A4(new_n987), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n797), .A2(KEYINPUT122), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(KEYINPUT122), .B1(new_n797), .B2(new_n988), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n986), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n228), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n307), .A2(new_n308), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT121), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n523), .A2(new_n525), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n994), .B(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n981), .B1(new_n992), .B2(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(new_n996), .ZN(new_n998));
  AOI211_X1 g812(.A(KEYINPUT123), .B(new_n998), .C1(new_n991), .C2(new_n228), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n718), .A2(new_n644), .A3(new_n887), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n750), .B1(new_n770), .B2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n811), .A2(new_n744), .A3(new_n746), .A4(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n797), .A2(new_n703), .A3(new_n853), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(KEYINPUT124), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n1005), .A2(KEYINPUT124), .ZN(new_n1008));
  OAI211_X1 g822(.A(new_n1004), .B(new_n228), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n996), .B1(G900), .B2(G953), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT125), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n228), .B1(G227), .B2(G900), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  OAI211_X1 g828(.A(new_n1000), .B(new_n1011), .C1(new_n1012), .C2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n985), .A2(new_n984), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n811), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n797), .A2(new_n988), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT122), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n797), .A2(KEYINPUT122), .A3(new_n988), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1017), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n996), .B1(new_n1022), .B2(G953), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1023), .A2(KEYINPUT123), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n992), .A2(new_n981), .A3(new_n996), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1024), .A2(new_n1025), .A3(new_n1012), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1024), .A2(new_n1025), .A3(new_n1011), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1026), .A2(new_n1027), .A3(new_n1013), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1015), .A2(new_n1028), .ZN(G72));
  NAND2_X1  g843(.A1(G472), .A2(G902), .ZN(new_n1030));
  XOR2_X1   g844(.A(new_n1030), .B(KEYINPUT63), .Z(new_n1031));
  INV_X1    g845(.A(new_n1031), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1032), .B1(new_n331), .B2(new_n323), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1033), .B1(new_n869), .B2(new_n871), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1008), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1003), .B1(new_n1035), .B2(new_n1006), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1032), .B1(new_n1036), .B2(new_n832), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n309), .A2(new_n311), .ZN(new_n1038));
  XNOR2_X1  g852(.A(new_n1038), .B(KEYINPUT126), .ZN(new_n1039));
  OR2_X1    g853(.A1(new_n1039), .A2(new_n258), .ZN(new_n1040));
  OAI211_X1 g854(.A(new_n934), .B(new_n1034), .C1(new_n1037), .C2(new_n1040), .ZN(new_n1041));
  INV_X1    g855(.A(KEYINPUT127), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n1032), .B1(new_n1022), .B2(new_n832), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1039), .A2(new_n258), .ZN(new_n1044));
  OAI21_X1  g858(.A(new_n1042), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OR3_X1    g859(.A1(new_n1043), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n1041), .B1(new_n1045), .B2(new_n1046), .ZN(G57));
endmodule


