

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U548 ( .A1(G8), .A2(n746), .ZN(n794) );
  XOR2_X1 U549 ( .A(n541), .B(n540), .Z(n517) );
  XOR2_X1 U550 ( .A(KEYINPUT31), .B(n743), .Z(n518) );
  NOR2_X4 U551 ( .A1(G651), .A2(G543), .ZN(n665) );
  NAND2_X1 U552 ( .A1(n608), .A2(n607), .ZN(n709) );
  AND2_X1 U553 ( .A1(n539), .A2(G2104), .ZN(n580) );
  BUF_X2 U554 ( .A(n664), .Z(n519) );
  NOR2_X1 U555 ( .A1(n637), .A2(n529), .ZN(n664) );
  INV_X1 U556 ( .A(G2105), .ZN(n539) );
  INV_X1 U557 ( .A(n708), .ZN(n730) );
  AND2_X1 U558 ( .A1(n760), .A2(n759), .ZN(n763) );
  XNOR2_X1 U559 ( .A(n757), .B(n756), .ZN(n783) );
  NAND2_X1 U560 ( .A1(n755), .A2(n754), .ZN(n757) );
  INV_X1 U561 ( .A(KEYINPUT33), .ZN(n775) );
  BUF_X1 U562 ( .A(n580), .Z(n907) );
  INV_X1 U563 ( .A(G2104), .ZN(n542) );
  NAND2_X1 U564 ( .A1(n661), .A2(G51), .ZN(n534) );
  NOR2_X1 U565 ( .A1(G2105), .A2(G2104), .ZN(n545) );
  INV_X1 U566 ( .A(KEYINPUT23), .ZN(n550) );
  NAND2_X1 U567 ( .A1(n580), .A2(G101), .ZN(n551) );
  XOR2_X1 U568 ( .A(KEYINPUT6), .B(n536), .Z(n520) );
  OR2_X1 U569 ( .A1(n794), .A2(n793), .ZN(n521) );
  AND2_X1 U570 ( .A1(n829), .A2(n840), .ZN(n522) );
  AND2_X1 U571 ( .A1(n577), .A2(G138), .ZN(n523) );
  INV_X1 U572 ( .A(KEYINPUT27), .ZN(n715) );
  XNOR2_X1 U573 ( .A(n716), .B(n715), .ZN(n718) );
  INV_X1 U574 ( .A(KEYINPUT30), .ZN(n736) );
  INV_X1 U575 ( .A(G168), .ZN(n738) );
  NOR2_X1 U576 ( .A1(G1966), .A2(n794), .ZN(n758) );
  INV_X1 U577 ( .A(KEYINPUT32), .ZN(n756) );
  INV_X1 U578 ( .A(KEYINPUT64), .ZN(n773) );
  NAND2_X1 U579 ( .A1(n813), .A2(n703), .ZN(n708) );
  INV_X1 U580 ( .A(n837), .ZN(n829) );
  INV_X1 U581 ( .A(KEYINPUT100), .ZN(n790) );
  INV_X1 U582 ( .A(KEYINPUT86), .ZN(n540) );
  INV_X1 U583 ( .A(KEYINPUT0), .ZN(n525) );
  XNOR2_X1 U584 ( .A(n525), .B(G543), .ZN(n637) );
  INV_X1 U585 ( .A(KEYINPUT17), .ZN(n544) );
  INV_X1 U586 ( .A(KEYINPUT65), .ZN(n532) );
  BUF_X1 U587 ( .A(n577), .Z(n908) );
  XNOR2_X1 U588 ( .A(n545), .B(n544), .ZN(n577) );
  XNOR2_X1 U589 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U590 ( .A(n549), .B(KEYINPUT87), .ZN(n701) );
  BUF_X1 U591 ( .A(n701), .Z(G164) );
  NAND2_X1 U592 ( .A1(n665), .A2(G89), .ZN(n524) );
  XNOR2_X1 U593 ( .A(n524), .B(KEYINPUT4), .ZN(n527) );
  INV_X1 U594 ( .A(G651), .ZN(n529) );
  NAND2_X1 U595 ( .A1(G76), .A2(n519), .ZN(n526) );
  NAND2_X1 U596 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n528), .B(KEYINPUT5), .ZN(n537) );
  NOR2_X1 U598 ( .A1(G543), .A2(n529), .ZN(n531) );
  XNOR2_X1 U599 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n530) );
  XNOR2_X1 U600 ( .A(n531), .B(n530), .ZN(n612) );
  BUF_X1 U601 ( .A(n612), .Z(n660) );
  NAND2_X1 U602 ( .A1(G63), .A2(n660), .ZN(n535) );
  NOR2_X1 U603 ( .A1(G651), .A2(n637), .ZN(n533) );
  XNOR2_X2 U604 ( .A(n533), .B(n532), .ZN(n661) );
  NAND2_X1 U605 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U606 ( .A1(n537), .A2(n520), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n538), .B(KEYINPUT7), .ZN(G168) );
  AND2_X1 U608 ( .A1(G2105), .A2(G2104), .ZN(n911) );
  NAND2_X1 U609 ( .A1(n911), .A2(G114), .ZN(n548) );
  NAND2_X1 U610 ( .A1(G102), .A2(n580), .ZN(n541) );
  AND2_X1 U611 ( .A1(n542), .A2(G2105), .ZN(n913) );
  NAND2_X1 U612 ( .A1(G126), .A2(n913), .ZN(n543) );
  NAND2_X1 U613 ( .A1(n517), .A2(n543), .ZN(n546) );
  NOR2_X1 U614 ( .A1(n546), .A2(n523), .ZN(n547) );
  NAND2_X1 U615 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U616 ( .A1(n911), .A2(G113), .ZN(n553) );
  NAND2_X1 U617 ( .A1(n553), .A2(n552), .ZN(n557) );
  NAND2_X1 U618 ( .A1(G125), .A2(n913), .ZN(n555) );
  NAND2_X1 U619 ( .A1(G137), .A2(n577), .ZN(n554) );
  NAND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X2 U621 ( .A1(n557), .A2(n556), .ZN(G160) );
  XNOR2_X1 U622 ( .A(G2427), .B(KEYINPUT104), .ZN(n567) );
  XOR2_X1 U623 ( .A(G2430), .B(G2446), .Z(n559) );
  XNOR2_X1 U624 ( .A(KEYINPUT105), .B(G2438), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n563) );
  XOR2_X1 U626 ( .A(G2435), .B(G2454), .Z(n561) );
  XNOR2_X1 U627 ( .A(G1348), .B(G1341), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U629 ( .A(n563), .B(n562), .Z(n565) );
  XNOR2_X1 U630 ( .A(G2451), .B(G2443), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  AND2_X1 U633 ( .A1(n568), .A2(G14), .ZN(G401) );
  NAND2_X1 U634 ( .A1(G64), .A2(n660), .ZN(n570) );
  NAND2_X1 U635 ( .A1(G52), .A2(n661), .ZN(n569) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n575) );
  NAND2_X1 U637 ( .A1(G77), .A2(n519), .ZN(n572) );
  NAND2_X1 U638 ( .A1(G90), .A2(n665), .ZN(n571) );
  NAND2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U640 ( .A(KEYINPUT9), .B(n573), .Z(n574) );
  NOR2_X1 U641 ( .A1(n575), .A2(n574), .ZN(G171) );
  AND2_X1 U642 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U643 ( .A1(G123), .A2(n913), .ZN(n576) );
  XNOR2_X1 U644 ( .A(n576), .B(KEYINPUT18), .ZN(n585) );
  NAND2_X1 U645 ( .A1(G111), .A2(n911), .ZN(n579) );
  NAND2_X1 U646 ( .A1(G135), .A2(n908), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U648 ( .A1(G99), .A2(n907), .ZN(n581) );
  XNOR2_X1 U649 ( .A(KEYINPUT75), .B(n581), .ZN(n582) );
  NOR2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n944) );
  XNOR2_X1 U652 ( .A(G2096), .B(n944), .ZN(n586) );
  OR2_X1 U653 ( .A1(G2100), .A2(n586), .ZN(G156) );
  INV_X1 U654 ( .A(G57), .ZN(G237) );
  INV_X1 U655 ( .A(G69), .ZN(G235) );
  INV_X1 U656 ( .A(G108), .ZN(G238) );
  INV_X1 U657 ( .A(G120), .ZN(G236) );
  INV_X1 U658 ( .A(G132), .ZN(G219) );
  INV_X1 U659 ( .A(G82), .ZN(G220) );
  NAND2_X1 U660 ( .A1(G78), .A2(n519), .ZN(n588) );
  NAND2_X1 U661 ( .A1(G91), .A2(n665), .ZN(n587) );
  NAND2_X1 U662 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U663 ( .A(KEYINPUT68), .B(n589), .Z(n593) );
  NAND2_X1 U664 ( .A1(G65), .A2(n660), .ZN(n591) );
  NAND2_X1 U665 ( .A1(G53), .A2(n661), .ZN(n590) );
  AND2_X1 U666 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U667 ( .A1(n593), .A2(n592), .ZN(G299) );
  XOR2_X1 U668 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U669 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n595) );
  NAND2_X1 U670 ( .A1(G7), .A2(G661), .ZN(n594) );
  XNOR2_X1 U671 ( .A(n595), .B(n594), .ZN(G223) );
  XOR2_X1 U672 ( .A(KEYINPUT11), .B(KEYINPUT70), .Z(n597) );
  INV_X1 U673 ( .A(G223), .ZN(n850) );
  NAND2_X1 U674 ( .A1(G567), .A2(n850), .ZN(n596) );
  XNOR2_X1 U675 ( .A(n597), .B(n596), .ZN(G234) );
  NAND2_X1 U676 ( .A1(G68), .A2(n519), .ZN(n600) );
  NAND2_X1 U677 ( .A1(n665), .A2(G81), .ZN(n598) );
  XNOR2_X1 U678 ( .A(n598), .B(KEYINPUT12), .ZN(n599) );
  NAND2_X1 U679 ( .A1(n600), .A2(n599), .ZN(n602) );
  XNOR2_X1 U680 ( .A(KEYINPUT13), .B(KEYINPUT71), .ZN(n601) );
  XNOR2_X1 U681 ( .A(n602), .B(n601), .ZN(n605) );
  NAND2_X1 U682 ( .A1(n612), .A2(G56), .ZN(n603) );
  XOR2_X1 U683 ( .A(KEYINPUT14), .B(n603), .Z(n604) );
  NOR2_X1 U684 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U685 ( .A(n606), .B(KEYINPUT72), .ZN(n608) );
  NAND2_X1 U686 ( .A1(G43), .A2(n661), .ZN(n607) );
  INV_X1 U687 ( .A(G860), .ZN(n623) );
  OR2_X1 U688 ( .A1(n709), .A2(n623), .ZN(G153) );
  INV_X1 U689 ( .A(G171), .ZN(G301) );
  NAND2_X1 U690 ( .A1(G868), .A2(G301), .ZN(n620) );
  NAND2_X1 U691 ( .A1(G79), .A2(n519), .ZN(n609) );
  XNOR2_X1 U692 ( .A(n609), .B(KEYINPUT74), .ZN(n617) );
  NAND2_X1 U693 ( .A1(G92), .A2(n665), .ZN(n611) );
  NAND2_X1 U694 ( .A1(G54), .A2(n661), .ZN(n610) );
  NAND2_X1 U695 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U696 ( .A1(G66), .A2(n612), .ZN(n613) );
  XNOR2_X1 U697 ( .A(KEYINPUT73), .B(n613), .ZN(n614) );
  NOR2_X1 U698 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U699 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U700 ( .A(KEYINPUT15), .B(n618), .ZN(n986) );
  OR2_X1 U701 ( .A1(n986), .A2(G868), .ZN(n619) );
  NAND2_X1 U702 ( .A1(n620), .A2(n619), .ZN(G284) );
  INV_X1 U703 ( .A(G868), .ZN(n683) );
  NOR2_X1 U704 ( .A1(G286), .A2(n683), .ZN(n622) );
  NOR2_X1 U705 ( .A1(G868), .A2(G299), .ZN(n621) );
  NOR2_X1 U706 ( .A1(n622), .A2(n621), .ZN(G297) );
  NAND2_X1 U707 ( .A1(n623), .A2(G559), .ZN(n624) );
  NAND2_X1 U708 ( .A1(n624), .A2(n986), .ZN(n625) );
  XNOR2_X1 U709 ( .A(n625), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U710 ( .A1(G868), .A2(n709), .ZN(n628) );
  NAND2_X1 U711 ( .A1(G868), .A2(n986), .ZN(n626) );
  NOR2_X1 U712 ( .A1(G559), .A2(n626), .ZN(n627) );
  NOR2_X1 U713 ( .A1(n628), .A2(n627), .ZN(G282) );
  NAND2_X1 U714 ( .A1(n986), .A2(G559), .ZN(n680) );
  XNOR2_X1 U715 ( .A(n709), .B(n680), .ZN(n629) );
  NOR2_X1 U716 ( .A1(n629), .A2(G860), .ZN(n636) );
  NAND2_X1 U717 ( .A1(G80), .A2(n519), .ZN(n631) );
  NAND2_X1 U718 ( .A1(G93), .A2(n665), .ZN(n630) );
  NAND2_X1 U719 ( .A1(n631), .A2(n630), .ZN(n635) );
  NAND2_X1 U720 ( .A1(G67), .A2(n660), .ZN(n633) );
  NAND2_X1 U721 ( .A1(G55), .A2(n661), .ZN(n632) );
  NAND2_X1 U722 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U723 ( .A1(n635), .A2(n634), .ZN(n682) );
  XNOR2_X1 U724 ( .A(n636), .B(n682), .ZN(G145) );
  NAND2_X1 U725 ( .A1(G74), .A2(G651), .ZN(n642) );
  NAND2_X1 U726 ( .A1(G49), .A2(n661), .ZN(n639) );
  NAND2_X1 U727 ( .A1(G87), .A2(n637), .ZN(n638) );
  NAND2_X1 U728 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U729 ( .A1(n660), .A2(n640), .ZN(n641) );
  NAND2_X1 U730 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U731 ( .A(n643), .B(KEYINPUT76), .ZN(G288) );
  NAND2_X1 U732 ( .A1(G85), .A2(n665), .ZN(n645) );
  NAND2_X1 U733 ( .A1(G60), .A2(n660), .ZN(n644) );
  NAND2_X1 U734 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U735 ( .A1(G72), .A2(n519), .ZN(n646) );
  XOR2_X1 U736 ( .A(KEYINPUT66), .B(n646), .Z(n647) );
  NOR2_X1 U737 ( .A1(n648), .A2(n647), .ZN(n650) );
  NAND2_X1 U738 ( .A1(n661), .A2(G47), .ZN(n649) );
  NAND2_X1 U739 ( .A1(n650), .A2(n649), .ZN(G290) );
  NAND2_X1 U740 ( .A1(n660), .A2(G61), .ZN(n651) );
  XNOR2_X1 U741 ( .A(KEYINPUT77), .B(n651), .ZN(n656) );
  NAND2_X1 U742 ( .A1(n519), .A2(G73), .ZN(n652) );
  XNOR2_X1 U743 ( .A(n652), .B(KEYINPUT2), .ZN(n654) );
  NAND2_X1 U744 ( .A1(G86), .A2(n665), .ZN(n653) );
  NAND2_X1 U745 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U746 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U747 ( .A(n657), .B(KEYINPUT78), .ZN(n659) );
  NAND2_X1 U748 ( .A1(n661), .A2(G48), .ZN(n658) );
  NAND2_X1 U749 ( .A1(n659), .A2(n658), .ZN(G305) );
  NAND2_X1 U750 ( .A1(G62), .A2(n660), .ZN(n663) );
  NAND2_X1 U751 ( .A1(G50), .A2(n661), .ZN(n662) );
  NAND2_X1 U752 ( .A1(n663), .A2(n662), .ZN(n670) );
  NAND2_X1 U753 ( .A1(G75), .A2(n519), .ZN(n667) );
  NAND2_X1 U754 ( .A1(G88), .A2(n665), .ZN(n666) );
  NAND2_X1 U755 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U756 ( .A(KEYINPUT79), .B(n668), .Z(n669) );
  NOR2_X1 U757 ( .A1(n670), .A2(n669), .ZN(G166) );
  XOR2_X1 U758 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n672) );
  XNOR2_X1 U759 ( .A(KEYINPUT19), .B(KEYINPUT80), .ZN(n671) );
  XNOR2_X1 U760 ( .A(n672), .B(n671), .ZN(n674) );
  XOR2_X1 U761 ( .A(G290), .B(G299), .Z(n673) );
  XNOR2_X1 U762 ( .A(n674), .B(n673), .ZN(n676) );
  XNOR2_X1 U763 ( .A(n709), .B(n682), .ZN(n675) );
  XNOR2_X1 U764 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U765 ( .A(G288), .B(n677), .ZN(n679) );
  XNOR2_X1 U766 ( .A(G305), .B(G166), .ZN(n678) );
  XNOR2_X1 U767 ( .A(n679), .B(n678), .ZN(n859) );
  XNOR2_X1 U768 ( .A(n859), .B(n680), .ZN(n681) );
  NOR2_X1 U769 ( .A1(n683), .A2(n681), .ZN(n685) );
  AND2_X1 U770 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U771 ( .A1(n685), .A2(n684), .ZN(G295) );
  NAND2_X1 U772 ( .A1(G2078), .A2(G2084), .ZN(n686) );
  XOR2_X1 U773 ( .A(KEYINPUT20), .B(n686), .Z(n687) );
  NAND2_X1 U774 ( .A1(G2090), .A2(n687), .ZN(n688) );
  XNOR2_X1 U775 ( .A(KEYINPUT21), .B(n688), .ZN(n689) );
  NAND2_X1 U776 ( .A1(n689), .A2(G2072), .ZN(n690) );
  XOR2_X1 U777 ( .A(KEYINPUT83), .B(n690), .Z(G158) );
  XNOR2_X1 U778 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U779 ( .A1(G220), .A2(G219), .ZN(n691) );
  XOR2_X1 U780 ( .A(KEYINPUT22), .B(n691), .Z(n692) );
  NOR2_X1 U781 ( .A1(G218), .A2(n692), .ZN(n693) );
  NAND2_X1 U782 ( .A1(G96), .A2(n693), .ZN(n857) );
  NAND2_X1 U783 ( .A1(n857), .A2(G2106), .ZN(n698) );
  NOR2_X1 U784 ( .A1(G236), .A2(G238), .ZN(n695) );
  NOR2_X1 U785 ( .A1(G235), .A2(G237), .ZN(n694) );
  NAND2_X1 U786 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U787 ( .A(KEYINPUT84), .B(n696), .ZN(n858) );
  NAND2_X1 U788 ( .A1(n858), .A2(G567), .ZN(n697) );
  NAND2_X1 U789 ( .A1(n698), .A2(n697), .ZN(n932) );
  NAND2_X1 U790 ( .A1(G483), .A2(G661), .ZN(n699) );
  NOR2_X1 U791 ( .A1(n932), .A2(n699), .ZN(n856) );
  NAND2_X1 U792 ( .A1(G36), .A2(n856), .ZN(n700) );
  XOR2_X1 U793 ( .A(KEYINPUT85), .B(n700), .Z(G176) );
  XOR2_X1 U794 ( .A(KEYINPUT88), .B(G166), .Z(G303) );
  INV_X1 U795 ( .A(n701), .ZN(n813) );
  NAND2_X1 U796 ( .A1(G160), .A2(G40), .ZN(n814) );
  INV_X1 U797 ( .A(n814), .ZN(n702) );
  INV_X1 U798 ( .A(G1384), .ZN(n812) );
  AND2_X1 U799 ( .A1(n702), .A2(n812), .ZN(n703) );
  BUF_X2 U800 ( .A(n708), .Z(n746) );
  NAND2_X1 U801 ( .A1(G1348), .A2(n746), .ZN(n705) );
  NAND2_X1 U802 ( .A1(G2067), .A2(n730), .ZN(n704) );
  NAND2_X1 U803 ( .A1(n705), .A2(n704), .ZN(n714) );
  INV_X1 U804 ( .A(G1996), .ZN(n965) );
  NOR2_X1 U805 ( .A1(n708), .A2(n965), .ZN(n707) );
  INV_X1 U806 ( .A(KEYINPUT26), .ZN(n706) );
  XNOR2_X1 U807 ( .A(n707), .B(n706), .ZN(n712) );
  AND2_X1 U808 ( .A1(n708), .A2(G1341), .ZN(n710) );
  NOR2_X1 U809 ( .A1(n710), .A2(n709), .ZN(n711) );
  AND2_X1 U810 ( .A1(n712), .A2(n711), .ZN(n721) );
  NOR2_X1 U811 ( .A1(n721), .A2(n986), .ZN(n713) );
  NOR2_X1 U812 ( .A1(n714), .A2(n713), .ZN(n720) );
  NAND2_X1 U813 ( .A1(n730), .A2(G2072), .ZN(n716) );
  NAND2_X1 U814 ( .A1(G1956), .A2(n746), .ZN(n717) );
  NAND2_X1 U815 ( .A1(n718), .A2(n717), .ZN(n725) );
  NOR2_X1 U816 ( .A1(G299), .A2(n725), .ZN(n719) );
  NOR2_X1 U817 ( .A1(n720), .A2(n719), .ZN(n723) );
  NAND2_X1 U818 ( .A1(n986), .A2(n721), .ZN(n722) );
  NAND2_X1 U819 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U820 ( .A(n724), .B(KEYINPUT95), .ZN(n728) );
  NAND2_X1 U821 ( .A1(G299), .A2(n725), .ZN(n726) );
  XOR2_X1 U822 ( .A(KEYINPUT28), .B(n726), .Z(n727) );
  NOR2_X1 U823 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U824 ( .A(n729), .B(KEYINPUT29), .ZN(n734) );
  XOR2_X1 U825 ( .A(G1961), .B(KEYINPUT94), .Z(n1017) );
  NAND2_X1 U826 ( .A1(n1017), .A2(n746), .ZN(n732) );
  XNOR2_X1 U827 ( .A(G2078), .B(KEYINPUT25), .ZN(n964) );
  NAND2_X1 U828 ( .A1(n730), .A2(n964), .ZN(n731) );
  NAND2_X1 U829 ( .A1(n732), .A2(n731), .ZN(n740) );
  NAND2_X1 U830 ( .A1(G171), .A2(n740), .ZN(n733) );
  NAND2_X1 U831 ( .A1(n734), .A2(n733), .ZN(n744) );
  NOR2_X1 U832 ( .A1(G2084), .A2(n746), .ZN(n761) );
  NOR2_X1 U833 ( .A1(n758), .A2(n761), .ZN(n735) );
  NAND2_X1 U834 ( .A1(G8), .A2(n735), .ZN(n737) );
  XNOR2_X1 U835 ( .A(n737), .B(n736), .ZN(n739) );
  AND2_X1 U836 ( .A1(n739), .A2(n738), .ZN(n742) );
  NOR2_X1 U837 ( .A1(G171), .A2(n740), .ZN(n741) );
  NOR2_X1 U838 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U839 ( .A1(n744), .A2(n518), .ZN(n745) );
  XNOR2_X1 U840 ( .A(n745), .B(KEYINPUT96), .ZN(n760) );
  NAND2_X1 U841 ( .A1(n760), .A2(G286), .ZN(n755) );
  INV_X1 U842 ( .A(G8), .ZN(n753) );
  NOR2_X1 U843 ( .A1(n746), .A2(G2090), .ZN(n747) );
  XNOR2_X1 U844 ( .A(n747), .B(KEYINPUT98), .ZN(n750) );
  NOR2_X1 U845 ( .A1(G1971), .A2(n794), .ZN(n748) );
  XOR2_X1 U846 ( .A(KEYINPUT97), .B(n748), .Z(n749) );
  NOR2_X1 U847 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U848 ( .A1(n751), .A2(G303), .ZN(n752) );
  OR2_X1 U849 ( .A1(n753), .A2(n752), .ZN(n754) );
  INV_X1 U850 ( .A(n758), .ZN(n759) );
  NAND2_X1 U851 ( .A1(G8), .A2(n761), .ZN(n762) );
  NAND2_X1 U852 ( .A1(n763), .A2(n762), .ZN(n782) );
  INV_X1 U853 ( .A(n794), .ZN(n765) );
  NAND2_X1 U854 ( .A1(G1976), .A2(G288), .ZN(n764) );
  XOR2_X1 U855 ( .A(KEYINPUT99), .B(n764), .Z(n999) );
  AND2_X1 U856 ( .A1(n765), .A2(n999), .ZN(n767) );
  AND2_X1 U857 ( .A1(n782), .A2(n767), .ZN(n766) );
  NAND2_X1 U858 ( .A1(n783), .A2(n766), .ZN(n772) );
  INV_X1 U859 ( .A(n767), .ZN(n770) );
  NOR2_X1 U860 ( .A1(G288), .A2(G1976), .ZN(n998) );
  NOR2_X1 U861 ( .A1(G303), .A2(G1971), .ZN(n768) );
  NOR2_X1 U862 ( .A1(n998), .A2(n768), .ZN(n769) );
  OR2_X1 U863 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U864 ( .A1(n772), .A2(n771), .ZN(n774) );
  XNOR2_X1 U865 ( .A(n774), .B(n773), .ZN(n776) );
  NAND2_X1 U866 ( .A1(n776), .A2(n775), .ZN(n781) );
  XOR2_X1 U867 ( .A(G1981), .B(G305), .Z(n983) );
  INV_X1 U868 ( .A(n983), .ZN(n779) );
  NAND2_X1 U869 ( .A1(n998), .A2(KEYINPUT33), .ZN(n777) );
  NOR2_X1 U870 ( .A1(n777), .A2(n794), .ZN(n778) );
  NOR2_X1 U871 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U872 ( .A1(n781), .A2(n780), .ZN(n789) );
  NAND2_X1 U873 ( .A1(n782), .A2(n783), .ZN(n786) );
  NOR2_X1 U874 ( .A1(G2090), .A2(G303), .ZN(n784) );
  NAND2_X1 U875 ( .A1(G8), .A2(n784), .ZN(n785) );
  NAND2_X1 U876 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n787), .A2(n794), .ZN(n788) );
  NAND2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n791) );
  XNOR2_X1 U879 ( .A(n791), .B(n790), .ZN(n795) );
  NOR2_X1 U880 ( .A1(G1981), .A2(G305), .ZN(n792) );
  XOR2_X1 U881 ( .A(n792), .B(KEYINPUT24), .Z(n793) );
  NAND2_X1 U882 ( .A1(n795), .A2(n521), .ZN(n830) );
  NAND2_X1 U883 ( .A1(G119), .A2(n913), .ZN(n797) );
  NAND2_X1 U884 ( .A1(G107), .A2(n911), .ZN(n796) );
  NAND2_X1 U885 ( .A1(n797), .A2(n796), .ZN(n800) );
  NAND2_X1 U886 ( .A1(n907), .A2(G95), .ZN(n798) );
  XOR2_X1 U887 ( .A(KEYINPUT92), .B(n798), .Z(n799) );
  NOR2_X1 U888 ( .A1(n800), .A2(n799), .ZN(n802) );
  NAND2_X1 U889 ( .A1(n908), .A2(G131), .ZN(n801) );
  NAND2_X1 U890 ( .A1(n802), .A2(n801), .ZN(n893) );
  NAND2_X1 U891 ( .A1(G1991), .A2(n893), .ZN(n811) );
  NAND2_X1 U892 ( .A1(G129), .A2(n913), .ZN(n804) );
  NAND2_X1 U893 ( .A1(G117), .A2(n911), .ZN(n803) );
  NAND2_X1 U894 ( .A1(n804), .A2(n803), .ZN(n807) );
  NAND2_X1 U895 ( .A1(n907), .A2(G105), .ZN(n805) );
  XOR2_X1 U896 ( .A(KEYINPUT38), .B(n805), .Z(n806) );
  NOR2_X1 U897 ( .A1(n807), .A2(n806), .ZN(n809) );
  NAND2_X1 U898 ( .A1(n908), .A2(G141), .ZN(n808) );
  NAND2_X1 U899 ( .A1(n809), .A2(n808), .ZN(n890) );
  NAND2_X1 U900 ( .A1(G1996), .A2(n890), .ZN(n810) );
  NAND2_X1 U901 ( .A1(n811), .A2(n810), .ZN(n934) );
  AND2_X1 U902 ( .A1(n813), .A2(n812), .ZN(n815) );
  NOR2_X1 U903 ( .A1(n815), .A2(n814), .ZN(n845) );
  NAND2_X1 U904 ( .A1(n934), .A2(n845), .ZN(n816) );
  XNOR2_X1 U905 ( .A(n816), .B(KEYINPUT93), .ZN(n837) );
  XNOR2_X1 U906 ( .A(KEYINPUT90), .B(KEYINPUT36), .ZN(n827) );
  NAND2_X1 U907 ( .A1(G128), .A2(n913), .ZN(n818) );
  NAND2_X1 U908 ( .A1(G116), .A2(n911), .ZN(n817) );
  NAND2_X1 U909 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U910 ( .A(n819), .B(KEYINPUT35), .ZN(n825) );
  XNOR2_X1 U911 ( .A(KEYINPUT89), .B(KEYINPUT34), .ZN(n823) );
  NAND2_X1 U912 ( .A1(G104), .A2(n907), .ZN(n821) );
  NAND2_X1 U913 ( .A1(G140), .A2(n908), .ZN(n820) );
  NAND2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U915 ( .A(n823), .B(n822), .ZN(n824) );
  NAND2_X1 U916 ( .A1(n825), .A2(n824), .ZN(n826) );
  XOR2_X1 U917 ( .A(n827), .B(n826), .Z(n923) );
  XNOR2_X1 U918 ( .A(KEYINPUT37), .B(G2067), .ZN(n842) );
  OR2_X1 U919 ( .A1(n923), .A2(n842), .ZN(n828) );
  XNOR2_X1 U920 ( .A(n828), .B(KEYINPUT91), .ZN(n956) );
  NAND2_X1 U921 ( .A1(n845), .A2(n956), .ZN(n840) );
  NAND2_X1 U922 ( .A1(n830), .A2(n522), .ZN(n831) );
  XNOR2_X1 U923 ( .A(n831), .B(KEYINPUT101), .ZN(n833) );
  XNOR2_X1 U924 ( .A(G1986), .B(G290), .ZN(n991) );
  NAND2_X1 U925 ( .A1(n845), .A2(n991), .ZN(n832) );
  NAND2_X1 U926 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U927 ( .A(n834), .B(KEYINPUT102), .ZN(n848) );
  NOR2_X1 U928 ( .A1(G1996), .A2(n890), .ZN(n942) );
  NOR2_X1 U929 ( .A1(G1986), .A2(G290), .ZN(n835) );
  NOR2_X1 U930 ( .A1(G1991), .A2(n893), .ZN(n946) );
  NOR2_X1 U931 ( .A1(n835), .A2(n946), .ZN(n836) );
  NOR2_X1 U932 ( .A1(n837), .A2(n836), .ZN(n838) );
  NOR2_X1 U933 ( .A1(n942), .A2(n838), .ZN(n839) );
  XNOR2_X1 U934 ( .A(KEYINPUT39), .B(n839), .ZN(n841) );
  NAND2_X1 U935 ( .A1(n841), .A2(n840), .ZN(n843) );
  NAND2_X1 U936 ( .A1(n923), .A2(n842), .ZN(n933) );
  NAND2_X1 U937 ( .A1(n843), .A2(n933), .ZN(n844) );
  NAND2_X1 U938 ( .A1(n845), .A2(n844), .ZN(n846) );
  XOR2_X1 U939 ( .A(KEYINPUT103), .B(n846), .Z(n847) );
  NAND2_X1 U940 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U941 ( .A(n849), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U942 ( .A1(G2106), .A2(n850), .ZN(G217) );
  INV_X1 U943 ( .A(G661), .ZN(n852) );
  NAND2_X1 U944 ( .A1(G2), .A2(G15), .ZN(n851) );
  NOR2_X1 U945 ( .A1(n852), .A2(n851), .ZN(n853) );
  XOR2_X1 U946 ( .A(KEYINPUT106), .B(n853), .Z(G259) );
  NAND2_X1 U947 ( .A1(G3), .A2(G1), .ZN(n854) );
  XOR2_X1 U948 ( .A(KEYINPUT107), .B(n854), .Z(n855) );
  NAND2_X1 U949 ( .A1(n856), .A2(n855), .ZN(G188) );
  INV_X1 U951 ( .A(G96), .ZN(G221) );
  NOR2_X1 U952 ( .A1(n858), .A2(n857), .ZN(G325) );
  INV_X1 U953 ( .A(G325), .ZN(G261) );
  XOR2_X1 U954 ( .A(n859), .B(G286), .Z(n861) );
  XNOR2_X1 U955 ( .A(G171), .B(n986), .ZN(n860) );
  XNOR2_X1 U956 ( .A(n861), .B(n860), .ZN(n862) );
  NOR2_X1 U957 ( .A1(G37), .A2(n862), .ZN(G397) );
  XNOR2_X1 U958 ( .A(G1996), .B(KEYINPUT41), .ZN(n872) );
  XOR2_X1 U959 ( .A(G1971), .B(G1961), .Z(n864) );
  XNOR2_X1 U960 ( .A(G1991), .B(G1986), .ZN(n863) );
  XNOR2_X1 U961 ( .A(n864), .B(n863), .ZN(n868) );
  XOR2_X1 U962 ( .A(G1976), .B(G1956), .Z(n866) );
  XNOR2_X1 U963 ( .A(G1981), .B(G1966), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U965 ( .A(n868), .B(n867), .Z(n870) );
  XNOR2_X1 U966 ( .A(KEYINPUT110), .B(G2474), .ZN(n869) );
  XNOR2_X1 U967 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U968 ( .A(n872), .B(n871), .ZN(G229) );
  XOR2_X1 U969 ( .A(KEYINPUT109), .B(G2678), .Z(n874) );
  XNOR2_X1 U970 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n873) );
  XNOR2_X1 U971 ( .A(n874), .B(n873), .ZN(n878) );
  XOR2_X1 U972 ( .A(KEYINPUT42), .B(G2072), .Z(n876) );
  XNOR2_X1 U973 ( .A(G2067), .B(G2090), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U975 ( .A(n878), .B(n877), .Z(n880) );
  XNOR2_X1 U976 ( .A(G2096), .B(G2100), .ZN(n879) );
  XNOR2_X1 U977 ( .A(n880), .B(n879), .ZN(n882) );
  XOR2_X1 U978 ( .A(G2078), .B(G2084), .Z(n881) );
  XNOR2_X1 U979 ( .A(n882), .B(n881), .ZN(G227) );
  NAND2_X1 U980 ( .A1(n913), .A2(G124), .ZN(n883) );
  XNOR2_X1 U981 ( .A(n883), .B(KEYINPUT44), .ZN(n885) );
  NAND2_X1 U982 ( .A1(G112), .A2(n911), .ZN(n884) );
  NAND2_X1 U983 ( .A1(n885), .A2(n884), .ZN(n889) );
  NAND2_X1 U984 ( .A1(G100), .A2(n907), .ZN(n887) );
  NAND2_X1 U985 ( .A1(G136), .A2(n908), .ZN(n886) );
  NAND2_X1 U986 ( .A1(n887), .A2(n886), .ZN(n888) );
  NOR2_X1 U987 ( .A1(n889), .A2(n888), .ZN(G162) );
  XNOR2_X1 U988 ( .A(G162), .B(n890), .ZN(n891) );
  XNOR2_X1 U989 ( .A(n891), .B(n944), .ZN(n898) );
  XOR2_X1 U990 ( .A(KEYINPUT48), .B(KEYINPUT112), .Z(n892) );
  XNOR2_X1 U991 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U992 ( .A(n894), .B(KEYINPUT46), .Z(n896) );
  XNOR2_X1 U993 ( .A(G164), .B(KEYINPUT114), .ZN(n895) );
  XNOR2_X1 U994 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U995 ( .A(n898), .B(n897), .Z(n922) );
  NAND2_X1 U996 ( .A1(G106), .A2(n907), .ZN(n900) );
  NAND2_X1 U997 ( .A1(G142), .A2(n908), .ZN(n899) );
  NAND2_X1 U998 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n901), .B(KEYINPUT45), .ZN(n906) );
  NAND2_X1 U1000 ( .A1(G130), .A2(n913), .ZN(n903) );
  NAND2_X1 U1001 ( .A1(G118), .A2(n911), .ZN(n902) );
  NAND2_X1 U1002 ( .A1(n903), .A2(n902), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(KEYINPUT111), .B(n904), .ZN(n905) );
  NAND2_X1 U1004 ( .A1(n906), .A2(n905), .ZN(n919) );
  NAND2_X1 U1005 ( .A1(G103), .A2(n907), .ZN(n910) );
  NAND2_X1 U1006 ( .A1(G139), .A2(n908), .ZN(n909) );
  NAND2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(n918) );
  NAND2_X1 U1008 ( .A1(n911), .A2(G115), .ZN(n912) );
  XOR2_X1 U1009 ( .A(KEYINPUT113), .B(n912), .Z(n915) );
  NAND2_X1 U1010 ( .A1(n913), .A2(G127), .ZN(n914) );
  NAND2_X1 U1011 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1012 ( .A(KEYINPUT47), .B(n916), .Z(n917) );
  NOR2_X1 U1013 ( .A1(n918), .A2(n917), .ZN(n936) );
  XNOR2_X1 U1014 ( .A(n919), .B(n936), .ZN(n920) );
  XNOR2_X1 U1015 ( .A(G160), .B(n920), .ZN(n921) );
  XNOR2_X1 U1016 ( .A(n922), .B(n921), .ZN(n924) );
  XOR2_X1 U1017 ( .A(n924), .B(n923), .Z(n925) );
  NOR2_X1 U1018 ( .A1(G37), .A2(n925), .ZN(G395) );
  NOR2_X1 U1019 ( .A1(G401), .A2(n932), .ZN(n929) );
  NOR2_X1 U1020 ( .A1(G229), .A2(G227), .ZN(n926) );
  XNOR2_X1 U1021 ( .A(KEYINPUT49), .B(n926), .ZN(n927) );
  NOR2_X1 U1022 ( .A1(G397), .A2(n927), .ZN(n928) );
  NAND2_X1 U1023 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1024 ( .A1(n930), .A2(G395), .ZN(n931) );
  XNOR2_X1 U1025 ( .A(n931), .B(KEYINPUT115), .ZN(G225) );
  XOR2_X1 U1026 ( .A(KEYINPUT116), .B(G225), .Z(G308) );
  INV_X1 U1027 ( .A(n932), .ZN(G319) );
  INV_X1 U1028 ( .A(n933), .ZN(n935) );
  NOR2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n954) );
  XNOR2_X1 U1030 ( .A(G2072), .B(n936), .ZN(n939) );
  XNOR2_X1 U1031 ( .A(G164), .B(G2078), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(n937), .B(KEYINPUT118), .ZN(n938) );
  NAND2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1034 ( .A(n940), .B(KEYINPUT50), .ZN(n952) );
  XOR2_X1 U1035 ( .A(G2090), .B(G162), .Z(n941) );
  NOR2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1037 ( .A(KEYINPUT51), .B(n943), .Z(n950) );
  XNOR2_X1 U1038 ( .A(G160), .B(G2084), .ZN(n945) );
  NAND2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n947) );
  NOR2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1041 ( .A(KEYINPUT117), .B(n948), .Z(n949) );
  NAND2_X1 U1042 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1043 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1044 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1045 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1046 ( .A(KEYINPUT52), .B(n957), .Z(n958) );
  NOR2_X1 U1047 ( .A1(KEYINPUT55), .A2(n958), .ZN(n959) );
  XNOR2_X1 U1048 ( .A(KEYINPUT119), .B(n959), .ZN(n960) );
  NAND2_X1 U1049 ( .A1(n960), .A2(G29), .ZN(n1040) );
  XNOR2_X1 U1050 ( .A(G29), .B(KEYINPUT121), .ZN(n981) );
  XOR2_X1 U1051 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n979) );
  XNOR2_X1 U1052 ( .A(G2090), .B(G35), .ZN(n974) );
  XOR2_X1 U1053 ( .A(G1991), .B(G25), .Z(n961) );
  NAND2_X1 U1054 ( .A1(n961), .A2(G28), .ZN(n971) );
  XNOR2_X1 U1055 ( .A(G2067), .B(G26), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(G33), .B(G2072), .ZN(n962) );
  NOR2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n969) );
  XOR2_X1 U1058 ( .A(n964), .B(G27), .Z(n967) );
  XOR2_X1 U1059 ( .A(n965), .B(G32), .Z(n966) );
  NOR2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1063 ( .A(KEYINPUT53), .B(n972), .ZN(n973) );
  NOR2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n977) );
  XOR2_X1 U1065 ( .A(G2084), .B(G34), .Z(n975) );
  XNOR2_X1 U1066 ( .A(KEYINPUT54), .B(n975), .ZN(n976) );
  NAND2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1068 ( .A(n979), .B(n978), .ZN(n980) );
  NAND2_X1 U1069 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1070 ( .A1(n982), .A2(G11), .ZN(n1038) );
  XNOR2_X1 U1071 ( .A(G16), .B(KEYINPUT56), .ZN(n1007) );
  XNOR2_X1 U1072 ( .A(G168), .B(G1966), .ZN(n984) );
  NAND2_X1 U1073 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1074 ( .A(n985), .B(KEYINPUT57), .ZN(n1005) );
  XOR2_X1 U1075 ( .A(G1348), .B(n986), .Z(n988) );
  XNOR2_X1 U1076 ( .A(n709), .B(G1341), .ZN(n987) );
  NOR2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n997) );
  XNOR2_X1 U1078 ( .A(G1971), .B(G303), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(n989), .B(KEYINPUT123), .ZN(n993) );
  XNOR2_X1 U1080 ( .A(G1961), .B(G301), .ZN(n990) );
  NOR2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n995) );
  XNOR2_X1 U1083 ( .A(G1956), .B(G299), .ZN(n994) );
  NOR2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n1003) );
  INV_X1 U1086 ( .A(n998), .ZN(n1000) );
  NAND2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(KEYINPUT122), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1089 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1090 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1091 ( .A1(n1007), .A2(n1006), .ZN(n1036) );
  INV_X1 U1092 ( .A(G16), .ZN(n1034) );
  XNOR2_X1 U1093 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n1032) );
  XOR2_X1 U1094 ( .A(G1956), .B(G20), .Z(n1012) );
  XNOR2_X1 U1095 ( .A(G1981), .B(G6), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(G1341), .B(G19), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(KEYINPUT124), .B(n1010), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1015) );
  XOR2_X1 U1100 ( .A(KEYINPUT59), .B(G1348), .Z(n1013) );
  XNOR2_X1 U1101 ( .A(G4), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(KEYINPUT60), .B(n1016), .ZN(n1019) );
  XNOR2_X1 U1104 ( .A(n1017), .B(G5), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(G21), .B(G1966), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1108 ( .A(KEYINPUT125), .B(n1022), .Z(n1030) );
  XOR2_X1 U1109 ( .A(G1971), .B(G22), .Z(n1025) );
  XOR2_X1 U1110 ( .A(G23), .B(KEYINPUT126), .Z(n1023) );
  XNOR2_X1 U1111 ( .A(n1023), .B(G1976), .ZN(n1024) );
  NAND2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1027) );
  XNOR2_X1 U1113 ( .A(G24), .B(G1986), .ZN(n1026) );
  NOR2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1115 ( .A(KEYINPUT58), .B(n1028), .ZN(n1029) );
  NAND2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1117 ( .A(n1032), .B(n1031), .ZN(n1033) );
  NAND2_X1 U1118 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1119 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NOR2_X1 U1120 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NAND2_X1 U1121 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XOR2_X1 U1122 ( .A(KEYINPUT62), .B(n1041), .Z(G311) );
  INV_X1 U1123 ( .A(G311), .ZN(G150) );
endmodule

