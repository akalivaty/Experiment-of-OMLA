

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589;

  NOR2_X2 U323 ( .A1(n587), .A2(n541), .ZN(n388) );
  XNOR2_X1 U324 ( .A(KEYINPUT47), .B(KEYINPUT109), .ZN(n385) );
  XNOR2_X1 U325 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n394) );
  XNOR2_X1 U326 ( .A(n328), .B(KEYINPUT71), .ZN(n291) );
  XNOR2_X1 U327 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U328 ( .A(n319), .B(n318), .ZN(n322) );
  XNOR2_X1 U329 ( .A(n386), .B(n385), .ZN(n393) );
  XNOR2_X1 U330 ( .A(n416), .B(n291), .ZN(n329) );
  XNOR2_X1 U331 ( .A(n395), .B(n394), .ZN(n528) );
  XNOR2_X1 U332 ( .A(n330), .B(n329), .ZN(n387) );
  INV_X1 U333 ( .A(G190GAT), .ZN(n452) );
  XOR2_X1 U334 ( .A(n310), .B(n446), .Z(n529) );
  XNOR2_X1 U335 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U336 ( .A(n455), .B(n454), .ZN(G1351GAT) );
  INV_X1 U337 ( .A(KEYINPUT121), .ZN(n451) );
  XOR2_X1 U338 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n293) );
  XNOR2_X1 U339 ( .A(KEYINPUT81), .B(G183GAT), .ZN(n292) );
  XNOR2_X1 U340 ( .A(n293), .B(n292), .ZN(n294) );
  XNOR2_X1 U341 ( .A(KEYINPUT18), .B(n294), .ZN(n406) );
  XOR2_X1 U342 ( .A(KEYINPUT20), .B(G99GAT), .Z(n296) );
  XNOR2_X1 U343 ( .A(G43GAT), .B(G190GAT), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U345 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n298) );
  XNOR2_X1 U346 ( .A(G169GAT), .B(G15GAT), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U348 ( .A(n300), .B(n299), .Z(n305) );
  XOR2_X1 U349 ( .A(G120GAT), .B(G71GAT), .Z(n328) );
  XOR2_X1 U350 ( .A(KEYINPUT82), .B(G176GAT), .Z(n302) );
  NAND2_X1 U351 ( .A1(G227GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U352 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U353 ( .A(n328), .B(n303), .ZN(n304) );
  XNOR2_X1 U354 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U355 ( .A(n406), .B(n306), .Z(n310) );
  XOR2_X1 U356 ( .A(KEYINPUT0), .B(G134GAT), .Z(n308) );
  XNOR2_X1 U357 ( .A(KEYINPUT78), .B(G127GAT), .ZN(n307) );
  XNOR2_X1 U358 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U359 ( .A(G113GAT), .B(n309), .Z(n446) );
  XNOR2_X1 U360 ( .A(G176GAT), .B(G92GAT), .ZN(n311) );
  XNOR2_X1 U361 ( .A(n311), .B(G64GAT), .ZN(n399) );
  INV_X1 U362 ( .A(n399), .ZN(n312) );
  XOR2_X1 U363 ( .A(G99GAT), .B(G85GAT), .Z(n351) );
  NAND2_X1 U364 ( .A1(n312), .A2(n351), .ZN(n315) );
  INV_X1 U365 ( .A(n351), .ZN(n313) );
  NAND2_X1 U366 ( .A1(n399), .A2(n313), .ZN(n314) );
  NAND2_X1 U367 ( .A1(n315), .A2(n314), .ZN(n319) );
  NAND2_X1 U368 ( .A1(G230GAT), .A2(G233GAT), .ZN(n317) );
  INV_X1 U369 ( .A(KEYINPUT31), .ZN(n316) );
  XNOR2_X1 U370 ( .A(G57GAT), .B(KEYINPUT68), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n320), .B(KEYINPUT13), .ZN(n367) );
  XNOR2_X1 U372 ( .A(n367), .B(KEYINPUT33), .ZN(n321) );
  XNOR2_X1 U373 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U374 ( .A(n323), .B(KEYINPUT32), .ZN(n330) );
  XNOR2_X1 U375 ( .A(G148GAT), .B(KEYINPUT70), .ZN(n324) );
  XNOR2_X1 U376 ( .A(n324), .B(KEYINPUT69), .ZN(n325) );
  XOR2_X1 U377 ( .A(n325), .B(G204GAT), .Z(n327) );
  XNOR2_X1 U378 ( .A(G78GAT), .B(G106GAT), .ZN(n326) );
  XOR2_X1 U379 ( .A(n327), .B(n326), .Z(n416) );
  XOR2_X1 U380 ( .A(KEYINPUT41), .B(n387), .Z(n563) );
  XOR2_X1 U381 ( .A(KEYINPUT67), .B(KEYINPUT7), .Z(n332) );
  XNOR2_X1 U382 ( .A(G43GAT), .B(G29GAT), .ZN(n331) );
  XNOR2_X1 U383 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U384 ( .A(KEYINPUT8), .B(n333), .Z(n362) );
  XOR2_X1 U385 ( .A(G169GAT), .B(G8GAT), .Z(n396) );
  XOR2_X1 U386 ( .A(n396), .B(KEYINPUT29), .Z(n335) );
  NAND2_X1 U387 ( .A1(G229GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U389 ( .A(G15GAT), .B(G1GAT), .Z(n372) );
  XOR2_X1 U390 ( .A(n336), .B(n372), .Z(n344) );
  XOR2_X1 U391 ( .A(G22GAT), .B(G113GAT), .Z(n338) );
  XNOR2_X1 U392 ( .A(G36GAT), .B(G50GAT), .ZN(n337) );
  XNOR2_X1 U393 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U394 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n340) );
  XNOR2_X1 U395 ( .A(G141GAT), .B(G197GAT), .ZN(n339) );
  XNOR2_X1 U396 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U397 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U398 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U399 ( .A(n362), .B(n345), .Z(n533) );
  INV_X1 U400 ( .A(n533), .ZN(n574) );
  AND2_X1 U401 ( .A1(n563), .A2(n574), .ZN(n347) );
  XNOR2_X1 U402 ( .A(KEYINPUT46), .B(KEYINPUT108), .ZN(n346) );
  XNOR2_X1 U403 ( .A(n347), .B(n346), .ZN(n384) );
  XOR2_X1 U404 ( .A(KEYINPUT74), .B(KEYINPUT9), .Z(n349) );
  XNOR2_X1 U405 ( .A(KEYINPUT72), .B(KEYINPUT10), .ZN(n348) );
  XNOR2_X1 U406 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U407 ( .A(n350), .B(G92GAT), .Z(n353) );
  XNOR2_X1 U408 ( .A(G106GAT), .B(n351), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n358) );
  XNOR2_X1 U410 ( .A(G36GAT), .B(G190GAT), .ZN(n354) );
  XNOR2_X1 U411 ( .A(n354), .B(G218GAT), .ZN(n403) );
  XOR2_X1 U412 ( .A(G50GAT), .B(G162GAT), .Z(n412) );
  XOR2_X1 U413 ( .A(n403), .B(n412), .Z(n356) );
  NAND2_X1 U414 ( .A1(G232GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U416 ( .A(n358), .B(n357), .Z(n364) );
  XOR2_X1 U417 ( .A(KEYINPUT65), .B(KEYINPUT73), .Z(n360) );
  XNOR2_X1 U418 ( .A(G134GAT), .B(KEYINPUT11), .ZN(n359) );
  XNOR2_X1 U419 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U421 ( .A(n364), .B(n363), .Z(n545) );
  XOR2_X1 U422 ( .A(G78GAT), .B(G71GAT), .Z(n366) );
  XNOR2_X1 U423 ( .A(G183GAT), .B(G127GAT), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n366), .B(n365), .ZN(n371) );
  XOR2_X1 U425 ( .A(n367), .B(KEYINPUT12), .Z(n369) );
  NAND2_X1 U426 ( .A1(G231GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U427 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U428 ( .A(n371), .B(n370), .Z(n374) );
  XOR2_X1 U429 ( .A(G22GAT), .B(G155GAT), .Z(n411) );
  XNOR2_X1 U430 ( .A(n372), .B(n411), .ZN(n373) );
  XNOR2_X1 U431 ( .A(n374), .B(n373), .ZN(n382) );
  XOR2_X1 U432 ( .A(KEYINPUT77), .B(G64GAT), .Z(n376) );
  XNOR2_X1 U433 ( .A(G8GAT), .B(G211GAT), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n376), .B(n375), .ZN(n380) );
  XOR2_X1 U435 ( .A(KEYINPUT76), .B(KEYINPUT75), .Z(n378) );
  XNOR2_X1 U436 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n377) );
  XNOR2_X1 U437 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U438 ( .A(n380), .B(n379), .Z(n381) );
  XOR2_X1 U439 ( .A(n382), .B(n381), .Z(n582) );
  INV_X1 U440 ( .A(n582), .ZN(n541) );
  NAND2_X1 U441 ( .A1(n545), .A2(n541), .ZN(n383) );
  OR2_X1 U442 ( .A1(n384), .A2(n383), .ZN(n386) );
  XNOR2_X1 U443 ( .A(n545), .B(KEYINPUT36), .ZN(n587) );
  XOR2_X1 U444 ( .A(KEYINPUT45), .B(n388), .Z(n389) );
  NOR2_X1 U445 ( .A1(n387), .A2(n389), .ZN(n390) );
  XNOR2_X1 U446 ( .A(KEYINPUT110), .B(n390), .ZN(n391) );
  NAND2_X1 U447 ( .A1(n391), .A2(n533), .ZN(n392) );
  NAND2_X1 U448 ( .A1(n393), .A2(n392), .ZN(n395) );
  XOR2_X1 U449 ( .A(G204GAT), .B(n396), .Z(n398) );
  NAND2_X1 U450 ( .A1(G226GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U451 ( .A(n398), .B(n397), .ZN(n400) );
  XOR2_X1 U452 ( .A(n400), .B(n399), .Z(n405) );
  XOR2_X1 U453 ( .A(G211GAT), .B(KEYINPUT84), .Z(n402) );
  XNOR2_X1 U454 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n401) );
  XNOR2_X1 U455 ( .A(n402), .B(n401), .ZN(n425) );
  XNOR2_X1 U456 ( .A(n425), .B(n403), .ZN(n404) );
  XNOR2_X1 U457 ( .A(n405), .B(n404), .ZN(n407) );
  XOR2_X1 U458 ( .A(n407), .B(n406), .Z(n505) );
  INV_X1 U459 ( .A(n505), .ZN(n518) );
  AND2_X1 U460 ( .A1(n528), .A2(n518), .ZN(n410) );
  XNOR2_X1 U461 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n408) );
  XOR2_X1 U462 ( .A(n408), .B(KEYINPUT119), .Z(n409) );
  XNOR2_X1 U463 ( .A(n410), .B(n409), .ZN(n571) );
  XOR2_X1 U464 ( .A(KEYINPUT24), .B(G218GAT), .Z(n414) );
  XNOR2_X1 U465 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U466 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U467 ( .A(n416), .B(n415), .ZN(n418) );
  NAND2_X1 U468 ( .A1(G228GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U469 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U470 ( .A(KEYINPUT86), .B(KEYINPUT83), .Z(n420) );
  XNOR2_X1 U471 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n419) );
  XNOR2_X1 U472 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U473 ( .A(n422), .B(n421), .Z(n427) );
  XOR2_X1 U474 ( .A(KEYINPUT2), .B(KEYINPUT85), .Z(n424) );
  XNOR2_X1 U475 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n423) );
  XNOR2_X1 U476 ( .A(n424), .B(n423), .ZN(n437) );
  XNOR2_X1 U477 ( .A(n437), .B(n425), .ZN(n426) );
  XNOR2_X1 U478 ( .A(n427), .B(n426), .ZN(n466) );
  XOR2_X1 U479 ( .A(KEYINPUT5), .B(KEYINPUT88), .Z(n429) );
  NAND2_X1 U480 ( .A1(G225GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U481 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U482 ( .A(KEYINPUT4), .B(n430), .ZN(n444) );
  XOR2_X1 U483 ( .A(KEYINPUT1), .B(KEYINPUT87), .Z(n432) );
  XNOR2_X1 U484 ( .A(G148GAT), .B(G155GAT), .ZN(n431) );
  XNOR2_X1 U485 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U486 ( .A(KEYINPUT89), .B(G57GAT), .Z(n434) );
  XNOR2_X1 U487 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n433) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U489 ( .A(n436), .B(n435), .Z(n442) );
  XOR2_X1 U490 ( .A(G85GAT), .B(G162GAT), .Z(n439) );
  XNOR2_X1 U491 ( .A(G29GAT), .B(n437), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U493 ( .A(G120GAT), .B(n440), .ZN(n441) );
  XNOR2_X1 U494 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U495 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U496 ( .A(n446), .B(n445), .Z(n516) );
  NOR2_X1 U497 ( .A1(n466), .A2(n516), .ZN(n447) );
  AND2_X1 U498 ( .A1(n571), .A2(n447), .ZN(n448) );
  XNOR2_X1 U499 ( .A(n448), .B(KEYINPUT55), .ZN(n449) );
  NOR2_X1 U500 ( .A1(n529), .A2(n449), .ZN(n450) );
  XNOR2_X1 U501 ( .A(n451), .B(n450), .ZN(n567) );
  INV_X1 U502 ( .A(n545), .ZN(n557) );
  NAND2_X1 U503 ( .A1(n567), .A2(n557), .ZN(n455) );
  XOR2_X1 U504 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n453) );
  XOR2_X1 U505 ( .A(KEYINPUT34), .B(KEYINPUT95), .Z(n457) );
  XNOR2_X1 U506 ( .A(G1GAT), .B(KEYINPUT94), .ZN(n456) );
  XNOR2_X1 U507 ( .A(n457), .B(n456), .ZN(n476) );
  INV_X1 U508 ( .A(n516), .ZN(n570) );
  NOR2_X1 U509 ( .A1(n533), .A2(n387), .ZN(n487) );
  NOR2_X1 U510 ( .A1(n529), .A2(n505), .ZN(n458) );
  NOR2_X1 U511 ( .A1(n466), .A2(n458), .ZN(n459) );
  XOR2_X1 U512 ( .A(n459), .B(KEYINPUT25), .Z(n460) );
  XNOR2_X1 U513 ( .A(KEYINPUT92), .B(n460), .ZN(n464) );
  XOR2_X1 U514 ( .A(KEYINPUT91), .B(KEYINPUT26), .Z(n462) );
  NAND2_X1 U515 ( .A1(n466), .A2(n529), .ZN(n461) );
  XNOR2_X1 U516 ( .A(n462), .B(n461), .ZN(n573) );
  XNOR2_X1 U517 ( .A(n505), .B(KEYINPUT27), .ZN(n467) );
  NOR2_X1 U518 ( .A1(n573), .A2(n467), .ZN(n463) );
  NOR2_X1 U519 ( .A1(n464), .A2(n463), .ZN(n465) );
  NOR2_X1 U520 ( .A1(n516), .A2(n465), .ZN(n471) );
  INV_X1 U521 ( .A(n529), .ZN(n521) );
  XNOR2_X1 U522 ( .A(n466), .B(KEYINPUT28), .ZN(n524) );
  INV_X1 U523 ( .A(n524), .ZN(n531) );
  NOR2_X1 U524 ( .A1(n570), .A2(n467), .ZN(n468) );
  XNOR2_X1 U525 ( .A(n468), .B(KEYINPUT90), .ZN(n527) );
  NAND2_X1 U526 ( .A1(n531), .A2(n527), .ZN(n469) );
  NOR2_X1 U527 ( .A1(n521), .A2(n469), .ZN(n470) );
  NOR2_X1 U528 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U529 ( .A(KEYINPUT93), .B(n472), .ZN(n485) );
  NAND2_X1 U530 ( .A1(n582), .A2(n545), .ZN(n473) );
  XOR2_X1 U531 ( .A(KEYINPUT16), .B(n473), .Z(n474) );
  AND2_X1 U532 ( .A1(n485), .A2(n474), .ZN(n499) );
  NAND2_X1 U533 ( .A1(n487), .A2(n499), .ZN(n481) );
  NOR2_X1 U534 ( .A1(n570), .A2(n481), .ZN(n475) );
  XOR2_X1 U535 ( .A(n476), .B(n475), .Z(G1324GAT) );
  NOR2_X1 U536 ( .A1(n505), .A2(n481), .ZN(n477) );
  XOR2_X1 U537 ( .A(KEYINPUT96), .B(n477), .Z(n478) );
  XNOR2_X1 U538 ( .A(G8GAT), .B(n478), .ZN(G1325GAT) );
  NOR2_X1 U539 ( .A1(n529), .A2(n481), .ZN(n480) );
  XNOR2_X1 U540 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n480), .B(n479), .ZN(G1326GAT) );
  NOR2_X1 U542 ( .A1(n531), .A2(n481), .ZN(n483) );
  XNOR2_X1 U543 ( .A(G22GAT), .B(KEYINPUT97), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n483), .B(n482), .ZN(G1327GAT) );
  NOR2_X1 U545 ( .A1(n582), .A2(n587), .ZN(n484) );
  NAND2_X1 U546 ( .A1(n485), .A2(n484), .ZN(n486) );
  XNOR2_X1 U547 ( .A(KEYINPUT37), .B(n486), .ZN(n513) );
  NAND2_X1 U548 ( .A1(n487), .A2(n513), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n488), .B(KEYINPUT38), .ZN(n496) );
  NOR2_X1 U550 ( .A1(n496), .A2(n570), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n489), .B(KEYINPUT39), .ZN(n490) );
  XNOR2_X1 U552 ( .A(G29GAT), .B(n490), .ZN(G1328GAT) );
  NOR2_X1 U553 ( .A1(n496), .A2(n505), .ZN(n491) );
  XOR2_X1 U554 ( .A(KEYINPUT98), .B(n491), .Z(n492) );
  XNOR2_X1 U555 ( .A(G36GAT), .B(n492), .ZN(G1329GAT) );
  NOR2_X1 U556 ( .A1(n496), .A2(n529), .ZN(n494) );
  XNOR2_X1 U557 ( .A(KEYINPUT99), .B(KEYINPUT40), .ZN(n493) );
  XNOR2_X1 U558 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  NOR2_X1 U560 ( .A1(n531), .A2(n496), .ZN(n497) );
  XOR2_X1 U561 ( .A(KEYINPUT100), .B(n497), .Z(n498) );
  XNOR2_X1 U562 ( .A(G50GAT), .B(n498), .ZN(G1331GAT) );
  INV_X1 U563 ( .A(n563), .ZN(n537) );
  NOR2_X1 U564 ( .A1(n537), .A2(n574), .ZN(n514) );
  NAND2_X1 U565 ( .A1(n514), .A2(n499), .ZN(n508) );
  NOR2_X1 U566 ( .A1(n570), .A2(n508), .ZN(n504) );
  XOR2_X1 U567 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n501) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n500) );
  XNOR2_X1 U569 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U570 ( .A(KEYINPUT101), .B(n502), .ZN(n503) );
  XNOR2_X1 U571 ( .A(n504), .B(n503), .ZN(G1332GAT) );
  NOR2_X1 U572 ( .A1(n505), .A2(n508), .ZN(n506) );
  XOR2_X1 U573 ( .A(G64GAT), .B(n506), .Z(G1333GAT) );
  NOR2_X1 U574 ( .A1(n529), .A2(n508), .ZN(n507) );
  XOR2_X1 U575 ( .A(G71GAT), .B(n507), .Z(G1334GAT) );
  NOR2_X1 U576 ( .A1(n508), .A2(n531), .ZN(n512) );
  XOR2_X1 U577 ( .A(KEYINPUT105), .B(KEYINPUT43), .Z(n510) );
  XNOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT104), .ZN(n509) );
  XNOR2_X1 U579 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U580 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  NAND2_X1 U581 ( .A1(n514), .A2(n513), .ZN(n515) );
  XOR2_X1 U582 ( .A(KEYINPUT106), .B(n515), .Z(n523) );
  NAND2_X1 U583 ( .A1(n516), .A2(n523), .ZN(n517) );
  XNOR2_X1 U584 ( .A(G85GAT), .B(n517), .ZN(G1336GAT) );
  XOR2_X1 U585 ( .A(G92GAT), .B(KEYINPUT107), .Z(n520) );
  NAND2_X1 U586 ( .A1(n518), .A2(n523), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n520), .B(n519), .ZN(G1337GAT) );
  NAND2_X1 U588 ( .A1(n523), .A2(n521), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n522), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U590 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n526) );
  NAND2_X1 U591 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(G1339GAT) );
  NAND2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n549) );
  NOR2_X1 U594 ( .A1(n529), .A2(n549), .ZN(n530) );
  NAND2_X1 U595 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U596 ( .A(KEYINPUT111), .B(n532), .Z(n544) );
  NOR2_X1 U597 ( .A1(n533), .A2(n544), .ZN(n535) );
  XNOR2_X1 U598 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U600 ( .A(G113GAT), .B(n536), .ZN(G1340GAT) );
  NOR2_X1 U601 ( .A1(n537), .A2(n544), .ZN(n539) );
  XNOR2_X1 U602 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U604 ( .A(G120GAT), .B(n540), .ZN(G1341GAT) );
  NOR2_X1 U605 ( .A1(n541), .A2(n544), .ZN(n542) );
  XOR2_X1 U606 ( .A(KEYINPUT50), .B(n542), .Z(n543) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  NOR2_X1 U608 ( .A1(n545), .A2(n544), .ZN(n547) );
  XNOR2_X1 U609 ( .A(KEYINPUT115), .B(KEYINPUT51), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U611 ( .A(G134GAT), .B(n548), .Z(G1343GAT) );
  NOR2_X1 U612 ( .A1(n573), .A2(n549), .ZN(n558) );
  NAND2_X1 U613 ( .A1(n558), .A2(n574), .ZN(n550) );
  XNOR2_X1 U614 ( .A(G141GAT), .B(n550), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT117), .Z(n552) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U618 ( .A(KEYINPUT116), .B(n553), .Z(n555) );
  NAND2_X1 U619 ( .A1(n558), .A2(n563), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  NAND2_X1 U621 ( .A1(n558), .A2(n582), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n559), .B(KEYINPUT118), .ZN(n560) );
  XNOR2_X1 U625 ( .A(G162GAT), .B(n560), .ZN(G1347GAT) );
  NAND2_X1 U626 ( .A1(n567), .A2(n574), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(KEYINPUT122), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(n562), .ZN(G1348GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n565) );
  NAND2_X1 U630 ( .A1(n567), .A2(n563), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(G176GAT), .B(n566), .ZN(G1349GAT) );
  XOR2_X1 U633 ( .A(G183GAT), .B(KEYINPUT123), .Z(n569) );
  NAND2_X1 U634 ( .A1(n567), .A2(n582), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G1350GAT) );
  XOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT60), .Z(n576) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n585) );
  NAND2_X1 U639 ( .A1(n585), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(n578) );
  XOR2_X1 U641 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n580) );
  NAND2_X1 U644 ( .A1(n585), .A2(n387), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(n581), .ZN(G1353GAT) );
  XOR2_X1 U647 ( .A(G211GAT), .B(KEYINPUT127), .Z(n584) );
  NAND2_X1 U648 ( .A1(n585), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1354GAT) );
  INV_X1 U650 ( .A(n585), .ZN(n586) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(n588), .Z(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

