//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 1 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n781, new_n782, new_n783, new_n785, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978, new_n979;
  INV_X1    g000(.A(KEYINPUT1), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT69), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT69), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT67), .ZN(new_n207));
  XNOR2_X1  g006(.A(G113gat), .B(G120gat), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G120gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G113gat), .ZN(new_n211));
  INV_X1    g010(.A(G113gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G120gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT67), .ZN(new_n215));
  AND2_X1   g014(.A1(G127gat), .A2(G134gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(G127gat), .A2(G134gat), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT68), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G127gat), .ZN(new_n219));
  INV_X1    g018(.A(G134gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT68), .ZN(new_n222));
  NAND2_X1  g021(.A1(G127gat), .A2(G134gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n209), .A2(new_n215), .A3(new_n218), .A4(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT4), .ZN(new_n226));
  XNOR2_X1  g025(.A(G155gat), .B(G162gat), .ZN(new_n227));
  INV_X1    g026(.A(G148gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G141gat), .ZN(new_n229));
  INV_X1    g028(.A(G141gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G148gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT2), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT77), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT77), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT2), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n227), .B1(new_n232), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G155gat), .ZN(new_n239));
  INV_X1    g038(.A(G162gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n233), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G155gat), .A2(G162gat), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n241), .A2(new_n242), .B1(new_n229), .B2(new_n231), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n221), .B(new_n223), .C1(new_n208), .C2(KEYINPUT1), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n225), .A2(new_n226), .A3(new_n244), .A4(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT81), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n218), .B(new_n224), .C1(new_n207), .C2(new_n208), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n203), .B(new_n205), .C1(new_n214), .C2(KEYINPUT67), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n245), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n242), .ZN(new_n252));
  NOR2_X1   g051(.A1(G155gat), .A2(G162gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G141gat), .B(G148gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT77), .B(KEYINPUT2), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(new_n232), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT4), .B1(new_n251), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n248), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n225), .A2(new_n245), .A3(new_n244), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n263), .A2(new_n247), .A3(KEYINPUT4), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT3), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n257), .A2(new_n265), .A3(new_n259), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT3), .B1(new_n238), .B2(new_n243), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n251), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT78), .ZN(new_n269));
  NOR3_X1   g068(.A1(new_n238), .A2(KEYINPUT3), .A3(new_n243), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n265), .B1(new_n257), .B2(new_n259), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT78), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n272), .A2(new_n273), .A3(new_n251), .ZN(new_n274));
  AOI22_X1  g073(.A1(new_n262), .A2(new_n264), .B1(new_n269), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n276));
  NAND2_X1  g075(.A1(G225gat), .A2(G233gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n251), .A2(new_n260), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n279), .A3(KEYINPUT79), .ZN(new_n280));
  INV_X1    g079(.A(new_n277), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT79), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n251), .A2(new_n282), .A3(new_n260), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n280), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  AND2_X1   g083(.A1(new_n284), .A2(KEYINPUT5), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n261), .A2(new_n246), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n273), .B1(new_n272), .B2(new_n251), .ZN(new_n287));
  AND4_X1   g086(.A1(new_n273), .A2(new_n251), .A3(new_n266), .A4(new_n267), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n286), .B(new_n277), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT80), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  AND4_X1   g089(.A1(KEYINPUT80), .A2(new_n289), .A3(KEYINPUT5), .A4(new_n284), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n278), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G1gat), .B(G29gat), .ZN(new_n293));
  INV_X1    g092(.A(G85gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT0), .B(G57gat), .ZN(new_n296));
  XOR2_X1   g095(.A(new_n295), .B(new_n296), .Z(new_n297));
  NAND2_X1  g096(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT82), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n299), .A2(KEYINPUT6), .ZN(new_n300));
  INV_X1    g099(.A(new_n297), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n301), .B(new_n278), .C1(new_n290), .C2(new_n291), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n298), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n292), .B(new_n297), .C1(new_n299), .C2(KEYINPUT6), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G227gat), .A2(G233gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT70), .ZN(new_n308));
  INV_X1    g107(.A(G190gat), .ZN(new_n309));
  INV_X1    g108(.A(G183gat), .ZN(new_n310));
  OAI211_X1 g109(.A(KEYINPUT65), .B(new_n309), .C1(new_n310), .C2(KEYINPUT27), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT28), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT27), .ZN(new_n314));
  AOI21_X1  g113(.A(G190gat), .B1(new_n314), .B2(G183gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n310), .A2(KEYINPUT27), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n311), .A2(new_n315), .A3(new_n312), .A4(new_n316), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G183gat), .A2(G190gat), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(G169gat), .A2(G176gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NOR3_X1   g123(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n325));
  OAI211_X1 g124(.A(KEYINPUT66), .B(new_n321), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT26), .ZN(new_n328));
  INV_X1    g127(.A(G169gat), .ZN(new_n329));
  INV_X1    g128(.A(G176gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n331), .A2(new_n323), .A3(new_n322), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT66), .B1(new_n332), .B2(new_n321), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n320), .A2(new_n327), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n335), .B1(G183gat), .B2(G190gat), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n329), .A2(new_n330), .A3(KEYINPUT23), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n340), .B1(G169gat), .B2(G176gat), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n339), .A2(new_n341), .A3(KEYINPUT25), .A4(new_n323), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  AND3_X1   g142(.A1(new_n339), .A2(new_n341), .A3(new_n323), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT64), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT24), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n321), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n310), .A2(new_n309), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n335), .A3(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n337), .A2(new_n345), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n344), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT25), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n343), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n334), .A2(new_n353), .ZN(new_n354));
  AOI211_X1 g153(.A(new_n217), .B(new_n216), .C1(new_n214), .C2(new_n202), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n218), .A2(new_n224), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n208), .A2(new_n207), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n355), .B1(new_n358), .B2(new_n209), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n308), .B1(new_n354), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n251), .B1(new_n334), .B2(new_n353), .ZN(new_n361));
  OR2_X1    g160(.A1(new_n338), .A2(new_n342), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n339), .A2(new_n341), .A3(new_n323), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n347), .A2(new_n335), .A3(new_n348), .ZN(new_n364));
  INV_X1    g163(.A(new_n350), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n362), .B1(new_n366), .B2(KEYINPUT25), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n321), .B1(new_n324), .B2(new_n325), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT66), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n370), .A2(new_n326), .A3(new_n318), .A4(new_n319), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n367), .A2(new_n359), .A3(new_n308), .A4(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n361), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n307), .B1(new_n360), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT33), .ZN(new_n375));
  XNOR2_X1  g174(.A(G15gat), .B(G43gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(G71gat), .B(G99gat), .ZN(new_n377));
  XOR2_X1   g176(.A(new_n376), .B(new_n377), .Z(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n374), .B(KEYINPUT32), .C1(new_n375), .C2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n379), .B1(new_n374), .B2(KEYINPUT32), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT71), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n374), .A2(new_n375), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n382), .B1(new_n381), .B2(new_n383), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n380), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n360), .A2(new_n373), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n306), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n388), .B(KEYINPUT34), .Z(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n389), .B(new_n380), .C1(new_n385), .C2(new_n384), .ZN(new_n392));
  XNOR2_X1  g191(.A(G8gat), .B(G36gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(G64gat), .B(G92gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G211gat), .B(G218gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  AND2_X1   g196(.A1(G197gat), .A2(G204gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(G197gat), .A2(G204gat), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OR2_X1    g199(.A1(KEYINPUT74), .A2(G218gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(KEYINPUT74), .A2(G218gat), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(G211gat), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT22), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n400), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT75), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n397), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(KEYINPUT74), .A2(G218gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(KEYINPUT74), .A2(G218gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT22), .B1(new_n410), .B2(G211gat), .ZN(new_n411));
  OAI211_X1 g210(.A(KEYINPUT75), .B(new_n396), .C1(new_n411), .C2(new_n400), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT76), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n367), .A2(new_n371), .ZN(new_n416));
  INV_X1    g215(.A(G226gat), .ZN(new_n417));
  INV_X1    g216(.A(G233gat), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT29), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n419), .B1(new_n416), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n415), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  OAI22_X1  g223(.A1(new_n354), .A2(KEYINPUT29), .B1(new_n417), .B2(new_n418), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT76), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n414), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n421), .A2(new_n423), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n414), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n395), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n395), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n423), .A2(new_n415), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n425), .A2(new_n420), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n433), .B1(new_n434), .B2(new_n415), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n429), .B(new_n432), .C1(new_n435), .C2(new_n414), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n431), .A2(new_n436), .A3(KEYINPUT30), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n427), .A2(new_n430), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT30), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(new_n439), .A3(new_n432), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n305), .A2(new_n391), .A3(new_n392), .A4(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(G22gat), .ZN(new_n443));
  INV_X1    g242(.A(G228gat), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n444), .A2(new_n418), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n405), .A2(new_n397), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n422), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n405), .A2(new_n397), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n265), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n260), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n266), .A2(new_n422), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n413), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n445), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT84), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n407), .A2(new_n412), .B1(new_n266), .B2(new_n422), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT83), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n445), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n413), .A2(new_n457), .A3(new_n451), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n265), .B1(new_n413), .B2(KEYINPUT29), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n260), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n455), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n445), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n464), .B1(new_n452), .B2(KEYINPUT83), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n456), .A2(new_n457), .ZN(new_n466));
  AND4_X1   g265(.A1(new_n455), .A2(new_n462), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n443), .B(new_n454), .C1(new_n463), .C2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT86), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n454), .B1(new_n463), .B2(new_n467), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(G22gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n471), .A2(new_n469), .A3(G22gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(G78gat), .B(G106gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(KEYINPUT31), .B(G50gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n475), .B(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n473), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n477), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n452), .A2(KEYINPUT83), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n480), .A2(new_n466), .A3(new_n445), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n461), .A2(new_n260), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT84), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n462), .A2(new_n465), .A3(new_n455), .A4(new_n466), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n443), .B1(new_n485), .B2(new_n454), .ZN(new_n486));
  AOI211_X1 g285(.A(G22gat), .B(new_n453), .C1(new_n483), .C2(new_n484), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n479), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT85), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT85), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n490), .B(new_n479), .C1(new_n486), .C2(new_n487), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n478), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT35), .B1(new_n442), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT92), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n489), .A2(new_n491), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT35), .B1(new_n496), .B2(new_n478), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT73), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n498), .B1(new_n386), .B2(new_n390), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n391), .A2(new_n392), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n499), .B1(new_n500), .B2(new_n498), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n292), .A2(KEYINPUT6), .A3(new_n297), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT6), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n298), .A2(new_n503), .A3(new_n302), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n502), .B1(new_n504), .B2(KEYINPUT90), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT90), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n298), .A2(new_n506), .A3(new_n503), .A4(new_n302), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n437), .A2(KEYINPUT87), .A3(new_n440), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT87), .B1(new_n437), .B2(new_n440), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n497), .A2(new_n501), .A3(new_n508), .A4(new_n511), .ZN(new_n512));
  OAI211_X1 g311(.A(KEYINPUT92), .B(KEYINPUT35), .C1(new_n442), .C2(new_n492), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n495), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT36), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT72), .B1(new_n500), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT72), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n391), .A2(new_n392), .A3(new_n517), .A4(KEYINPUT36), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n516), .B(new_n518), .C1(new_n501), .C2(KEYINPUT36), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n424), .A2(new_n426), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n414), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT37), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n522), .B1(new_n428), .B2(new_n413), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT38), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n522), .B(new_n429), .C1(new_n435), .C2(new_n414), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(new_n395), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT91), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT91), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n524), .A2(new_n528), .A3(new_n395), .A4(new_n525), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT37), .B1(new_n427), .B2(new_n430), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n531), .A2(new_n395), .A3(new_n525), .ZN(new_n532));
  AOI22_X1  g331(.A1(new_n532), .A2(KEYINPUT38), .B1(new_n438), .B2(new_n432), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n505), .A2(new_n530), .A3(new_n533), .A4(new_n507), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n262), .A2(new_n264), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n287), .A2(new_n288), .ZN(new_n536));
  OAI211_X1 g335(.A(KEYINPUT88), .B(new_n281), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT88), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n538), .B1(new_n275), .B2(new_n277), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT39), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n280), .A2(new_n283), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n541), .B1(new_n543), .B2(new_n277), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n544), .A2(KEYINPUT89), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(KEYINPUT89), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n545), .A2(new_n537), .A3(new_n539), .A4(new_n546), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n542), .A2(new_n547), .A3(KEYINPUT40), .A4(new_n301), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n548), .A2(new_n298), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n542), .A2(new_n301), .A3(new_n547), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT40), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n549), .B(new_n552), .C1(new_n509), .C2(new_n510), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n492), .B1(new_n534), .B2(new_n553), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n492), .A2(new_n305), .A3(new_n441), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n519), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n514), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NOR3_X1   g358(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n560));
  INV_X1    g359(.A(G29gat), .ZN(new_n561));
  INV_X1    g360(.A(G36gat), .ZN(new_n562));
  OAI22_X1  g361(.A1(new_n559), .A2(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(G43gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(G50gat), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT15), .B1(new_n565), .B2(KEYINPUT93), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G43gat), .B(G50gat), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT15), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n563), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n567), .A2(new_n569), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n574), .A2(KEYINPUT17), .ZN(new_n575));
  XNOR2_X1  g374(.A(G15gat), .B(G22gat), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT16), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n576), .B1(new_n577), .B2(G1gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n578), .B(new_n579), .C1(G1gat), .C2(new_n576), .ZN(new_n580));
  NOR2_X1   g379(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n574), .A2(KEYINPUT17), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n575), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G229gat), .A2(G233gat), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n574), .A2(new_n582), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT18), .ZN(new_n588));
  OR2_X1    g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n588), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT95), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n591), .B1(new_n574), .B2(new_n582), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n586), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n585), .B(KEYINPUT13), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n586), .A2(new_n592), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n593), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n589), .A2(new_n590), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G113gat), .B(G141gat), .ZN(new_n599));
  INV_X1    g398(.A(G197gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT11), .B(G169gat), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n601), .B(new_n602), .Z(new_n603));
  XOR2_X1   g402(.A(new_n603), .B(KEYINPUT12), .Z(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n598), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n589), .A2(new_n590), .A3(new_n597), .A4(new_n604), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n607), .A2(KEYINPUT96), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(KEYINPUT96), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n606), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G71gat), .B(G78gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT98), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(G57gat), .B(G64gat), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT97), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n613), .B(new_n617), .C1(new_n616), .C2(new_n615), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT99), .ZN(new_n619));
  INV_X1    g418(.A(new_n612), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT9), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n620), .B1(new_n621), .B2(new_n615), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G85gat), .A2(G92gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT7), .ZN(new_n626));
  INV_X1    g425(.A(G99gat), .ZN(new_n627));
  INV_X1    g426(.A(G106gat), .ZN(new_n628));
  OAI21_X1  g427(.A(KEYINPUT8), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n626), .B(new_n629), .C1(G85gat), .C2(G92gat), .ZN(new_n630));
  XOR2_X1   g429(.A(G99gat), .B(G106gat), .Z(new_n631));
  XOR2_X1   g430(.A(new_n630), .B(new_n631), .Z(new_n632));
  NAND2_X1  g431(.A1(new_n624), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT10), .ZN(new_n634));
  INV_X1    g433(.A(new_n632), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n623), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n624), .A2(KEYINPUT10), .A3(new_n632), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G230gat), .A2(G233gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT102), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G120gat), .B(G148gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(G176gat), .B(G204gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n642), .B1(new_n633), .B2(new_n636), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n646), .B1(new_n647), .B2(KEYINPUT103), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n643), .B(new_n648), .C1(KEYINPUT103), .C2(new_n647), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n646), .B(KEYINPUT104), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n641), .B1(new_n637), .B2(new_n638), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n650), .B1(new_n651), .B2(new_n647), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n611), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n635), .A2(new_n574), .ZN(new_n655));
  NAND2_X1  g454(.A1(G232gat), .A2(G233gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT100), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n655), .B1(KEYINPUT41), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n575), .A2(new_n583), .A3(new_n635), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(G190gat), .B(G218gat), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n658), .A2(KEYINPUT41), .ZN(new_n664));
  XOR2_X1   g463(.A(G134gat), .B(G162gat), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n659), .A2(new_n662), .A3(new_n660), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n666), .B1(new_n667), .B2(KEYINPUT101), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n663), .B(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT21), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n623), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g471(.A(G127gat), .B(G155gat), .Z(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(G231gat), .A2(G233gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(new_n310), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G211gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n674), .B(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n582), .B1(new_n623), .B2(new_n671), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n678), .A2(new_n682), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n557), .A2(new_n654), .A3(new_n670), .A4(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n305), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g494(.A1(new_n691), .A2(new_n511), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT16), .B(G8gat), .Z(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT42), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n696), .A2(KEYINPUT42), .A3(new_n697), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n702));
  INV_X1    g501(.A(G8gat), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n702), .B1(new_n696), .B2(new_n703), .ZN(new_n704));
  OAI211_X1 g503(.A(KEYINPUT106), .B(G8gat), .C1(new_n691), .C2(new_n511), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n700), .A2(new_n701), .A3(new_n704), .A4(new_n705), .ZN(G1325gat));
  INV_X1    g505(.A(new_n519), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n692), .A2(G15gat), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(G15gat), .B1(new_n692), .B2(new_n501), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(G1326gat));
  INV_X1    g509(.A(new_n492), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n691), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g511(.A(KEYINPUT43), .B(G22gat), .Z(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1327gat));
  NAND2_X1  g513(.A1(new_n557), .A2(new_n669), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n654), .A2(new_n685), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n717), .A2(new_n561), .A3(new_n693), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT45), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n720), .B1(new_n557), .B2(new_n669), .ZN(new_n721));
  AOI211_X1 g520(.A(KEYINPUT44), .B(new_n670), .C1(new_n514), .C2(new_n556), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n723), .A2(new_n716), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n693), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n725), .A2(KEYINPUT107), .ZN(new_n726));
  OAI21_X1  g525(.A(G29gat), .B1(new_n725), .B2(KEYINPUT107), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n719), .B1(new_n726), .B2(new_n727), .ZN(G1328gat));
  INV_X1    g527(.A(new_n511), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n717), .A2(new_n562), .A3(new_n729), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n730), .B(KEYINPUT46), .Z(new_n731));
  NAND2_X1  g530(.A1(new_n724), .A2(new_n729), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n731), .B1(new_n733), .B2(new_n562), .ZN(G1329gat));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n736));
  INV_X1    g535(.A(new_n716), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n707), .B(new_n737), .C1(new_n721), .C2(new_n722), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n736), .B1(new_n738), .B2(G43gat), .ZN(new_n739));
  INV_X1    g538(.A(new_n501), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(G43gat), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n717), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT47), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n738), .A2(new_n736), .A3(G43gat), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n742), .ZN(new_n749));
  INV_X1    g548(.A(new_n738), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n564), .B1(new_n750), .B2(KEYINPUT109), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n738), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n749), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n735), .B(new_n748), .C1(new_n754), .C2(new_n743), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n715), .A2(KEYINPUT44), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n670), .B1(new_n514), .B2(new_n556), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n720), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n759), .A2(KEYINPUT109), .A3(new_n707), .A4(new_n737), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(new_n753), .A3(G43gat), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n743), .B1(new_n761), .B2(new_n742), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n746), .A2(new_n739), .A3(new_n744), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT110), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n755), .A2(new_n764), .ZN(G1330gat));
  NAND2_X1  g564(.A1(new_n724), .A2(new_n492), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n711), .A2(G50gat), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n766), .A2(G50gat), .B1(new_n717), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g568(.A1(new_n685), .A2(new_n610), .A3(new_n669), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n557), .A2(new_n653), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT111), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n693), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g574(.A1(new_n772), .A2(new_n511), .ZN(new_n776));
  NOR2_X1   g575(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n777));
  AND2_X1   g576(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(new_n776), .B2(new_n777), .ZN(G1333gat));
  NAND3_X1  g579(.A1(new_n773), .A2(G71gat), .A3(new_n707), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n772), .A2(new_n740), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n781), .B1(new_n782), .B2(G71gat), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g583(.A1(new_n772), .A2(new_n711), .ZN(new_n785));
  XNOR2_X1  g584(.A(KEYINPUT112), .B(G78gat), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(G1335gat));
  INV_X1    g586(.A(new_n653), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n611), .A2(new_n685), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(KEYINPUT113), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n757), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n788), .B1(new_n791), .B2(KEYINPUT51), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n757), .A2(new_n793), .A3(new_n790), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(G85gat), .B1(new_n795), .B2(new_n693), .ZN(new_n796));
  INV_X1    g595(.A(new_n790), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(new_n788), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n759), .A2(KEYINPUT114), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT114), .B1(new_n759), .B2(new_n798), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n305), .A2(new_n294), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n796), .B1(new_n802), .B2(new_n803), .ZN(G1336gat));
  NOR2_X1   g603(.A1(new_n511), .A2(G92gat), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n792), .A2(new_n794), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT115), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n792), .A2(new_n808), .A3(new_n794), .A4(new_n805), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n729), .B1(new_n800), .B2(new_n801), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n810), .B1(new_n811), .B2(G92gat), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813));
  INV_X1    g612(.A(G92gat), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n723), .A2(new_n788), .A3(new_n797), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n814), .B1(new_n815), .B2(new_n729), .ZN(new_n816));
  XNOR2_X1  g615(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n806), .A2(new_n817), .ZN(new_n818));
  OAI22_X1  g617(.A1(new_n812), .A2(new_n813), .B1(new_n816), .B2(new_n818), .ZN(G1337gat));
  AOI21_X1  g618(.A(G99gat), .B1(new_n795), .B2(new_n501), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n519), .A2(new_n627), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n820), .B1(new_n802), .B2(new_n821), .ZN(G1338gat));
  OAI21_X1  g621(.A(new_n492), .B1(new_n800), .B2(new_n801), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n711), .A2(G106gat), .ZN(new_n824));
  AOI22_X1  g623(.A1(new_n823), .A2(G106gat), .B1(new_n795), .B2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n628), .B1(new_n815), .B2(new_n492), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n795), .A2(new_n824), .ZN(new_n828));
  XNOR2_X1  g627(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI22_X1  g629(.A1(new_n825), .A2(new_n826), .B1(new_n827), .B2(new_n830), .ZN(G1339gat));
  NAND3_X1  g630(.A1(new_n637), .A2(new_n641), .A3(new_n638), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n643), .A2(new_n832), .A3(KEYINPUT54), .ZN(new_n833));
  INV_X1    g632(.A(new_n646), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n834), .B1(new_n651), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n833), .A2(KEYINPUT55), .A3(new_n836), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n837), .A2(new_n649), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n833), .A2(new_n836), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n838), .A2(new_n610), .A3(new_n841), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n607), .B(KEYINPUT96), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n595), .B1(new_n593), .B2(new_n596), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n585), .B1(new_n584), .B2(new_n586), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n844), .B1(KEYINPUT118), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n846), .B1(KEYINPUT118), .B2(new_n845), .ZN(new_n847));
  INV_X1    g646(.A(new_n603), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n843), .A2(new_n653), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n669), .B1(new_n842), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n838), .A2(new_n669), .A3(new_n841), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n843), .A2(new_n849), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n685), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n770), .A2(new_n788), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n857), .A2(new_n500), .A3(new_n492), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n858), .A2(new_n693), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n859), .A2(new_n511), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n212), .A3(new_n610), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n857), .A2(new_n740), .A3(new_n492), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(new_n693), .A3(new_n511), .ZN(new_n863));
  OAI21_X1  g662(.A(G113gat), .B1(new_n863), .B2(new_n611), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n861), .A2(new_n864), .ZN(G1340gat));
  NAND3_X1  g664(.A1(new_n860), .A2(new_n210), .A3(new_n653), .ZN(new_n866));
  OAI21_X1  g665(.A(G120gat), .B1(new_n863), .B2(new_n788), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT119), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n867), .A2(new_n868), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(G1341gat));
  NOR3_X1   g670(.A1(new_n863), .A2(new_n219), .A3(new_n685), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n860), .A2(new_n686), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(new_n219), .ZN(G1342gat));
  NOR2_X1   g673(.A1(new_n729), .A2(new_n670), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n859), .A2(new_n220), .A3(new_n875), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n876), .A2(KEYINPUT56), .ZN(new_n877));
  OAI21_X1  g676(.A(G134gat), .B1(new_n863), .B2(new_n670), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(KEYINPUT56), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(G1343gat));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n841), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n839), .A2(KEYINPUT120), .A3(new_n840), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n882), .A2(new_n838), .A3(new_n610), .A4(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n669), .B1(new_n884), .B2(new_n850), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n685), .B1(new_n885), .B2(new_n854), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n886), .A2(new_n856), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT57), .B1(new_n887), .B2(new_n711), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n707), .A2(new_n305), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n511), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n711), .B1(new_n855), .B2(new_n856), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n888), .A2(new_n610), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n230), .B1(new_n894), .B2(KEYINPUT122), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n895), .B1(KEYINPUT122), .B2(new_n894), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n891), .A2(new_n889), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n511), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n898), .A2(G141gat), .A3(new_n611), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(KEYINPUT58), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n894), .A2(KEYINPUT121), .A3(G141gat), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT121), .B1(new_n894), .B2(G141gat), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n902), .A2(new_n903), .A3(new_n899), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT58), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n901), .B1(new_n904), .B2(new_n905), .ZN(G1344gat));
  INV_X1    g705(.A(new_n898), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n228), .A3(new_n653), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n888), .A2(new_n893), .ZN(new_n909));
  AOI211_X1 g708(.A(KEYINPUT59), .B(new_n228), .C1(new_n909), .C2(new_n653), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n891), .A2(KEYINPUT57), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n711), .B1(new_n886), .B2(new_n856), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n912), .B1(new_n913), .B2(KEYINPUT57), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n914), .A2(new_n511), .A3(new_n653), .A4(new_n889), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n911), .B1(new_n915), .B2(G148gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n908), .B1(new_n910), .B2(new_n916), .ZN(G1345gat));
  AOI21_X1  g716(.A(G155gat), .B1(new_n907), .B2(new_n686), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n685), .A2(new_n239), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n909), .B2(new_n919), .ZN(G1346gat));
  NAND3_X1  g719(.A1(new_n897), .A2(new_n240), .A3(new_n875), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n909), .A2(new_n669), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n922), .B2(new_n240), .ZN(G1347gat));
  NOR2_X1   g722(.A1(new_n511), .A2(new_n693), .ZN(new_n924));
  XOR2_X1   g723(.A(new_n924), .B(KEYINPUT123), .Z(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n862), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(G169gat), .B1(new_n927), .B2(new_n611), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n858), .A2(new_n924), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n610), .A2(new_n329), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(G1348gat));
  NOR3_X1   g730(.A1(new_n927), .A2(new_n330), .A3(new_n788), .ZN(new_n932));
  INV_X1    g731(.A(new_n929), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(new_n653), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n932), .B1(new_n330), .B2(new_n934), .ZN(G1349gat));
  OAI21_X1  g734(.A(G183gat), .B1(new_n927), .B2(new_n685), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n314), .A2(G183gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n686), .A2(new_n937), .A3(new_n316), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n936), .B1(new_n929), .B2(new_n938), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g739(.A1(new_n862), .A2(new_n669), .A3(new_n926), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G190gat), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT124), .ZN(new_n943));
  OR3_X1    g742(.A1(new_n942), .A2(new_n943), .A3(KEYINPUT61), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n942), .B2(KEYINPUT61), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n942), .A2(KEYINPUT61), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n933), .A2(new_n309), .A3(new_n669), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(G1351gat));
  NAND2_X1  g748(.A1(new_n926), .A2(new_n519), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT126), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n950), .A2(KEYINPUT126), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n914), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(G197gat), .B1(new_n953), .B2(new_n611), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n857), .A2(new_n693), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n519), .A2(new_n729), .A3(new_n492), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n956), .A2(KEYINPUT125), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(KEYINPUT125), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n955), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n960), .A2(new_n600), .A3(new_n610), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n954), .A2(new_n961), .ZN(G1352gat));
  NOR3_X1   g761(.A1(new_n959), .A2(G204gat), .A3(new_n788), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT62), .ZN(new_n964));
  OAI21_X1  g763(.A(G204gat), .B1(new_n953), .B2(new_n788), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1353gat));
  INV_X1    g765(.A(G211gat), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n950), .A2(new_n685), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n967), .B1(new_n914), .B2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n970));
  OR3_X1    g769(.A1(new_n969), .A2(new_n970), .A3(KEYINPUT63), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n970), .B1(new_n969), .B2(KEYINPUT63), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n969), .A2(KEYINPUT63), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n960), .A2(new_n967), .A3(new_n686), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(G1354gat));
  AOI21_X1  g775(.A(G218gat), .B1(new_n960), .B2(new_n669), .ZN(new_n977));
  INV_X1    g776(.A(new_n953), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n669), .A2(new_n410), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(G1355gat));
endmodule


