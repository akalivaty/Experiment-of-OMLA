//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 0 1 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n547, new_n548, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n457));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  AOI21_X1  g035(.A(G2105), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G137), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND3_X1   g038(.A1(new_n463), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT66), .B1(new_n463), .B2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G101), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(G125), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n463), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n467), .A2(new_n472), .ZN(G160));
  NOR2_X1   g048(.A1(new_n468), .A2(new_n469), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(new_n463), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  OAI21_X1  g051(.A(KEYINPUT67), .B1(G100), .B2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NOR3_X1   g053(.A1(KEYINPUT67), .A2(G100), .A3(G2105), .ZN(new_n479));
  OAI221_X1 g054(.A(G2104), .B1(G112), .B2(new_n463), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n461), .A2(G136), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n476), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  OAI211_X1 g058(.A(G138), .B(new_n463), .C1(new_n468), .C2(new_n469), .ZN(new_n484));
  NAND2_X1  g059(.A1(KEYINPUT68), .A2(KEYINPUT4), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(G126), .A2(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n463), .A2(G138), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(new_n485), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n459), .A2(new_n460), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OR2_X1    g066(.A1(new_n463), .A2(G114), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n486), .A2(new_n491), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT69), .B1(new_n498), .B2(G651), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n500));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT6), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n498), .A2(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G50), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(new_n506), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n505), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G88), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n510), .A2(new_n511), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n516), .A2(new_n501), .ZN(new_n517));
  AND3_X1   g092(.A1(new_n508), .A2(new_n514), .A3(new_n517), .ZN(G166));
  AND2_X1   g093(.A1(new_n503), .A2(new_n504), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n519), .A2(G89), .A3(new_n515), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(G51), .A3(G543), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n522), .A2(KEYINPUT7), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(KEYINPUT7), .ZN(new_n524));
  AND2_X1   g099(.A1(G63), .A2(G651), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n523), .A2(new_n524), .B1(new_n515), .B2(new_n525), .ZN(new_n526));
  AND3_X1   g101(.A1(new_n520), .A2(new_n521), .A3(new_n526), .ZN(G168));
  NAND3_X1  g102(.A1(new_n519), .A2(G90), .A3(new_n515), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n519), .A2(G52), .A3(G543), .ZN(new_n529));
  NAND2_X1  g104(.A1(G77), .A2(G543), .ZN(new_n530));
  INV_X1    g105(.A(G64), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n512), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G651), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n528), .A2(new_n529), .A3(new_n533), .ZN(G171));
  AOI22_X1  g109(.A1(G43), .A2(new_n507), .B1(new_n513), .B2(G81), .ZN(new_n535));
  NAND2_X1  g110(.A1(G68), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G56), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n512), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT70), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g115(.A(KEYINPUT70), .B(new_n536), .C1(new_n512), .C2(new_n537), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n540), .A2(G651), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n535), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  NAND4_X1  g120(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  NAND4_X1  g124(.A1(new_n503), .A2(G53), .A3(G543), .A4(new_n504), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT9), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(KEYINPUT71), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n550), .B(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(G78), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G65), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n512), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n513), .A2(G91), .B1(new_n556), .B2(G651), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n553), .A2(new_n557), .ZN(G299));
  NAND3_X1  g133(.A1(new_n528), .A2(new_n529), .A3(new_n533), .ZN(G301));
  NAND3_X1  g134(.A1(new_n520), .A2(new_n521), .A3(new_n526), .ZN(G286));
  NAND3_X1  g135(.A1(new_n508), .A2(new_n514), .A3(new_n517), .ZN(G303));
  INV_X1    g136(.A(G49), .ZN(new_n562));
  NOR4_X1   g137(.A1(new_n505), .A2(KEYINPUT72), .A3(new_n562), .A4(new_n506), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT72), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n562), .A2(new_n506), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n564), .B1(new_n519), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n515), .A2(G74), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G651), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n519), .A2(new_n515), .ZN(new_n570));
  INV_X1    g145(.A(G87), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G288));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n512), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G651), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n503), .A2(G48), .A3(G543), .A4(new_n504), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n503), .A2(G86), .A3(new_n504), .A4(new_n515), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(KEYINPUT73), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT73), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n578), .A2(new_n583), .A3(new_n579), .A4(new_n580), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n582), .A2(new_n584), .ZN(G305));
  NAND3_X1  g160(.A1(new_n519), .A2(G85), .A3(new_n515), .ZN(new_n586));
  NAND2_X1  g161(.A1(G72), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G60), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n512), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G651), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n503), .A2(G47), .A3(G543), .A4(new_n504), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n586), .A2(new_n590), .A3(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  XNOR2_X1  g168(.A(KEYINPUT74), .B(KEYINPUT10), .ZN(new_n594));
  XOR2_X1   g169(.A(new_n594), .B(KEYINPUT75), .Z(new_n595));
  INV_X1    g170(.A(G92), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n570), .B2(new_n596), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n594), .B(KEYINPUT75), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n513), .A2(new_n598), .A3(G92), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n512), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n507), .A2(G54), .B1(new_n602), .B2(G651), .ZN(new_n603));
  AND3_X1   g178(.A1(new_n597), .A2(new_n599), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n593), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n593), .B1(new_n604), .B2(G868), .ZN(G321));
  NAND2_X1  g181(.A1(G286), .A2(G868), .ZN(new_n607));
  INV_X1    g182(.A(G299), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G297));
  OAI21_X1  g184(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND3_X1  g187(.A1(new_n597), .A2(new_n603), .A3(new_n599), .ZN(new_n613));
  OAI21_X1  g188(.A(G868), .B1(new_n613), .B2(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G868), .B2(new_n544), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g191(.A1(new_n464), .A2(new_n465), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(new_n490), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT76), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT13), .Z(new_n621));
  INV_X1    g196(.A(G2100), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n475), .A2(G123), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  INV_X1    g201(.A(G111), .ZN(new_n627));
  AOI22_X1  g202(.A1(new_n626), .A2(KEYINPUT77), .B1(new_n627), .B2(G2105), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(KEYINPUT77), .B2(new_n626), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n461), .A2(G135), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n625), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G2096), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n623), .A2(new_n624), .A3(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2427), .B(G2430), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(KEYINPUT14), .ZN(new_n639));
  AND2_X1   g214(.A1(new_n639), .A2(KEYINPUT78), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n639), .A2(KEYINPUT78), .ZN(new_n641));
  OAI22_X1  g216(.A1(new_n640), .A2(new_n641), .B1(new_n636), .B2(new_n637), .ZN(new_n642));
  XOR2_X1   g217(.A(G2451), .B(G2454), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n642), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT79), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G1341), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G1348), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(G14), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n645), .A2(new_n649), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(G401));
  INV_X1    g228(.A(KEYINPUT18), .ZN(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(KEYINPUT17), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n655), .A2(new_n656), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n654), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(new_n622), .ZN(new_n661));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(new_n657), .B2(KEYINPUT18), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(new_n632), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n661), .B(new_n664), .ZN(G227));
  XNOR2_X1  g240(.A(G1981), .B(G1986), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT19), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1956), .B(G2474), .Z(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  AND2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT20), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n671), .A2(new_n672), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n670), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT80), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  OR3_X1    g254(.A1(new_n670), .A2(new_n673), .A3(new_n676), .ZN(new_n680));
  AND3_X1   g255(.A1(new_n675), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1991), .B(G1996), .Z(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n667), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n683), .A2(new_n684), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n683), .A2(new_n684), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n688), .A2(new_n666), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(G229));
  AOI22_X1  g267(.A1(new_n617), .A2(G105), .B1(G141), .B2(new_n461), .ZN(new_n693));
  NAND3_X1  g268(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT26), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(G129), .B2(new_n475), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n699), .B2(G32), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT27), .B(G1996), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  INV_X1    g279(.A(G34), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(KEYINPUT24), .ZN(new_n706));
  AOI21_X1  g281(.A(G29), .B1(new_n705), .B2(KEYINPUT24), .ZN(new_n707));
  AOI22_X1  g282(.A1(G160), .A2(G29), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n704), .B1(G2084), .B2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G1961), .ZN(new_n710));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  NOR2_X1   g286(.A1(G171), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G5), .B2(new_n711), .ZN(new_n713));
  AOI211_X1 g288(.A(new_n703), .B(new_n709), .C1(new_n710), .C2(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(G29), .A2(G35), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G162), .B2(G29), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT29), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(G2090), .Z(new_n718));
  AND2_X1   g293(.A1(new_n699), .A2(G33), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT25), .ZN(new_n720));
  NAND2_X1  g295(.A1(G103), .A2(G2104), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(G2105), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n463), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n461), .A2(G139), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n490), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n463), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n719), .B1(new_n726), .B2(G29), .ZN(new_n727));
  INV_X1    g302(.A(G2072), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(G164), .A2(new_n699), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G27), .B2(new_n699), .ZN(new_n731));
  INV_X1    g306(.A(G2078), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n727), .A2(new_n728), .ZN(new_n735));
  AND4_X1   g310(.A1(new_n729), .A2(new_n733), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n708), .A2(G2084), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT88), .Z(new_n738));
  NAND4_X1  g313(.A1(new_n714), .A2(new_n718), .A3(new_n736), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT91), .B(KEYINPUT23), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n711), .A2(G20), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G299), .B2(G16), .ZN(new_n743));
  INV_X1    g318(.A(G1956), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT31), .B(G11), .Z(new_n746));
  INV_X1    g321(.A(KEYINPUT30), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n699), .B1(new_n747), .B2(G28), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n749), .A2(KEYINPUT89), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n749), .A2(KEYINPUT89), .B1(new_n747), .B2(G28), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n746), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n631), .B2(new_n699), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n711), .A2(G21), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G168), .B2(new_n711), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n753), .B1(new_n755), .B2(G1966), .ZN(new_n756));
  OAI221_X1 g331(.A(new_n756), .B1(G1966), .B2(new_n755), .C1(new_n713), .C2(new_n710), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT90), .ZN(new_n758));
  NOR3_X1   g333(.A1(new_n739), .A2(new_n745), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n475), .A2(G128), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n461), .A2(G140), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n463), .A2(G116), .ZN(new_n762));
  OAI21_X1  g337(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n760), .B(new_n761), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G29), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n699), .A2(G26), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT28), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G2067), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n604), .A2(G16), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G4), .B2(G16), .ZN(new_n772));
  INV_X1    g347(.A(G1348), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n773), .B2(new_n772), .ZN(new_n775));
  NOR2_X1   g350(.A1(G16), .A2(G19), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n544), .B2(G16), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT86), .Z(new_n778));
  AND2_X1   g353(.A1(new_n778), .A2(G1341), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n778), .A2(G1341), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n775), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT87), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n759), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n711), .A2(G23), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n573), .B2(new_n711), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT84), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT33), .B(G1976), .Z(new_n789));
  OR2_X1    g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT32), .B(G1981), .ZN(new_n791));
  MUX2_X1   g366(.A(G6), .B(G305), .S(G16), .Z(new_n792));
  AOI22_X1  g367(.A1(new_n788), .A2(new_n789), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n711), .A2(G22), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G166), .B2(new_n711), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(G1971), .Z(new_n796));
  OR2_X1    g371(.A1(new_n792), .A2(new_n791), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n790), .A2(new_n793), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n798), .A2(KEYINPUT34), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(KEYINPUT34), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n475), .A2(G119), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n461), .A2(G131), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n463), .A2(G107), .ZN(new_n803));
  OAI21_X1  g378(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n801), .B(new_n802), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(G29), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n699), .A2(G25), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT81), .Z(new_n808));
  NAND2_X1  g383(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT35), .B(G1991), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT82), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n809), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n711), .A2(G24), .ZN(new_n813));
  AND3_X1   g388(.A1(new_n586), .A2(new_n590), .A3(new_n591), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(new_n711), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT83), .Z(new_n816));
  OAI21_X1  g391(.A(new_n812), .B1(new_n816), .B2(G1986), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(G1986), .B2(new_n816), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n799), .A2(new_n800), .A3(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT85), .B(KEYINPUT36), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n819), .A2(new_n821), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n785), .B1(new_n822), .B2(new_n823), .ZN(G311));
  INV_X1    g399(.A(G311), .ZN(G150));
  NAND2_X1  g400(.A1(G80), .A2(G543), .ZN(new_n826));
  INV_X1    g401(.A(G67), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n512), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(G651), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n503), .A2(G93), .A3(new_n504), .A4(new_n515), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n503), .A2(G55), .A3(G543), .A4(new_n504), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(KEYINPUT92), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT92), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n829), .A2(new_n834), .A3(new_n830), .A4(new_n831), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n543), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n832), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n837), .A2(new_n535), .A3(new_n834), .A4(new_n542), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT38), .Z(new_n840));
  NAND2_X1  g415(.A1(new_n604), .A2(G559), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT93), .B(G860), .Z(new_n845));
  NAND3_X1  g420(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n837), .A2(new_n845), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT37), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(G145));
  XNOR2_X1  g424(.A(new_n620), .B(new_n805), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n697), .B(new_n726), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n764), .B(G164), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n475), .A2(G130), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n461), .A2(G142), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n463), .A2(G118), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n854), .B(new_n855), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n853), .B(new_n858), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n852), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n852), .A2(new_n859), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(G160), .B(new_n482), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(new_n631), .Z(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(G37), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n860), .A2(new_n864), .A3(new_n861), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g445(.A(G290), .B1(new_n567), .B2(new_n572), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n519), .A2(new_n565), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(KEYINPUT72), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n519), .A2(new_n564), .A3(new_n565), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI22_X1  g450(.A1(new_n513), .A2(G87), .B1(G651), .B2(new_n568), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n814), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n871), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(KEYINPUT94), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n582), .A2(G303), .A3(new_n584), .ZN(new_n880));
  AOI21_X1  g455(.A(G303), .B1(new_n582), .B2(new_n584), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT94), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n871), .A2(new_n877), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n879), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n871), .A2(new_n877), .A3(new_n883), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n886), .B1(new_n881), .B2(new_n880), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(KEYINPUT95), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT42), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n613), .A2(G559), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n839), .B(new_n892), .Z(new_n893));
  NAND2_X1  g468(.A1(new_n604), .A2(new_n608), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n613), .A2(G299), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n839), .B(new_n892), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT41), .B1(new_n894), .B2(new_n895), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n894), .A2(KEYINPUT41), .A3(new_n895), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n891), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n897), .A2(new_n891), .A3(new_n901), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n890), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n904), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n906), .A2(new_n889), .A3(new_n902), .ZN(new_n907));
  OAI21_X1  g482(.A(G868), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n837), .A2(G868), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(G295));
  INV_X1    g486(.A(KEYINPUT96), .ZN(new_n912));
  XNOR2_X1  g487(.A(G295), .B(new_n912), .ZN(G331));
  NOR2_X1   g488(.A1(new_n900), .A2(new_n899), .ZN(new_n914));
  OAI21_X1  g489(.A(KEYINPUT97), .B1(G171), .B2(G286), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT97), .ZN(new_n916));
  NAND3_X1  g491(.A1(G168), .A2(new_n916), .A3(G301), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT98), .B1(G168), .B2(G301), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT98), .ZN(new_n920));
  NAND3_X1  g495(.A1(G171), .A2(new_n920), .A3(G286), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT99), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n836), .A2(new_n924), .A3(new_n838), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n924), .B1(new_n836), .B2(new_n838), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n839), .A2(KEYINPUT99), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n915), .A2(new_n917), .B1(new_n919), .B2(new_n921), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n836), .A2(new_n924), .A3(new_n838), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n914), .A2(new_n927), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n896), .B1(new_n927), .B2(new_n931), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n888), .ZN(new_n935));
  AOI21_X1  g510(.A(G37), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT102), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n888), .A2(KEYINPUT101), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT101), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n885), .A2(new_n887), .A3(new_n939), .ZN(new_n940));
  AOI22_X1  g515(.A1(new_n932), .A2(new_n937), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n927), .A2(new_n931), .ZN(new_n942));
  INV_X1    g517(.A(new_n896), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n914), .A2(new_n927), .A3(new_n931), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(KEYINPUT102), .A3(new_n945), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n941), .A2(KEYINPUT103), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT103), .B1(new_n941), .B2(new_n946), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n936), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT100), .B1(new_n932), .B2(new_n933), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT100), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n944), .A2(new_n953), .A3(new_n945), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n938), .A2(new_n940), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n952), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n934), .A2(new_n935), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n867), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT44), .B1(new_n951), .B2(new_n960), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n950), .B(new_n936), .C1(new_n947), .C2(new_n948), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT43), .B1(new_n956), .B2(new_n958), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n961), .A2(new_n966), .ZN(G397));
  XNOR2_X1  g542(.A(new_n764), .B(new_n769), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G1996), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n969), .B1(new_n970), .B2(new_n698), .ZN(new_n971));
  XNOR2_X1  g546(.A(KEYINPUT104), .B(G1384), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT45), .B1(new_n496), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G40), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n467), .A2(new_n974), .A3(new_n472), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n977), .A2(G1996), .A3(new_n697), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT106), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n978), .A2(new_n979), .ZN(new_n981));
  OAI22_X1  g556(.A1(new_n971), .A2(new_n976), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT107), .ZN(new_n983));
  INV_X1    g558(.A(new_n810), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n805), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n805), .A2(new_n984), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n977), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n983), .A2(new_n987), .ZN(new_n988));
  OR3_X1    g563(.A1(new_n976), .A2(G1986), .A3(G290), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n977), .A2(G1986), .A3(G290), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT105), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1384), .ZN(new_n994));
  AND2_X1   g569(.A1(G126), .A2(G2105), .ZN(new_n995));
  INV_X1    g570(.A(G138), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n996), .A2(G2105), .ZN(new_n997));
  INV_X1    g572(.A(new_n485), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n995), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n495), .B1(new_n999), .B2(new_n474), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n998), .B1(new_n461), .B2(G138), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n994), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n489), .A2(new_n490), .B1(new_n492), .B2(new_n494), .ZN(new_n1006));
  AOI21_X1  g581(.A(G1384), .B1(new_n1006), .B2(new_n486), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT109), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1004), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n472), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1010), .A2(G40), .A3(new_n466), .A4(new_n462), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1011), .B1(KEYINPUT50), .B2(new_n1002), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT120), .B1(new_n1013), .B2(new_n710), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n972), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n975), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n732), .A2(KEYINPUT53), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n1017), .A2(new_n1018), .A3(new_n973), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n975), .A2(new_n1016), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT108), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(new_n1007), .B2(KEYINPUT45), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n1007), .A2(new_n1021), .A3(KEYINPUT45), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1020), .B(new_n732), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1019), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1013), .A2(KEYINPUT120), .A3(new_n710), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1015), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT123), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT120), .ZN(new_n1031));
  AOI211_X1 g606(.A(new_n1031), .B(G1961), .C1(new_n1009), .C2(new_n1012), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1014), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT123), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(new_n1034), .A3(new_n1027), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1030), .A2(G171), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT124), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1030), .A2(new_n1035), .A3(KEYINPUT124), .A4(G171), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1013), .A2(new_n710), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT112), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT45), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1042), .B1(new_n1043), .B2(new_n1011), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT45), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1002), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  AOI211_X1 g622(.A(new_n1003), .B(G1384), .C1(new_n1006), .C2(new_n486), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT109), .B1(new_n496), .B2(new_n994), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1045), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1050), .A2(KEYINPUT112), .A3(new_n975), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1044), .A2(new_n1047), .A3(new_n1051), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1040), .B(new_n1041), .C1(new_n1052), .C2(new_n1018), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(G171), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1038), .A2(new_n1039), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT125), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1038), .A2(KEYINPUT125), .A3(new_n1039), .A4(new_n1056), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1004), .A2(new_n1008), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1011), .B1(new_n1062), .B2(new_n1045), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1046), .B1(new_n1063), .B2(KEYINPUT112), .ZN(new_n1064));
  AOI21_X1  g639(.A(G1966), .B1(new_n1064), .B2(new_n1044), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1013), .A2(G2084), .ZN(new_n1066));
  OAI211_X1 g641(.A(G8), .B(G286), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT118), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G8), .ZN(new_n1070));
  INV_X1    g645(.A(G1966), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1051), .A2(new_n1047), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT112), .B1(new_n1050), .B2(new_n975), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1071), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1066), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1070), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1076), .A2(KEYINPUT118), .A3(G286), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1069), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT51), .B1(new_n1076), .B2(KEYINPUT119), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1066), .B1(new_n1052), .B2(new_n1071), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1070), .B1(new_n1080), .B2(G168), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(new_n1080), .B2(new_n1070), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1065), .A2(G286), .A3(new_n1066), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1084), .B(KEYINPUT51), .C1(new_n1085), .C2(new_n1070), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1078), .A2(new_n1082), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT114), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1011), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1089), .B1(new_n1090), .B2(new_n1005), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1002), .A2(KEYINPUT108), .A3(new_n1045), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1017), .B1(new_n1022), .B2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT56), .B(G2072), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1091), .A2(new_n744), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n553), .A2(new_n1096), .A3(new_n557), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1096), .B1(new_n553), .B2(new_n557), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1088), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1020), .B(new_n1094), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n975), .B1(new_n1002), .B2(KEYINPUT50), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1102), .B1(new_n1062), .B2(KEYINPUT50), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1101), .B1(new_n1103), .B2(G1956), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1099), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1104), .A2(KEYINPUT114), .A3(new_n1105), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1099), .B(new_n1101), .C1(new_n1103), .C2(G1956), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1100), .A2(KEYINPUT61), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT61), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT116), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1104), .A2(new_n1110), .A3(new_n1105), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1107), .A2(KEYINPUT116), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1091), .A2(new_n744), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1099), .B1(new_n1113), .B2(new_n1101), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1109), .B(new_n1111), .C1(new_n1112), .C2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1093), .A2(new_n970), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1004), .A2(new_n975), .A3(new_n1008), .ZN(new_n1117));
  XOR2_X1   g692(.A(KEYINPUT58), .B(G1341), .Z(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT59), .B1(new_n1120), .B2(new_n544), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n1122));
  AOI211_X1 g697(.A(new_n1122), .B(new_n543), .C1(new_n1116), .C2(new_n1119), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1108), .A2(new_n1115), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1013), .A2(new_n773), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT113), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n1117), .B2(G2067), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1090), .A2(KEYINPUT113), .A3(new_n769), .A4(new_n975), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1126), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT60), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT117), .B1(new_n1132), .B2(new_n613), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n613), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT117), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1133), .A2(new_n1134), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1134), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1140));
  AOI211_X1 g715(.A(KEYINPUT117), .B(new_n613), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1125), .B1(new_n1138), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1130), .A2(new_n604), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1100), .A2(new_n1144), .A3(new_n1106), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n1107), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT115), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT115), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1145), .A2(new_n1148), .A3(new_n1107), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1087), .B1(new_n1143), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(KEYINPUT121), .B1(new_n1029), .B2(G171), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1053), .A2(G171), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT121), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1033), .A2(new_n1154), .A3(G301), .A4(new_n1027), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1152), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n1055), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1156), .A2(KEYINPUT122), .A3(new_n1055), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n573), .A2(KEYINPUT110), .A3(G1976), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n875), .A2(G1976), .A3(new_n876), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT110), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1070), .B1(new_n1090), .B2(new_n975), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1161), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n573), .A2(G1976), .ZN(new_n1167));
  OR3_X1    g742(.A1(new_n1166), .A2(KEYINPUT52), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1166), .A2(KEYINPUT52), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(G303), .A2(G8), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT55), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1093), .A2(G1971), .ZN(new_n1173));
  INV_X1    g748(.A(G2090), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1173), .B1(new_n1174), .B2(new_n1103), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1172), .B1(new_n1175), .B2(new_n1070), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1013), .A2(G2090), .ZN(new_n1177));
  OAI21_X1  g752(.A(G8), .B1(new_n1177), .B2(new_n1173), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1178), .A2(new_n1172), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT49), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n581), .B(G1981), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(new_n1181), .ZN(new_n1183));
  AND2_X1   g758(.A1(new_n1183), .A2(KEYINPUT111), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1183), .A2(KEYINPUT111), .ZN(new_n1185));
  OAI221_X1 g760(.A(new_n1165), .B1(new_n1181), .B2(new_n1182), .C1(new_n1184), .C2(new_n1185), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1170), .A2(new_n1176), .A3(new_n1180), .A4(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1159), .A2(new_n1160), .A3(new_n1188), .ZN(new_n1189));
  NOR3_X1   g764(.A1(new_n1061), .A2(new_n1151), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1087), .A2(KEYINPUT62), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT62), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1078), .A2(new_n1082), .A3(new_n1086), .A4(new_n1192), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1187), .A2(new_n1153), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1191), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n581), .A2(G1981), .ZN(new_n1196));
  NOR2_X1   g771(.A1(G288), .A2(G1976), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1196), .B1(new_n1186), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1165), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1186), .A2(new_n1169), .A3(new_n1168), .ZN(new_n1200));
  OAI22_X1  g775(.A1(new_n1198), .A2(new_n1199), .B1(new_n1200), .B2(new_n1180), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1200), .A2(new_n1179), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT63), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1203), .B1(new_n1178), .B2(new_n1172), .ZN(new_n1204));
  NAND4_X1  g779(.A1(new_n1202), .A2(G168), .A3(new_n1076), .A4(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1076), .A2(G168), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1203), .B1(new_n1187), .B2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1201), .B1(new_n1205), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1195), .A2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n993), .B1(new_n1190), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT46), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n698), .B1(new_n1211), .B2(G1996), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n977), .B1(new_n969), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n977), .A2(new_n970), .ZN(new_n1214));
  AND3_X1   g789(.A1(new_n1214), .A2(KEYINPUT126), .A3(new_n1211), .ZN(new_n1215));
  AOI21_X1  g790(.A(KEYINPUT126), .B1(new_n1214), .B2(new_n1211), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1213), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  XOR2_X1   g792(.A(new_n1217), .B(KEYINPUT47), .Z(new_n1218));
  NAND2_X1  g793(.A1(new_n983), .A2(new_n986), .ZN(new_n1219));
  OR2_X1    g794(.A1(new_n764), .A2(G2067), .ZN(new_n1220));
  AOI21_X1  g795(.A(new_n976), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g796(.A(new_n989), .B(KEYINPUT48), .ZN(new_n1222));
  AOI211_X1 g797(.A(new_n1218), .B(new_n1221), .C1(new_n988), .C2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1210), .A2(new_n1223), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g799(.A(KEYINPUT127), .ZN(new_n1226));
  INV_X1    g800(.A(G319), .ZN(new_n1227));
  NOR3_X1   g801(.A1(G401), .A2(new_n1227), .A3(G227), .ZN(new_n1228));
  NAND3_X1  g802(.A1(new_n869), .A2(new_n1228), .A3(new_n691), .ZN(new_n1229));
  INV_X1    g803(.A(new_n1229), .ZN(new_n1230));
  AOI21_X1  g804(.A(new_n1226), .B1(new_n964), .B2(new_n1230), .ZN(new_n1231));
  AOI211_X1 g805(.A(KEYINPUT127), .B(new_n1229), .C1(new_n962), .C2(new_n963), .ZN(new_n1232));
  NOR2_X1   g806(.A1(new_n1231), .A2(new_n1232), .ZN(G308));
  NAND2_X1  g807(.A1(new_n964), .A2(new_n1230), .ZN(G225));
endmodule


