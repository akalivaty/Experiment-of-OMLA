//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n188), .A2(G143), .ZN(new_n194));
  AOI22_X1  g008(.A1(new_n192), .A2(new_n193), .B1(KEYINPUT1), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n189), .A2(new_n191), .A3(new_n196), .A4(G128), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(G125), .ZN(new_n199));
  XNOR2_X1  g013(.A(G143), .B(G146), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT0), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(new_n193), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT0), .A2(G128), .ZN(new_n203));
  XNOR2_X1  g017(.A(new_n202), .B(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n199), .B1(new_n204), .B2(G125), .ZN(new_n205));
  INV_X1    g019(.A(G953), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G224), .ZN(new_n207));
  XNOR2_X1  g021(.A(new_n205), .B(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT67), .ZN(new_n209));
  XNOR2_X1  g023(.A(G116), .B(G119), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT2), .B(G113), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n209), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n212), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(KEYINPUT67), .A3(new_n210), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G104), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT3), .B1(new_n217), .B2(G107), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n219));
  INV_X1    g033(.A(G107), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(G104), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n217), .A2(G107), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n218), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  XOR2_X1   g037(.A(KEYINPUT81), .B(G101), .Z(new_n224));
  NAND2_X1  g038(.A1(new_n220), .A2(G104), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n222), .ZN(new_n226));
  AOI22_X1  g040(.A1(new_n223), .A2(new_n224), .B1(G101), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT5), .ZN(new_n228));
  INV_X1    g042(.A(G119), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n229), .A3(G116), .ZN(new_n230));
  OAI211_X1 g044(.A(G113), .B(new_n230), .C1(new_n211), .C2(new_n228), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n216), .A2(new_n227), .A3(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n218), .A2(new_n221), .A3(new_n222), .ZN(new_n233));
  AOI21_X1  g047(.A(KEYINPUT4), .B1(new_n233), .B2(G101), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n224), .A2(new_n218), .A3(new_n221), .A4(new_n222), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(G101), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n234), .B1(new_n237), .B2(KEYINPUT4), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT66), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n210), .B1(new_n214), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n212), .A2(KEYINPUT66), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n213), .A2(new_n215), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n232), .B1(new_n238), .B2(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(G110), .B(G122), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n232), .B(new_n244), .C1(new_n238), .C2(new_n242), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(KEYINPUT6), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT6), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n243), .A2(new_n249), .A3(new_n245), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n208), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT85), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT85), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n208), .A2(new_n248), .A3(new_n253), .A4(new_n250), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n207), .B1(KEYINPUT86), .B2(KEYINPUT7), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n256), .B1(KEYINPUT86), .B2(KEYINPUT7), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n205), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n206), .A2(KEYINPUT87), .A3(G224), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT7), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT87), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n260), .B1(new_n261), .B2(new_n207), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n258), .B1(new_n205), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n216), .A2(new_n231), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n226), .A2(G101), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n235), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n232), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n244), .B(KEYINPUT8), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n263), .A2(new_n247), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G902), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(G210), .B1(G237), .B2(G902), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n255), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n274), .B1(new_n255), .B2(new_n273), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n187), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT84), .B(G469), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT82), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n197), .A2(new_n279), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n200), .A2(KEYINPUT82), .A3(new_n196), .A4(G128), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n195), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n227), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT83), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT83), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n282), .A2(new_n227), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n198), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n284), .A2(new_n286), .B1(new_n266), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G131), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT11), .ZN(new_n290));
  INV_X1    g104(.A(G137), .ZN(new_n291));
  AND2_X1   g105(.A1(KEYINPUT64), .A2(G134), .ZN(new_n292));
  NOR2_X1   g106(.A1(KEYINPUT64), .A2(G134), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n290), .B(new_n291), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n290), .B1(G134), .B2(new_n291), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n292), .A2(new_n293), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G137), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n289), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT65), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT64), .ZN(new_n302));
  INV_X1    g116(.A(G134), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(KEYINPUT64), .A2(G134), .ZN(new_n305));
  AOI21_X1  g119(.A(G137), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n295), .B1(new_n306), .B2(new_n290), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n304), .A2(new_n305), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n289), .B1(new_n308), .B2(new_n291), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n301), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(G131), .B1(new_n298), .B2(G137), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n297), .A2(new_n311), .A3(KEYINPUT65), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n300), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT12), .B1(new_n288), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n198), .A2(KEYINPUT10), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n315), .A2(new_n266), .ZN(new_n316));
  INV_X1    g130(.A(new_n238), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n202), .A2(new_n203), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n202), .A2(new_n203), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n316), .B1(new_n317), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT10), .ZN(new_n322));
  INV_X1    g136(.A(new_n286), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n285), .B1(new_n282), .B2(new_n227), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n321), .A2(new_n325), .A3(new_n313), .ZN(new_n326));
  OAI22_X1  g140(.A1(new_n323), .A2(new_n324), .B1(new_n227), .B2(new_n198), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT12), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n297), .A2(new_n299), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G131), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n297), .A2(new_n311), .A3(KEYINPUT65), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT65), .B1(new_n297), .B2(new_n311), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n327), .A2(new_n328), .A3(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(G110), .B(G140), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n206), .A2(G227), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n335), .B(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n314), .A2(new_n326), .A3(new_n334), .A4(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT10), .B1(new_n284), .B2(new_n286), .ZN(new_n341));
  OAI22_X1  g155(.A1(new_n238), .A2(new_n204), .B1(new_n266), .B2(new_n315), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n333), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n338), .B1(new_n343), .B2(new_n326), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n272), .B(new_n278), .C1(new_n340), .C2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n314), .A2(new_n326), .A3(new_n334), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n337), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n343), .A2(new_n326), .A3(new_n338), .ZN(new_n348));
  AOI21_X1  g162(.A(G902), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G469), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n345), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G221), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT9), .B(G234), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n352), .B1(new_n354), .B2(new_n272), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n277), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G237), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n359), .A2(new_n206), .A3(G214), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n360), .B(new_n190), .ZN(new_n361));
  NAND2_X1  g175(.A1(KEYINPUT18), .A2(G131), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n361), .B(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G140), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G125), .ZN(new_n365));
  INV_X1    g179(.A(G125), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G140), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT78), .ZN(new_n369));
  XNOR2_X1  g183(.A(G125), .B(G140), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT78), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n369), .A2(new_n372), .A3(new_n188), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT77), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n366), .A2(KEYINPUT77), .A3(G140), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(G146), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT88), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n373), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n378), .B1(new_n373), .B2(new_n377), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n363), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n375), .A2(KEYINPUT16), .A3(new_n376), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT16), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n365), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G146), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n361), .A2(G131), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT17), .ZN(new_n389));
  OR2_X1    g203(.A1(new_n360), .A2(new_n190), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n360), .A2(new_n190), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n289), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n388), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n383), .A2(new_n188), .A3(new_n385), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n361), .A2(KEYINPUT17), .A3(G131), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n387), .A2(new_n393), .A3(new_n394), .A4(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(G113), .B(G122), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(new_n217), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n382), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n398), .B1(new_n382), .B2(new_n396), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n272), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G475), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT20), .ZN(new_n403));
  NOR2_X1   g217(.A1(G475), .A2(G902), .ZN(new_n404));
  AOI22_X1  g218(.A1(new_n386), .A2(G146), .B1(new_n388), .B2(new_n392), .ZN(new_n405));
  XNOR2_X1  g219(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n369), .A2(new_n372), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT90), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n375), .A2(KEYINPUT19), .A3(new_n376), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT90), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n369), .A2(new_n372), .A3(new_n410), .A4(new_n406), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n408), .A2(new_n188), .A3(new_n409), .A4(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n405), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n398), .B1(new_n413), .B2(new_n382), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n403), .B(new_n404), .C1(new_n399), .C2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n382), .A2(new_n396), .A3(new_n398), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n373), .A2(new_n377), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT88), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n379), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n420), .A2(new_n363), .B1(new_n405), .B2(new_n412), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n417), .B1(new_n421), .B2(new_n398), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n403), .B1(new_n422), .B2(new_n404), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n402), .B1(new_n416), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT91), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g240(.A(KEYINPUT91), .B(new_n402), .C1(new_n416), .C2(new_n423), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(KEYINPUT93), .A2(G952), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(KEYINPUT93), .A2(G952), .ZN(new_n431));
  AOI21_X1  g245(.A(G953), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G234), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n432), .B1(new_n433), .B2(new_n359), .ZN(new_n434));
  XOR2_X1   g248(.A(KEYINPUT21), .B(G898), .Z(new_n435));
  AOI211_X1 g249(.A(new_n272), .B(new_n206), .C1(G234), .C2(G237), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n434), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G116), .B(G122), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(new_n220), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n190), .A2(G128), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT13), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n193), .A2(G143), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n441), .A2(new_n442), .ZN(new_n446));
  OAI21_X1  g260(.A(G134), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n298), .A2(new_n441), .A3(new_n444), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n440), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n441), .A2(new_n444), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n308), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G116), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(KEYINPUT14), .A3(G122), .ZN(new_n454));
  INV_X1    g268(.A(new_n439), .ZN(new_n455));
  OAI211_X1 g269(.A(G107), .B(new_n454), .C1(new_n455), .C2(KEYINPUT14), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n452), .B(new_n456), .C1(G107), .C2(new_n455), .ZN(new_n457));
  INV_X1    g271(.A(G217), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n353), .A2(new_n458), .A3(G953), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n449), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n459), .B1(new_n457), .B2(new_n449), .ZN(new_n461));
  OR2_X1    g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT92), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(new_n463), .A3(new_n272), .ZN(new_n464));
  INV_X1    g278(.A(G478), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(KEYINPUT15), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n464), .B(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n428), .A2(new_n438), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n358), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(G119), .B(G128), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(KEYINPUT74), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT24), .B(G110), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n193), .A2(KEYINPUT23), .A3(G119), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n229), .A2(G128), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n229), .A2(G128), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n475), .B(new_n476), .C1(new_n477), .C2(KEYINPUT23), .ZN(new_n478));
  OAI22_X1  g292(.A1(new_n472), .A2(new_n474), .B1(G110), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n387), .A2(new_n479), .A3(new_n373), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n387), .A2(new_n394), .ZN(new_n481));
  INV_X1    g295(.A(new_n472), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n481), .B1(new_n482), .B2(new_n473), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT75), .ZN(new_n484));
  OR2_X1    g298(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n478), .A2(new_n484), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(G110), .A3(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(KEYINPUT76), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n480), .B1(new_n483), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT22), .B(G137), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n352), .A2(new_n433), .A3(G953), .ZN(new_n491));
  XOR2_X1   g305(.A(new_n490), .B(new_n491), .Z(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n480), .B(new_n492), .C1(new_n483), .C2(new_n488), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n494), .A2(new_n272), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT25), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n494), .A2(KEYINPUT25), .A3(new_n272), .A4(new_n495), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n458), .B1(G234), .B2(new_n272), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n494), .A2(new_n495), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n501), .A2(G902), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(KEYINPUT79), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT28), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n303), .A2(G137), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n298), .B2(G137), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n197), .A2(new_n195), .B1(new_n512), .B2(G131), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n513), .B1(new_n331), .B2(new_n332), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n514), .B1(new_n313), .B2(new_n204), .ZN(new_n515));
  INV_X1    g329(.A(new_n242), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n242), .B(new_n514), .C1(new_n313), .C2(new_n204), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n510), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n510), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n359), .A2(new_n206), .A3(G210), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n523), .B(KEYINPUT27), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT26), .B(G101), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n524), .B(new_n525), .ZN(new_n526));
  OAI211_X1 g340(.A(KEYINPUT30), .B(new_n514), .C1(new_n313), .C2(new_n204), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n310), .A2(new_n312), .ZN(new_n528));
  AOI22_X1  g342(.A1(new_n333), .A2(new_n320), .B1(new_n528), .B2(new_n513), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n527), .B(new_n516), .C1(new_n529), .C2(KEYINPUT30), .ZN(new_n530));
  INV_X1    g344(.A(new_n526), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n531), .B1(new_n529), .B2(new_n242), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  OAI22_X1  g347(.A1(new_n522), .A2(new_n526), .B1(KEYINPUT31), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT68), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n530), .A2(new_n536), .A3(new_n532), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n536), .B1(new_n530), .B2(new_n532), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT69), .B1(new_n539), .B2(KEYINPUT31), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n533), .A2(KEYINPUT68), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n530), .A2(new_n536), .A3(new_n532), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n541), .A2(KEYINPUT69), .A3(KEYINPUT31), .A4(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n535), .B1(new_n540), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT70), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n541), .A2(KEYINPUT31), .A3(new_n542), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT69), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n543), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT70), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(new_n551), .A3(new_n535), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n546), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(G472), .A2(G902), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT32), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n554), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT32), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n551), .B1(new_n550), .B2(new_n535), .ZN(new_n559));
  AOI211_X1 g373(.A(KEYINPUT70), .B(new_n534), .C1(new_n549), .C2(new_n543), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT71), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT29), .ZN(new_n563));
  INV_X1    g377(.A(new_n518), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT30), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n515), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n565), .B1(new_n528), .B2(new_n513), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n333), .A2(new_n320), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n242), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n564), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n563), .B1(new_n570), .B2(new_n526), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n519), .A2(new_n521), .A3(new_n531), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n562), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n242), .B1(new_n568), .B2(new_n514), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT28), .B1(new_n564), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(new_n520), .A3(new_n526), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n530), .A2(new_n518), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n531), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n576), .A2(new_n578), .A3(KEYINPUT71), .A4(new_n563), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n531), .A2(new_n563), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n520), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT72), .B1(new_n519), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n580), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n518), .B2(new_n510), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT72), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n575), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(G902), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n573), .A2(new_n579), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(G472), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT73), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n588), .A2(KEYINPUT73), .A3(G472), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n561), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n509), .B1(new_n555), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT80), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n556), .B1(new_n546), .B2(new_n552), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n561), .B(new_n593), .C1(new_n598), .C2(KEYINPUT32), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n599), .A2(KEYINPUT80), .A3(new_n509), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n470), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(new_n224), .ZN(G3));
  OAI21_X1  g416(.A(new_n272), .B1(new_n559), .B2(new_n560), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n598), .B1(G472), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n357), .A2(new_n508), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n428), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT94), .ZN(new_n608));
  AOI21_X1  g422(.A(KEYINPUT33), .B1(new_n462), .B2(new_n608), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n608), .B(KEYINPUT33), .C1(new_n460), .C2(new_n461), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  OAI211_X1 g425(.A(G478), .B(new_n272), .C1(new_n609), .C2(new_n611), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n462), .A2(new_n272), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n612), .B1(G478), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n607), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n277), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n438), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n606), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT34), .B(G104), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G6));
  INV_X1    g434(.A(new_n606), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n617), .A2(new_n424), .A3(new_n468), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT35), .B(G107), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G9));
  INV_X1    g439(.A(new_n470), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n489), .A2(KEYINPUT95), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT95), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n628), .B(new_n480), .C1(new_n483), .C2(new_n488), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n493), .A2(KEYINPUT36), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n627), .A2(new_n631), .A3(new_n629), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n500), .A2(new_n501), .B1(new_n635), .B2(new_n506), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n604), .A2(new_n626), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT37), .B(G110), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G12));
  INV_X1    g454(.A(new_n424), .ZN(new_n641));
  INV_X1    g455(.A(new_n434), .ZN(new_n642));
  INV_X1    g456(.A(G900), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n642), .B1(new_n643), .B2(new_n436), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n641), .A2(new_n467), .A3(new_n645), .ZN(new_n646));
  NOR4_X1   g460(.A1(new_n277), .A2(new_n357), .A3(new_n636), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n599), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G128), .ZN(G30));
  NAND2_X1  g463(.A1(new_n255), .A2(new_n273), .ZN(new_n650));
  INV_X1    g464(.A(new_n274), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n255), .A2(new_n273), .A3(new_n274), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT38), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n652), .A2(KEYINPUT38), .A3(new_n653), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n607), .A2(new_n467), .ZN(new_n660));
  INV_X1    g474(.A(new_n187), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n660), .A2(new_n661), .A3(new_n637), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(new_n644), .B(KEYINPUT39), .Z(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n357), .A2(new_n665), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n666), .A2(KEYINPUT40), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(KEYINPUT40), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n663), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n554), .B1(new_n559), .B2(new_n560), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n557), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n526), .B1(new_n517), .B2(new_n518), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n537), .A2(new_n538), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g487(.A(G472), .B1(new_n673), .B2(G902), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n671), .A2(new_n561), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n669), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(KEYINPUT96), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT96), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n669), .A2(new_n678), .A3(new_n675), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(new_n190), .ZN(G45));
  NAND4_X1  g495(.A1(new_n426), .A2(new_n614), .A3(new_n427), .A4(new_n645), .ZN(new_n682));
  NOR4_X1   g496(.A1(new_n277), .A2(new_n357), .A3(new_n682), .A4(new_n636), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n599), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G146), .ZN(G48));
  AND2_X1   g499(.A1(new_n561), .A2(new_n593), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n508), .B1(new_n686), .B2(new_n671), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n617), .A2(new_n615), .ZN(new_n688));
  INV_X1    g502(.A(new_n345), .ZN(new_n689));
  INV_X1    g503(.A(new_n344), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n339), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n350), .B1(new_n691), .B2(new_n272), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n356), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n687), .A2(new_n688), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT41), .B(G113), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G15));
  NAND3_X1  g512(.A1(new_n687), .A2(new_n622), .A3(new_n695), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G116), .ZN(G18));
  NOR2_X1   g514(.A1(new_n694), .A2(new_n277), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n701), .A2(new_n469), .A3(new_n637), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n599), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT97), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT97), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n599), .A2(new_n705), .A3(new_n702), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT98), .B(G119), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G21));
  INV_X1    g523(.A(new_n660), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n701), .A2(new_n438), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n603), .A2(G472), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n556), .B1(new_n535), .B2(new_n547), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n508), .B(KEYINPUT99), .ZN(new_n715));
  AND4_X1   g529(.A1(KEYINPUT100), .A2(new_n712), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n713), .B1(new_n603), .B2(G472), .ZN(new_n717));
  AOI21_X1  g531(.A(KEYINPUT100), .B1(new_n717), .B2(new_n715), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n711), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G122), .ZN(G24));
  NOR3_X1   g534(.A1(new_n694), .A2(new_n277), .A3(new_n682), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n712), .A2(new_n637), .A3(new_n714), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G125), .ZN(G27));
  INV_X1    g537(.A(new_n682), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n652), .A2(new_n187), .A3(new_n653), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n348), .A2(KEYINPUT101), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT101), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n343), .A2(new_n326), .A3(new_n728), .A4(new_n338), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n347), .A2(new_n727), .A3(G469), .A4(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(G469), .A2(G902), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n345), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n356), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT102), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n732), .A2(KEYINPUT102), .A3(new_n356), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n726), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n599), .A2(new_n509), .A3(new_n724), .A4(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT42), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n737), .A2(new_n740), .A3(new_n682), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n561), .A2(KEYINPUT103), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT103), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n553), .A2(new_n744), .A3(new_n558), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n671), .A2(new_n593), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n715), .B(new_n742), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n741), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G131), .ZN(G33));
  INV_X1    g564(.A(new_n646), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n599), .A2(new_n509), .A3(new_n751), .A4(new_n738), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G134), .ZN(G36));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n428), .A2(new_n614), .ZN(new_n755));
  OR2_X1    g569(.A1(new_n755), .A2(KEYINPUT43), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(KEYINPUT43), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n637), .A3(new_n757), .ZN(new_n758));
  OR3_X1    g572(.A1(new_n604), .A2(new_n754), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n726), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT105), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n754), .B1(new_n604), .B2(new_n758), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n759), .A2(KEYINPUT105), .A3(new_n726), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT106), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n347), .A2(new_n727), .A3(KEYINPUT45), .A4(new_n729), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n347), .A2(new_n348), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n768), .B(G469), .C1(new_n769), .C2(KEYINPUT45), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n770), .A2(new_n731), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n771), .A2(KEYINPUT46), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n345), .B1(new_n771), .B2(KEYINPUT46), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n356), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n774), .A2(new_n665), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT104), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n762), .A2(KEYINPUT106), .A3(new_n763), .A4(new_n764), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n767), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G137), .ZN(G39));
  OR4_X1    g593(.A1(new_n599), .A2(new_n509), .A3(new_n682), .A4(new_n725), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n774), .B(KEYINPUT47), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(new_n364), .ZN(G42));
  NAND3_X1  g597(.A1(new_n715), .A2(new_n356), .A3(new_n187), .ZN(new_n784));
  INV_X1    g598(.A(new_n693), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n755), .B1(new_n785), .B2(KEYINPUT49), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n786), .B1(KEYINPUT49), .B2(new_n785), .ZN(new_n787));
  OR4_X1    g601(.A1(new_n675), .A2(new_n784), .A3(new_n659), .A4(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT51), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n756), .A2(new_n757), .ZN(new_n790));
  INV_X1    g604(.A(new_n718), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n717), .A2(KEYINPUT100), .A3(new_n715), .ZN(new_n792));
  AOI211_X1 g606(.A(new_n434), .B(new_n790), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n793), .A2(new_n726), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n693), .A2(new_n355), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT111), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n781), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n694), .A2(new_n725), .A3(new_n434), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n757), .A3(new_n756), .ZN(new_n800));
  XOR2_X1   g614(.A(new_n800), .B(KEYINPUT114), .Z(new_n801));
  NAND3_X1  g615(.A1(new_n801), .A2(new_n637), .A3(new_n717), .ZN(new_n802));
  XOR2_X1   g616(.A(new_n802), .B(KEYINPUT115), .Z(new_n803));
  NAND2_X1  g617(.A1(new_n799), .A2(new_n509), .ZN(new_n804));
  NOR4_X1   g618(.A1(new_n675), .A2(new_n607), .A3(new_n614), .A4(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT116), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n694), .A2(new_n187), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n658), .B1(new_n808), .B2(KEYINPUT112), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(KEYINPUT112), .B2(new_n808), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n793), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT50), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n793), .A2(KEYINPUT50), .A3(new_n810), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n813), .A2(KEYINPUT113), .A3(new_n814), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n807), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n798), .B1(new_n819), .B2(KEYINPUT117), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n821));
  AOI211_X1 g635(.A(new_n821), .B(new_n807), .C1(new_n817), .C2(new_n818), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n789), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(KEYINPUT107), .B1(new_n601), .B2(new_n618), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n599), .A2(KEYINPUT80), .A3(new_n509), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT80), .B1(new_n599), .B2(new_n509), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n626), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT107), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n621), .A2(new_n688), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n467), .B(KEYINPUT108), .Z(new_n831));
  OR2_X1    g645(.A1(new_n831), .A2(new_n607), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n617), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n638), .B1(new_n606), .B2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n824), .A2(new_n830), .A3(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n637), .A2(new_n831), .A3(new_n641), .A4(new_n645), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n838), .A2(new_n357), .A3(new_n725), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n599), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n717), .A2(new_n637), .A3(new_n724), .A4(new_n738), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n752), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n749), .A2(new_n842), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n687), .B(new_n695), .C1(new_n688), .C2(new_n622), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n707), .A2(new_n844), .A3(new_n719), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  OAI22_X1  g660(.A1(new_n555), .A2(new_n594), .B1(new_n647), .B2(new_n683), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n636), .A2(new_n645), .ZN(new_n848));
  NOR4_X1   g662(.A1(new_n660), .A2(new_n848), .A3(new_n277), .A4(new_n733), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n561), .A2(new_n674), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n849), .B1(new_n555), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n847), .A2(new_n851), .A3(new_n722), .ZN(new_n852));
  XOR2_X1   g666(.A(KEYINPUT109), .B(KEYINPUT52), .Z(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT52), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n847), .A2(new_n851), .A3(new_n856), .A4(new_n722), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n854), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n837), .A2(new_n846), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n827), .A2(new_n829), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n835), .B1(new_n860), .B2(KEYINPUT107), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n852), .B(new_n856), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n861), .A2(new_n846), .A3(new_n830), .A4(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  OAI211_X1 g678(.A(KEYINPUT54), .B(new_n859), .C1(new_n864), .C2(new_n855), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n854), .A2(KEYINPUT53), .A3(new_n857), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n843), .A2(new_n866), .A3(new_n845), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n837), .A2(new_n867), .A3(KEYINPUT110), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT110), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n854), .A2(KEYINPUT53), .A3(new_n857), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n707), .A2(new_n719), .A3(new_n844), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n752), .A2(new_n840), .A3(new_n841), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n748), .B2(new_n741), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n870), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n824), .A2(new_n830), .A3(new_n836), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n869), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n868), .A2(new_n876), .B1(new_n855), .B2(new_n863), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n746), .A2(new_n747), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n880), .A2(new_n715), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n801), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT48), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n793), .A2(new_n701), .ZN(new_n884));
  OR3_X1    g698(.A1(new_n675), .A2(new_n615), .A3(new_n804), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n883), .A2(new_n432), .A3(new_n884), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n781), .A2(new_n795), .ZN(new_n887));
  AOI211_X1 g701(.A(new_n789), .B(new_n807), .C1(new_n794), .C2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n886), .B1(new_n888), .B2(new_n815), .ZN(new_n889));
  AND4_X1   g703(.A1(new_n823), .A2(new_n865), .A3(new_n879), .A4(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(G952), .A2(G953), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n788), .B1(new_n890), .B2(new_n891), .ZN(G75));
  INV_X1    g706(.A(KEYINPUT56), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n868), .A2(new_n876), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n863), .A2(new_n855), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(G902), .ZN(new_n897));
  INV_X1    g711(.A(G210), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n893), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n248), .A2(new_n250), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(new_n208), .ZN(new_n901));
  XNOR2_X1  g715(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n901), .B(new_n902), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n899), .A2(new_n903), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n206), .A2(G952), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(G51));
  NAND2_X1  g721(.A1(new_n896), .A2(KEYINPUT54), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n908), .A2(new_n879), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n731), .B(KEYINPUT57), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n691), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n897), .A2(new_n770), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n906), .B1(new_n911), .B2(new_n912), .ZN(G54));
  NAND4_X1  g727(.A1(new_n896), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n914));
  INV_X1    g728(.A(new_n422), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n916), .A2(new_n917), .A3(new_n906), .ZN(G60));
  NAND2_X1  g732(.A1(G478), .A2(G902), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT59), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n920), .B1(new_n609), .B2(new_n611), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n908), .B2(new_n879), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT119), .B1(new_n922), .B2(new_n906), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n879), .A2(new_n865), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n920), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n609), .A2(new_n611), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n922), .A2(KEYINPUT119), .A3(new_n906), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(G63));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n931));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT121), .ZN(new_n933));
  XOR2_X1   g747(.A(KEYINPUT120), .B(KEYINPUT60), .Z(new_n934));
  XOR2_X1   g748(.A(new_n933), .B(new_n934), .Z(new_n935));
  AOI21_X1  g749(.A(new_n503), .B1(new_n896), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(KEYINPUT124), .B1(new_n936), .B2(new_n906), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT124), .ZN(new_n938));
  INV_X1    g752(.A(new_n906), .ZN(new_n939));
  INV_X1    g753(.A(new_n935), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n894), .B2(new_n895), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n938), .B(new_n939), .C1(new_n941), .C2(new_n503), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n937), .A2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT122), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n941), .B2(new_n635), .ZN(new_n945));
  INV_X1    g759(.A(new_n635), .ZN(new_n946));
  NOR4_X1   g760(.A1(new_n877), .A2(KEYINPUT122), .A3(new_n946), .A4(new_n940), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n945), .A2(new_n947), .A3(KEYINPUT123), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n931), .B1(new_n943), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT61), .B1(new_n936), .B2(new_n906), .ZN(new_n950));
  OAI221_X1 g764(.A(new_n950), .B1(KEYINPUT123), .B2(KEYINPUT61), .C1(new_n947), .C2(new_n945), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n951), .ZN(G66));
  NAND2_X1  g766(.A1(new_n837), .A2(new_n871), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT125), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n954), .A2(G953), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n206), .B1(new_n435), .B2(G224), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(G898), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n900), .B1(new_n958), .B2(G953), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n957), .B(new_n959), .ZN(G69));
  AND2_X1   g774(.A1(new_n847), .A2(new_n722), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n677), .A2(new_n679), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(KEYINPUT62), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n597), .A2(new_n600), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n666), .A2(new_n726), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n965), .B1(new_n615), .B2(new_n832), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n782), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n963), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n962), .A2(KEYINPUT62), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n778), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n970), .A2(KEYINPUT126), .A3(new_n778), .ZN(new_n974));
  AOI21_X1  g788(.A(G953), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n566), .A2(new_n527), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n976), .B(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(KEYINPUT127), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n974), .ZN(new_n980));
  AOI21_X1  g794(.A(KEYINPUT126), .B1(new_n970), .B2(new_n778), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n206), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT127), .ZN(new_n983));
  INV_X1    g797(.A(new_n978), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n776), .A2(new_n616), .A3(new_n710), .A4(new_n881), .ZN(new_n986));
  INV_X1    g800(.A(new_n752), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n782), .A2(new_n987), .ZN(new_n988));
  AND4_X1   g802(.A1(new_n749), .A2(new_n986), .A3(new_n961), .A4(new_n988), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n989), .A2(new_n778), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n206), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n991), .B(new_n978), .C1(new_n643), .C2(new_n206), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n979), .A2(new_n985), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n206), .B1(G227), .B2(G900), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n994), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n979), .A2(new_n985), .A3(new_n996), .A4(new_n992), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n995), .A2(new_n997), .ZN(G72));
  NAND3_X1  g812(.A1(new_n954), .A2(new_n973), .A3(new_n974), .ZN(new_n999));
  NAND2_X1  g813(.A1(G472), .A2(G902), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT63), .Z(new_n1001));
  AOI211_X1 g815(.A(new_n531), .B(new_n570), .C1(new_n999), .C2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1001), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1003), .B1(new_n954), .B2(new_n990), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n1004), .A2(new_n526), .A3(new_n577), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1003), .B1(new_n539), .B2(new_n578), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n859), .B(new_n1006), .C1(new_n864), .C2(new_n855), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(new_n939), .ZN(new_n1008));
  NOR3_X1   g822(.A1(new_n1002), .A2(new_n1005), .A3(new_n1008), .ZN(G57));
endmodule


