//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 1 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1204, new_n1205, new_n1206, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  XOR2_X1   g0008(.A(KEYINPUT67), .B(G244), .Z(new_n209));
  AOI22_X1  g0009(.A1(new_n209), .A2(G77), .B1(G116), .B2(G270), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G107), .A2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n210), .B(new_n211), .C1(new_n201), .C2(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G68), .B2(G238), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G97), .A2(G257), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G87), .A2(G250), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G58), .A2(G232), .ZN(new_n217));
  NAND4_X1  g0017(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G20), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT68), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(G50), .B1(G58), .B2(G68), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT66), .Z(new_n228));
  AOI21_X1  g0028(.A(new_n223), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(new_n219), .ZN(new_n230));
  INV_X1    g0030(.A(G13), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n230), .A2(KEYINPUT64), .A3(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(KEYINPUT64), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n233), .B1(new_n219), .B2(G13), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n235), .B(G250), .C1(G257), .C2(G264), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT65), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT0), .ZN(new_n238));
  NAND3_X1  g0038(.A1(new_n222), .A2(new_n229), .A3(new_n238), .ZN(new_n239));
  INV_X1    g0039(.A(new_n239), .ZN(G361));
  XOR2_X1   g0040(.A(G226), .B(G232), .Z(new_n241));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT70), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G250), .B(G257), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G264), .B(G270), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G358));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n251), .B(new_n252), .Z(new_n253));
  XNOR2_X1  g0053(.A(G68), .B(G77), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G50), .B(G58), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XOR2_X1   g0056(.A(new_n253), .B(new_n256), .Z(G351));
  NAND2_X1  g0057(.A1(new_n204), .A2(G20), .ZN(new_n258));
  INV_X1    g0058(.A(G150), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n225), .A2(G33), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT8), .B(G58), .ZN(new_n263));
  OAI221_X1 g0063(.A(new_n258), .B1(new_n259), .B2(new_n261), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n224), .B1(new_n219), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G13), .A3(G20), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT72), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT72), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n271), .A2(new_n268), .A3(G13), .A4(G20), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n201), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n270), .A2(new_n272), .ZN(new_n275));
  INV_X1    g0075(.A(new_n266), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n275), .B(new_n276), .C1(G1), .C2(new_n225), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n267), .B(new_n274), .C1(new_n201), .C2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n278), .B(KEYINPUT9), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT3), .B(G33), .ZN(new_n280));
  INV_X1    g0080(.A(G223), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  AND2_X1   g0082(.A1(KEYINPUT71), .A2(G1698), .ZN(new_n283));
  NOR2_X1   g0083(.A1(KEYINPUT71), .A2(G1698), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G222), .ZN(new_n286));
  OAI221_X1 g0086(.A(new_n280), .B1(new_n281), .B2(new_n282), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G41), .ZN(new_n288));
  OAI211_X1 g0088(.A(G1), .B(G13), .C1(new_n265), .C2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n287), .B(new_n290), .C1(G77), .C2(new_n280), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n268), .B1(G41), .B2(G45), .ZN(new_n292));
  INV_X1    g0092(.A(G274), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n289), .A2(new_n292), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n291), .B(new_n295), .C1(new_n212), .C2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(G200), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n279), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT73), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n301), .A2(new_n305), .A3(new_n303), .ZN(new_n308));
  INV_X1    g0108(.A(G169), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n297), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n310), .B(new_n278), .C1(G179), .C2(new_n297), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n307), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT81), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G33), .A2(G87), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n212), .A2(new_n282), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT71), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n282), .ZN(new_n317));
  NAND2_X1  g0117(.A1(KEYINPUT71), .A2(G1698), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n315), .B1(new_n319), .B2(G223), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT3), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n321), .A2(KEYINPUT80), .A3(G33), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT80), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n323), .B1(KEYINPUT3), .B2(new_n265), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n322), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n314), .B1(new_n320), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n294), .B1(new_n327), .B2(new_n290), .ZN(new_n328));
  INV_X1    g0128(.A(G232), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n296), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n309), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT80), .B1(new_n321), .B2(G33), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n321), .A2(G33), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n281), .B1(new_n317), .B2(new_n318), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n322), .B(new_n335), .C1(new_n336), .C2(new_n315), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n289), .B1(new_n337), .B2(new_n314), .ZN(new_n338));
  INV_X1    g0138(.A(G179), .ZN(new_n339));
  NOR4_X1   g0139(.A1(new_n338), .A2(new_n339), .A3(new_n294), .A4(new_n330), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n313), .B1(new_n332), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n202), .A2(new_n203), .ZN(new_n342));
  NOR2_X1   g0142(.A1(G58), .A2(G68), .ZN(new_n343));
  OAI21_X1  g0143(.A(G20), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n260), .A2(G159), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(G20), .B1(new_n335), .B2(new_n322), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT7), .ZN(new_n349));
  OAI21_X1  g0149(.A(G68), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AND3_X1   g0150(.A1(new_n321), .A2(KEYINPUT80), .A3(G33), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n351), .B1(new_n334), .B2(new_n333), .ZN(new_n352));
  NOR3_X1   g0152(.A1(new_n352), .A2(KEYINPUT7), .A3(G20), .ZN(new_n353));
  OAI211_X1 g0153(.A(KEYINPUT16), .B(new_n347), .C1(new_n350), .C2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT16), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n349), .B1(new_n280), .B2(G20), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n334), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n203), .B1(new_n356), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n355), .B1(new_n360), .B2(new_n346), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n354), .A2(new_n266), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n263), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n277), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n273), .B2(new_n363), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  OAI22_X1  g0166(.A1(new_n285), .A2(new_n281), .B1(new_n212), .B2(new_n282), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n367), .A2(new_n352), .B1(G33), .B2(G87), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n295), .B(new_n331), .C1(new_n368), .C2(new_n289), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G169), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n328), .A2(G179), .A3(new_n331), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(KEYINPUT81), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n341), .A2(new_n366), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT18), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n328), .A2(G190), .A3(new_n331), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n369), .A2(G200), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n362), .A2(new_n375), .A3(new_n365), .A4(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT17), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n362), .A2(new_n365), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n380), .A2(KEYINPUT17), .A3(new_n375), .A4(new_n376), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT18), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n341), .A2(new_n366), .A3(new_n372), .A4(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n374), .A2(new_n379), .A3(new_n381), .A4(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G238), .ZN(new_n385));
  OAI221_X1 g0185(.A(new_n280), .B1(new_n385), .B2(new_n282), .C1(new_n285), .C2(new_n329), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n386), .B(new_n290), .C1(G107), .C2(new_n280), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n289), .A2(new_n292), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n209), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n387), .A2(new_n295), .A3(new_n389), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n390), .A2(G179), .ZN(new_n391));
  XOR2_X1   g0191(.A(KEYINPUT15), .B(G87), .Z(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n393), .A2(new_n262), .ZN(new_n394));
  INV_X1    g0194(.A(G77), .ZN(new_n395));
  OAI22_X1  g0195(.A1(new_n263), .A2(new_n261), .B1(new_n225), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n266), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n273), .A2(new_n395), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n397), .B(new_n398), .C1(new_n395), .C2(new_n277), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n390), .A2(new_n309), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n391), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n312), .A2(new_n384), .A3(new_n402), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n262), .A2(new_n395), .B1(new_n225), .B2(G68), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n404), .B(KEYINPUT77), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n201), .B2(new_n261), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT11), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n406), .A2(new_n407), .A3(new_n266), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n407), .B1(new_n406), .B2(new_n266), .ZN(new_n409));
  OR2_X1    g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OR2_X1    g0210(.A1(new_n277), .A2(new_n203), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n275), .A2(G68), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT12), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g0214(.A(new_n414), .B(KEYINPUT78), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n413), .B2(new_n412), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n410), .A2(new_n411), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n212), .B1(new_n317), .B2(new_n318), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n329), .A2(new_n282), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n280), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G33), .A2(G97), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n289), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n295), .B1(new_n296), .B2(new_n385), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT13), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT74), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT13), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n294), .B1(new_n388), .B2(G238), .ZN(new_n428));
  INV_X1    g0228(.A(new_n422), .ZN(new_n429));
  INV_X1    g0229(.A(new_n420), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n285), .B2(new_n212), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n429), .B1(new_n431), .B2(new_n280), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n427), .B(new_n428), .C1(new_n432), .C2(new_n289), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n425), .A2(new_n426), .A3(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n423), .A2(new_n424), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n435), .A2(KEYINPUT74), .A3(new_n427), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(G169), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT14), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n425), .A2(G179), .A3(new_n433), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT14), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n434), .A2(new_n436), .A3(new_n440), .A4(G169), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n438), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT79), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n438), .A2(KEYINPUT79), .A3(new_n439), .A4(new_n441), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n418), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n434), .A2(G200), .A3(new_n436), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT75), .ZN(new_n448));
  XNOR2_X1  g0248(.A(new_n447), .B(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n425), .A2(G190), .A3(new_n433), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT76), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(new_n418), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n446), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n399), .B1(G200), .B2(new_n390), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(new_n298), .B2(new_n390), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n403), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n275), .B(new_n276), .C1(G1), .C2(new_n265), .ZN(new_n459));
  INV_X1    g0259(.A(G107), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n357), .A2(new_n334), .A3(new_n225), .A4(G87), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT22), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT23), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n464), .B1(new_n225), .B2(G107), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n460), .A2(KEYINPUT23), .A3(G20), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n462), .A2(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G87), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n463), .A2(new_n468), .A3(G20), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n335), .A2(new_n322), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n225), .A2(G33), .A3(G116), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n467), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT88), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT88), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n467), .A2(new_n474), .A3(new_n470), .A4(new_n471), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n473), .A2(KEYINPUT24), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT24), .B1(new_n473), .B2(new_n475), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n461), .B1(new_n478), .B2(new_n266), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n273), .A2(new_n460), .ZN(new_n480));
  XNOR2_X1  g0280(.A(new_n480), .B(KEYINPUT89), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT25), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT89), .ZN(new_n483));
  XNOR2_X1  g0283(.A(new_n480), .B(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT25), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g0287(.A(KEYINPUT90), .B(G294), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G33), .ZN(new_n489));
  AND2_X1   g0289(.A1(G257), .A2(G1698), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n490), .B1(new_n319), .B2(G250), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n489), .B1(new_n491), .B2(new_n326), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT91), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT91), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n494), .B(new_n489), .C1(new_n491), .C2(new_n326), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n493), .A2(new_n495), .A3(new_n290), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n288), .A2(KEYINPUT5), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(G45), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n499), .A2(G1), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n288), .A2(KEYINPUT5), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n498), .A2(G274), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT5), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n268), .B(G45), .C1(new_n503), .C2(G41), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n504), .A2(new_n497), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(new_n290), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G264), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n496), .A2(new_n502), .A3(new_n507), .ZN(new_n508));
  OR2_X1    g0308(.A1(new_n508), .A2(new_n298), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(G200), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n479), .A2(new_n487), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT4), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n319), .A2(G244), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n326), .B2(new_n513), .ZN(new_n514));
  OAI211_X1 g0314(.A(KEYINPUT4), .B(G244), .C1(new_n283), .C2(new_n284), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G250), .A2(G1698), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n280), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G283), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n514), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n290), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n289), .B(G257), .C1(new_n504), .C2(new_n497), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n522), .A2(new_n502), .A3(KEYINPUT82), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(KEYINPUT82), .B1(new_n522), .B2(new_n502), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT83), .B1(new_n524), .B2(new_n525), .ZN(new_n529));
  INV_X1    g0329(.A(new_n525), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT83), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n531), .A3(new_n523), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n529), .A2(new_n532), .A3(new_n521), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n528), .A2(G190), .B1(new_n533), .B2(G200), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n356), .A2(new_n359), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G107), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n260), .A2(G77), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n460), .A2(KEYINPUT6), .A3(G97), .ZN(new_n538));
  INV_X1    g0338(.A(G97), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(new_n460), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n540), .A2(new_n206), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n538), .B1(new_n541), .B2(KEYINPUT6), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G20), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n536), .A2(new_n537), .A3(new_n543), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n544), .A2(new_n266), .B1(new_n539), .B2(new_n273), .ZN(new_n545));
  OR2_X1    g0345(.A1(new_n459), .A2(new_n539), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n545), .A2(new_n546), .B1(new_n527), .B2(new_n309), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n529), .A2(new_n532), .A3(new_n521), .A4(new_n339), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n534), .A2(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n519), .B(new_n225), .C1(G33), .C2(new_n539), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n551), .B(new_n266), .C1(new_n225), .C2(G116), .ZN(new_n552));
  XOR2_X1   g0352(.A(new_n552), .B(KEYINPUT20), .Z(new_n553));
  INV_X1    g0353(.A(G116), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n273), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n553), .B(new_n555), .C1(new_n554), .C2(new_n459), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n358), .A2(G303), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n319), .A2(G257), .B1(G264), .B2(G1698), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n557), .B1(new_n558), .B2(new_n326), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT86), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT86), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n561), .B(new_n557), .C1(new_n558), .C2(new_n326), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n560), .A2(new_n562), .A3(new_n290), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n506), .A2(G270), .B1(G274), .B2(new_n505), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n556), .B1(new_n565), .B2(G200), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n298), .B2(new_n565), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n511), .A2(new_n550), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n500), .A2(G274), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n289), .B(G250), .C1(G1), .C2(new_n499), .ZN(new_n570));
  OAI21_X1  g0370(.A(G238), .B1(new_n283), .B2(new_n284), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G244), .A2(G1698), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n352), .A2(new_n573), .B1(G33), .B2(G116), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n569), .B(new_n570), .C1(new_n574), .C2(new_n289), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT84), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n319), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n577));
  OAI22_X1  g0377(.A1(new_n577), .A2(new_n326), .B1(new_n265), .B2(new_n554), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n290), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT84), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n579), .A2(new_n580), .A3(new_n569), .A4(new_n570), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n576), .A2(new_n581), .A3(G200), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n352), .A2(new_n225), .A3(G68), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT19), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n225), .B1(new_n422), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(G87), .B2(new_n207), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n584), .B1(new_n262), .B2(new_n539), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n583), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n266), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n273), .A2(new_n393), .ZN(new_n590));
  OR2_X1    g0390(.A1(new_n459), .A2(new_n468), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n582), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT85), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n576), .A2(new_n581), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G190), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n582), .A2(new_n593), .A3(KEYINPUT85), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n596), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n597), .A2(new_n339), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n589), .B(new_n590), .C1(new_n393), .C2(new_n459), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n601), .B(new_n602), .C1(G169), .C2(new_n597), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT21), .ZN(new_n605));
  AOI211_X1 g0405(.A(new_n605), .B(new_n309), .C1(new_n563), .C2(new_n564), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n563), .A2(G179), .A3(new_n564), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n556), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n565), .A2(G169), .A3(new_n556), .ZN(new_n609));
  XNOR2_X1  g0409(.A(KEYINPUT87), .B(KEYINPUT21), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n473), .A2(new_n475), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT24), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n473), .A2(KEYINPUT24), .A3(new_n475), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(new_n266), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n461), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n616), .A2(new_n617), .A3(new_n487), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n508), .A2(new_n309), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(G179), .B2(new_n508), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n608), .B(new_n611), .C1(new_n618), .C2(new_n620), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n568), .A2(new_n604), .A3(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n458), .A2(new_n622), .ZN(G372));
  NAND2_X1  g0423(.A1(new_n381), .A2(new_n379), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n444), .A2(new_n445), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n417), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n453), .A2(new_n402), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n624), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n366), .B1(new_n332), .B2(new_n340), .ZN(new_n629));
  XNOR2_X1  g0429(.A(new_n629), .B(new_n382), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n308), .B(new_n307), .C1(new_n628), .C2(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n632), .A2(new_n311), .ZN(new_n633));
  INV_X1    g0433(.A(G200), .ZN(new_n634));
  INV_X1    g0434(.A(new_n575), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n593), .B(KEYINPUT92), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT92), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n635), .A2(new_n634), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n637), .B1(new_n638), .B2(new_n592), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n636), .A2(new_n598), .A3(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n621), .A2(new_n550), .A3(new_n511), .A4(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n548), .A2(new_n549), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n600), .A2(new_n643), .A3(new_n603), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT26), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n601), .B(new_n602), .C1(G169), .C2(new_n635), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT26), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n640), .A2(new_n643), .A3(new_n646), .A4(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n641), .A2(new_n645), .A3(new_n646), .A4(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n458), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n633), .A2(new_n650), .ZN(G369));
  NOR2_X1   g0451(.A1(new_n618), .A2(new_n620), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n225), .A2(G13), .ZN(new_n653));
  OR3_X1    g0453(.A1(new_n653), .A2(KEYINPUT27), .A3(G1), .ZN(new_n654));
  OAI21_X1  g0454(.A(KEYINPUT27), .B1(new_n653), .B2(G1), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(G213), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n618), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n652), .B1(new_n660), .B2(new_n511), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n618), .A2(new_n620), .A3(new_n658), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n608), .A2(new_n611), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n659), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n556), .A2(new_n658), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n664), .A2(new_n668), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(new_n567), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(G330), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n662), .B1(new_n663), .B2(new_n666), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(G399));
  INV_X1    g0476(.A(new_n235), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(G41), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(new_n268), .ZN(new_n679));
  NOR3_X1   g0479(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n680));
  INV_X1    g0480(.A(new_n227), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n679), .A2(new_n680), .B1(new_n681), .B2(new_n678), .ZN(new_n682));
  XOR2_X1   g0482(.A(new_n682), .B(KEYINPUT28), .Z(new_n683));
  AND2_X1   g0483(.A1(new_n641), .A2(new_n646), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n640), .A2(new_n643), .A3(new_n646), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(KEYINPUT26), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n600), .A2(new_n647), .A3(new_n643), .A4(new_n603), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n658), .B1(new_n684), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n690), .A2(KEYINPUT95), .A3(KEYINPUT29), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT95), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n649), .A2(new_n659), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT29), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AOI211_X1 g0495(.A(new_n694), .B(new_n658), .C1(new_n684), .C2(new_n689), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n691), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT31), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n496), .A2(new_n521), .A3(new_n507), .A4(new_n526), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n700), .A2(new_n607), .A3(KEYINPUT30), .A4(new_n597), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT93), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n563), .A2(G179), .A3(new_n564), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT93), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n704), .A2(new_n705), .A3(KEYINPUT30), .A4(new_n597), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n597), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n708), .A2(new_n703), .A3(new_n699), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT94), .B1(new_n709), .B2(KEYINPUT30), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n635), .A2(G179), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n711), .A2(new_n508), .A3(new_n533), .A4(new_n565), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n704), .A2(new_n597), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT94), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT30), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n707), .A2(new_n710), .A3(new_n712), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n658), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n698), .A2(new_n718), .B1(new_n622), .B2(new_n659), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n707), .B(new_n712), .C1(KEYINPUT30), .C2(new_n709), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n720), .A2(KEYINPUT31), .A3(new_n658), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n672), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n697), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n683), .B1(new_n724), .B2(G1), .ZN(G364));
  XNOR2_X1  g0525(.A(new_n653), .B(KEYINPUT96), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G45), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G1), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n678), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n671), .A2(new_n672), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n673), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G13), .A2(G33), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G20), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n730), .B1(new_n671), .B2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n224), .B1(G20), .B2(new_n309), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n225), .A2(new_n298), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n339), .A2(new_n634), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G326), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n339), .A2(G200), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G322), .ZN(new_n744));
  OAI22_X1  g0544(.A1(new_n740), .A2(new_n741), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n634), .A2(G179), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT99), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n225), .A2(G190), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G179), .A2(G200), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n225), .B1(new_n751), .B2(G190), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n750), .A2(G283), .B1(new_n488), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n747), .A2(new_n738), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G303), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n739), .A2(new_n748), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(KEYINPUT33), .B(G317), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n748), .A2(new_n751), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n759), .A2(new_n760), .B1(new_n762), .B2(G329), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n754), .A2(new_n358), .A3(new_n757), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n748), .A2(new_n742), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n745), .B(new_n764), .C1(G311), .C2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n756), .A2(G87), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(new_n201), .B2(new_n740), .ZN(new_n769));
  INV_X1    g0569(.A(G159), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n761), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT32), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n358), .B1(new_n766), .B2(G77), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n772), .B(new_n773), .C1(new_n460), .C2(new_n749), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n752), .A2(new_n539), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n202), .A2(new_n743), .B1(new_n758), .B2(new_n203), .ZN(new_n776));
  NOR4_X1   g0576(.A1(new_n769), .A2(new_n774), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n737), .B1(new_n767), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n677), .A2(new_n358), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n779), .A2(G355), .B1(new_n554), .B2(new_n677), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n235), .A2(new_n326), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT98), .Z(new_n782));
  NAND2_X1  g0582(.A1(new_n228), .A2(new_n499), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n256), .A2(G45), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT97), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n780), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n735), .A2(new_n737), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n736), .A2(new_n778), .A3(new_n789), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n732), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(G396));
  NAND2_X1  g0592(.A1(new_n399), .A2(new_n658), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n457), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n401), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n401), .A2(new_n658), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT101), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(new_n649), .B2(new_n659), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT102), .ZN(new_n801));
  INV_X1    g0601(.A(new_n798), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n649), .A2(new_n659), .A3(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OR3_X1    g0604(.A1(new_n801), .A2(new_n723), .A3(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n723), .B1(new_n801), .B2(new_n804), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n805), .A2(new_n730), .A3(new_n806), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G283), .A2(new_n759), .B1(new_n766), .B2(G116), .ZN(new_n808));
  INV_X1    g0608(.A(G294), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n808), .B1(new_n809), .B2(new_n743), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n750), .A2(G87), .ZN(new_n811));
  INV_X1    g0611(.A(G311), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n812), .B2(new_n761), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT100), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n775), .A2(new_n280), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n814), .B(new_n815), .C1(new_n460), .C2(new_n755), .ZN(new_n816));
  INV_X1    g0616(.A(new_n740), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n810), .B(new_n816), .C1(G303), .C2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n743), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G143), .A2(new_n819), .B1(new_n759), .B2(G150), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n817), .A2(G137), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n820), .B(new_n821), .C1(new_n770), .C2(new_n765), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT34), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n202), .B2(new_n752), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n822), .A2(new_n823), .B1(new_n201), .B2(new_n755), .ZN(new_n826));
  INV_X1    g0626(.A(G132), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n761), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n352), .B1(new_n749), .B2(new_n203), .ZN(new_n829));
  NOR4_X1   g0629(.A1(new_n825), .A2(new_n826), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n737), .B1(new_n818), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n798), .A2(new_n733), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n737), .A2(new_n733), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n395), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n831), .A2(new_n729), .A3(new_n832), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n807), .A2(new_n835), .ZN(G384));
  NAND2_X1  g0636(.A1(new_n417), .A2(new_n658), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n455), .A2(new_n837), .B1(new_n446), .B2(new_n658), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(new_n803), .B2(new_n797), .ZN(new_n839));
  INV_X1    g0639(.A(new_n656), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n347), .B1(new_n350), .B2(new_n353), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n841), .A2(new_n355), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n354), .A2(new_n266), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n365), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n384), .A2(new_n840), .A3(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT37), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n366), .A2(new_n840), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n373), .A2(new_n846), .A3(new_n377), .A4(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n370), .A2(new_n371), .A3(new_n656), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n850), .A2(new_n377), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n848), .B1(new_n851), .B2(new_n846), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n845), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT38), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n845), .A2(KEYINPUT38), .A3(new_n852), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n839), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n631), .A2(new_n656), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT104), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n629), .A2(new_n377), .A3(new_n847), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT106), .ZN(new_n864));
  AND3_X1   g0664(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT37), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n864), .B1(new_n863), .B2(KEYINPUT37), .ZN(new_n866));
  INV_X1    g0666(.A(new_n848), .ZN(new_n867));
  NOR3_X1   g0667(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n624), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n847), .B1(new_n630), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n854), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT39), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n871), .A2(new_n872), .A3(new_n856), .ZN(new_n873));
  INV_X1    g0673(.A(new_n856), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT38), .B1(new_n845), .B2(new_n852), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT39), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n446), .A2(KEYINPUT105), .A3(new_n659), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT105), .B1(new_n446), .B2(new_n659), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n858), .A2(KEYINPUT104), .A3(new_n859), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n862), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n691), .B(new_n458), .C1(new_n695), .C2(new_n696), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n633), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n885), .B(new_n887), .Z(new_n888));
  NAND2_X1  g0688(.A1(new_n718), .A2(new_n698), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n568), .A2(new_n604), .ZN(new_n890));
  INV_X1    g0690(.A(new_n621), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n890), .A2(new_n891), .A3(new_n659), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n717), .A2(KEYINPUT31), .A3(new_n658), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n889), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n626), .A2(new_n453), .A3(new_n837), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n446), .A2(new_n658), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n798), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n894), .A2(new_n857), .A3(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT40), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n871), .A2(new_n856), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n901), .A2(new_n894), .A3(KEYINPUT40), .A4(new_n897), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n900), .A2(G330), .A3(new_n902), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n458), .A2(new_n894), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(G330), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n900), .A2(new_n904), .A3(new_n902), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n888), .B(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n268), .B2(new_n726), .ZN(new_n910));
  OAI211_X1 g0710(.A(G116), .B(new_n226), .C1(new_n542), .C2(KEYINPUT35), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n911), .B(KEYINPUT103), .Z(new_n912));
  NAND2_X1  g0712(.A1(new_n542), .A2(KEYINPUT35), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT36), .ZN(new_n915));
  OAI21_X1  g0715(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n916), .A2(new_n227), .B1(G50), .B2(new_n203), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(G1), .A3(new_n231), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n910), .A2(new_n915), .A3(new_n918), .ZN(G367));
  INV_X1    g0719(.A(new_n675), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n550), .B1(new_n547), .B2(new_n659), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT42), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n920), .B(new_n922), .C1(new_n923), .C2(new_n662), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n663), .A2(new_n666), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT42), .B1(new_n925), .B2(new_n921), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n924), .B(new_n926), .C1(new_n642), .C2(new_n658), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n592), .A2(new_n658), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n640), .A2(new_n646), .A3(new_n928), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n929), .A2(KEYINPUT107), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(KEYINPUT107), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n930), .B(new_n931), .C1(new_n646), .C2(new_n928), .ZN(new_n932));
  XNOR2_X1  g0732(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n933));
  OR3_X1    g0733(.A1(new_n927), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n927), .B(new_n935), .C1(new_n932), .C2(new_n933), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n643), .A2(new_n658), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n921), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n937), .B1(new_n674), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n674), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n934), .A2(new_n942), .A3(new_n939), .A4(new_n936), .ZN(new_n943));
  XNOR2_X1  g0743(.A(KEYINPUT109), .B(KEYINPUT41), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n678), .B(new_n944), .Z(new_n945));
  NAND2_X1  g0745(.A1(new_n667), .A2(new_n673), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n674), .A2(new_n925), .A3(new_n946), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n724), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n675), .A2(new_n939), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT45), .ZN(new_n950));
  XOR2_X1   g0750(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n951));
  NAND3_X1  g0751(.A1(new_n920), .A2(new_n940), .A3(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n951), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n675), .B2(new_n939), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  OR3_X1    g0755(.A1(new_n950), .A2(new_n942), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n948), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n945), .B1(new_n957), .B2(new_n724), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n941), .B(new_n943), .C1(new_n958), .C2(new_n728), .ZN(new_n959));
  INV_X1    g0759(.A(new_n932), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n735), .ZN(new_n961));
  INV_X1    g0761(.A(new_n782), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n788), .B1(new_n235), .B2(new_n393), .C1(new_n962), .C2(new_n249), .ZN(new_n963));
  INV_X1    g0763(.A(G143), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n740), .A2(new_n964), .B1(new_n765), .B2(new_n201), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n749), .A2(new_n395), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n965), .B(new_n966), .C1(G137), .C2(new_n762), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n752), .A2(new_n203), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n358), .B(new_n968), .C1(new_n756), .C2(G58), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n970), .B1(new_n259), .B2(new_n743), .C1(new_n770), .C2(new_n758), .ZN(new_n971));
  INV_X1    g0771(.A(G283), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n765), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(G317), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n974), .A2(new_n761), .B1(new_n752), .B2(new_n460), .ZN(new_n975));
  OR3_X1    g0775(.A1(new_n755), .A2(KEYINPUT46), .A3(new_n554), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT46), .B1(new_n755), .B2(new_n554), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n750), .A2(G97), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n352), .B1(new_n488), .B2(new_n759), .ZN(new_n980));
  AOI22_X1  g0780(.A1(G311), .A2(new_n817), .B1(new_n819), .B2(G303), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n978), .A2(new_n979), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n971), .B1(new_n973), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT47), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n737), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n961), .A2(new_n729), .A3(new_n963), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n959), .A2(new_n986), .ZN(G387));
  NAND2_X1  g0787(.A1(new_n753), .A2(new_n392), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n201), .B2(new_n743), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n326), .B(new_n989), .C1(G150), .C2(new_n762), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n756), .A2(G77), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n363), .A2(new_n759), .B1(new_n766), .B2(G68), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n750), .A2(G97), .B1(G159), .B2(new_n817), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n990), .A2(new_n991), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  AOI22_X1  g0794(.A1(G311), .A2(new_n759), .B1(new_n819), .B2(G317), .ZN(new_n995));
  INV_X1    g0795(.A(G303), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n995), .B1(new_n996), .B2(new_n765), .C1(new_n744), .C2(new_n740), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT48), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n756), .A2(new_n488), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n998), .B(new_n999), .C1(new_n972), .C2(new_n752), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT49), .Z(new_n1001));
  OAI221_X1 g0801(.A(new_n326), .B1(new_n741), .B2(new_n761), .C1(new_n749), .C2(new_n554), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n994), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n737), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n735), .B1(new_n661), .B2(new_n662), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n245), .A2(G45), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT111), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n263), .A2(G50), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT50), .ZN(new_n1010));
  AOI21_X1  g0810(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1010), .A2(new_n680), .A3(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1008), .A2(new_n782), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n779), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1013), .B1(G107), .B2(new_n235), .C1(new_n680), .C2(new_n1014), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n730), .B(new_n1006), .C1(new_n788), .C2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(new_n947), .B2(new_n728), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n678), .B1(new_n724), .B2(new_n947), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1017), .B1(new_n948), .B2(new_n1018), .ZN(G393));
  OAI21_X1  g0819(.A(new_n942), .B1(new_n950), .B2(new_n955), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n956), .A2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n678), .B(new_n957), .C1(new_n1021), .C2(new_n948), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n940), .A2(new_n735), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n756), .A2(G283), .B1(G322), .B2(new_n762), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1025), .A2(KEYINPUT114), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n740), .A2(new_n974), .B1(new_n743), .B2(new_n812), .ZN(new_n1027));
  XOR2_X1   g0827(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n1028));
  XNOR2_X1  g0828(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n1025), .B2(KEYINPUT114), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n752), .A2(new_n554), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n750), .A2(G107), .B1(G294), .B2(new_n766), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1032), .B(new_n358), .C1(new_n996), .C2(new_n758), .ZN(new_n1033));
  NOR4_X1   g0833(.A1(new_n1026), .A2(new_n1030), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n759), .A2(G50), .B1(new_n753), .B2(G77), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1035), .B(new_n352), .C1(new_n263), .C2(new_n765), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n740), .A2(new_n259), .B1(new_n743), .B2(new_n770), .ZN(new_n1037));
  XOR2_X1   g0837(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n1038));
  XNOR2_X1  g0838(.A(new_n1037), .B(new_n1038), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1039), .B(new_n811), .C1(new_n203), .C2(new_n755), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1036), .B(new_n1040), .C1(G143), .C2(new_n762), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n737), .B1(new_n1034), .B2(new_n1041), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n788), .B1(new_n539), .B2(new_n235), .C1(new_n962), .C2(new_n253), .ZN(new_n1043));
  AND4_X1   g0843(.A1(new_n729), .A2(new_n1023), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n1021), .B2(new_n728), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1022), .A2(new_n1045), .ZN(G390));
  NAND2_X1  g0846(.A1(new_n641), .A2(new_n646), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n659), .B(new_n795), .C1(new_n1047), .C2(new_n688), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n797), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n894), .A2(G330), .A3(new_n799), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n838), .A2(new_n1051), .B1(new_n722), .B2(new_n897), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n889), .A2(new_n892), .A3(new_n721), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1053), .A2(G330), .A3(new_n802), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n838), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n894), .A2(new_n897), .A3(G330), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n803), .A2(new_n797), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1050), .A2(new_n1052), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n886), .A2(new_n633), .A3(new_n905), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n876), .B(new_n873), .C1(new_n839), .C2(new_n882), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n838), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1049), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT115), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n879), .B2(new_n880), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT105), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n626), .B2(new_n658), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1067), .A2(KEYINPUT115), .A3(new_n878), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1063), .A2(new_n1069), .A3(new_n901), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n722), .A2(new_n897), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n1061), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1056), .B1(new_n1061), .B2(new_n1070), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n1059), .A2(new_n1060), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1051), .A2(new_n838), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1075), .A2(new_n1071), .A3(new_n1050), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n894), .A2(new_n897), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1077), .A2(G330), .B1(new_n1054), .B2(new_n838), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1058), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1076), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1056), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1058), .A2(new_n1062), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n877), .B1(new_n1082), .B2(new_n881), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n838), .B1(new_n1048), .B2(new_n797), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n901), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1081), .B1(new_n1083), .B2(new_n1087), .ZN(new_n1088));
  AND3_X1   g0888(.A1(new_n886), .A2(new_n633), .A3(new_n905), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1061), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1080), .A2(new_n1088), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1074), .A2(new_n678), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT116), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1074), .A2(new_n1091), .A3(KEYINPUT116), .A4(new_n678), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n730), .B1(new_n263), .B2(new_n833), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT117), .Z(new_n1098));
  AOI22_X1  g0898(.A1(new_n759), .A2(G137), .B1(new_n753), .B2(G159), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n827), .B2(new_n743), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n358), .B(new_n1100), .C1(G50), .C2(new_n750), .ZN(new_n1101));
  XOR2_X1   g0901(.A(KEYINPUT54), .B(G143), .Z(new_n1102));
  NAND2_X1  g0902(.A1(new_n766), .A2(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n817), .A2(G128), .B1(new_n762), .B2(G125), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n755), .A2(new_n259), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT53), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1101), .A2(new_n1103), .A3(new_n1104), .A4(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n761), .A2(new_n809), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n743), .A2(new_n554), .B1(new_n752), .B2(new_n395), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT118), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1110), .A2(new_n280), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n817), .A2(G283), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n758), .A2(new_n460), .B1(new_n765), .B2(new_n539), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n750), .B2(G68), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1111), .A2(new_n768), .A3(new_n1112), .A4(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1107), .B1(new_n1108), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1098), .B1(new_n1116), .B2(new_n737), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT119), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n877), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1118), .B1(new_n1119), .B2(new_n733), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1120), .B1(new_n1122), .B2(new_n728), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1096), .A2(new_n1123), .ZN(G378));
  INV_X1    g0924(.A(KEYINPUT122), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n903), .A2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n900), .A2(KEYINPUT122), .A3(G330), .A4(new_n902), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n312), .B(KEYINPUT121), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n278), .A2(new_n840), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1128), .B(new_n1129), .ZN(new_n1130));
  XOR2_X1   g0930(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1131));
  XNOR2_X1  g0931(.A(new_n1130), .B(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1126), .A2(new_n1127), .A3(new_n1132), .ZN(new_n1133));
  OR2_X1    g0933(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n903), .A2(new_n1134), .A3(new_n1125), .A4(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n885), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n885), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1139), .A2(new_n1133), .A3(new_n1136), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1089), .B1(new_n1121), .B2(new_n1059), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1138), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT57), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1138), .A2(new_n1140), .A3(new_n1141), .A4(KEYINPUT57), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1144), .A2(new_n678), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1138), .A2(new_n1140), .A3(new_n728), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n730), .B1(new_n1132), .B2(new_n733), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n750), .A2(G58), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT120), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1150), .A2(new_n288), .A3(new_n326), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n393), .A2(new_n765), .B1(new_n539), .B2(new_n758), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n991), .B1(new_n460), .B2(new_n743), .C1(new_n554), .C2(new_n740), .ZN(new_n1153));
  NOR4_X1   g0953(.A1(new_n1151), .A2(new_n968), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n972), .B2(new_n761), .ZN(new_n1155));
  XOR2_X1   g0955(.A(new_n1155), .B(KEYINPUT58), .Z(new_n1156));
  AOI21_X1  g0956(.A(G50), .B1(new_n326), .B2(new_n288), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(G33), .B2(G41), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n756), .A2(new_n1102), .B1(G137), .B2(new_n766), .ZN(new_n1159));
  INV_X1    g0959(.A(G125), .ZN(new_n1160));
  INV_X1    g0960(.A(G128), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n740), .A2(new_n1160), .B1(new_n743), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(G150), .B2(new_n753), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1159), .B(new_n1163), .C1(new_n827), .C2(new_n758), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT59), .ZN(new_n1165));
  AOI211_X1 g0965(.A(G33), .B(G41), .C1(new_n762), .C2(G124), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n770), .B2(new_n749), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1158), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n737), .B1(new_n1156), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n833), .A2(new_n201), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1148), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1147), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1146), .A2(new_n1172), .ZN(G375));
  NAND2_X1  g0973(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n945), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1080), .A2(new_n1089), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n838), .A2(new_n733), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n326), .B1(G150), .B2(new_n766), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n759), .A2(new_n1102), .B1(new_n753), .B2(G50), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n817), .A2(G132), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n819), .A2(G137), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1150), .B1(new_n1161), .B2(new_n761), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(G159), .C2(new_n756), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n817), .A2(G294), .B1(new_n762), .B2(G303), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n280), .B1(new_n759), .B2(G116), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n972), .C2(new_n743), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n988), .B1(new_n755), .B2(new_n539), .C1(new_n395), .C2(new_n749), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(G107), .C2(new_n766), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n737), .B1(new_n1185), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n833), .A2(new_n203), .ZN(new_n1192));
  AND4_X1   g0992(.A1(new_n729), .A2(new_n1178), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n1080), .B2(new_n728), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1177), .A2(new_n1194), .ZN(G381));
  AND2_X1   g0995(.A1(new_n1123), .A2(new_n1092), .ZN(new_n1196));
  AND3_X1   g0996(.A1(new_n1146), .A2(new_n1172), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(G384), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n959), .A2(new_n986), .A3(new_n1045), .A4(new_n1022), .ZN(new_n1200));
  OR3_X1    g1000(.A1(new_n1200), .A2(G396), .A3(G393), .ZN(new_n1201));
  NOR3_X1   g1001(.A1(new_n1199), .A2(new_n1201), .A3(G381), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(G407));
  NAND2_X1  g1003(.A1(new_n1197), .A2(new_n657), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(G213), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1202), .A2(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT123), .ZN(G409));
  INV_X1    g1007(.A(KEYINPUT61), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(G393), .B(new_n791), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1200), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n959), .A2(new_n986), .B1(new_n1045), .B2(new_n1022), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1209), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1211), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1209), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1213), .A2(new_n1200), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1212), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1146), .A2(G378), .A3(new_n1172), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1147), .B(new_n1171), .C1(new_n1142), .C2(new_n945), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n1196), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n657), .A2(G213), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT60), .ZN(new_n1223));
  OAI211_X1 g1023(.A(KEYINPUT125), .B(new_n1223), .C1(new_n1080), .C2(new_n1089), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1224), .A2(new_n678), .A3(new_n1176), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1223), .B1(new_n1174), .B2(KEYINPUT125), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1194), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1227), .A2(new_n1198), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1198), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT63), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1216), .B1(new_n1222), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT124), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1220), .A2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1217), .A2(KEYINPUT124), .A3(new_n1219), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n1221), .A3(new_n1236), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n657), .A2(G213), .A3(G2897), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1230), .B(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1231), .B1(new_n1237), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1230), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1235), .A2(new_n1221), .A3(new_n1242), .A4(new_n1236), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1208), .B(new_n1233), .C1(new_n1241), .C2(new_n1244), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1228), .A2(KEYINPUT62), .A3(new_n1229), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1220), .A2(new_n1221), .A3(new_n1246), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1247), .B1(new_n1243), .B2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1208), .B1(new_n1222), .B2(new_n1239), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1216), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1245), .A2(new_n1251), .ZN(G405));
  INV_X1    g1052(.A(KEYINPUT127), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1230), .A2(new_n1253), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1216), .B(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(G375), .A2(new_n1196), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1256), .A2(new_n1217), .B1(new_n1253), .B2(new_n1230), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1255), .B(new_n1257), .ZN(G402));
endmodule


