//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n561, new_n562, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n582,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n639, new_n640, new_n643, new_n644, new_n646, new_n647,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1247, new_n1248, new_n1249, new_n1250;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n460), .A2(new_n462), .A3(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n459), .A2(KEYINPUT65), .A3(G2104), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n467), .A2(new_n462), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n470), .B1(new_n461), .B2(KEYINPUT3), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n468), .A2(G137), .A3(new_n469), .A4(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n469), .A2(G101), .A3(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n466), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  OAI21_X1  g050(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(G112), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(G2105), .ZN(new_n478));
  AND4_X1   g053(.A1(new_n469), .A2(new_n471), .A3(new_n467), .A4(new_n462), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n481));
  NAND4_X1  g056(.A1(new_n468), .A2(new_n481), .A3(G2105), .A4(new_n471), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n471), .A2(new_n467), .A3(G2105), .A4(new_n462), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT66), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  AOI211_X1 g061(.A(new_n478), .B(new_n480), .C1(new_n486), .C2(G124), .ZN(G162));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n471), .A2(new_n467), .A3(new_n489), .A4(new_n462), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n460), .A2(new_n462), .ZN(new_n491));
  NOR3_X1   g066(.A1(new_n488), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n492));
  AOI22_X1  g067(.A1(new_n490), .A2(KEYINPUT4), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(G114), .B2(new_n469), .ZN(new_n496));
  INV_X1    g071(.A(G126), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n483), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n493), .A2(new_n498), .ZN(G164));
  OR2_X1    g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  OR2_X1    g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT67), .B1(new_n506), .B2(G651), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT67), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(new_n504), .A3(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n510), .A2(G88), .A3(new_n502), .A4(new_n512), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n510), .A2(G50), .A3(G543), .A4(new_n512), .ZN(new_n514));
  AND3_X1   g089(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT68), .ZN(new_n515));
  AOI21_X1  g090(.A(KEYINPUT68), .B1(new_n513), .B2(new_n514), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n505), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(G166));
  INV_X1    g093(.A(G51), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n508), .B1(KEYINPUT6), .B2(new_n504), .ZN(new_n520));
  NOR3_X1   g095(.A1(new_n506), .A2(KEYINPUT67), .A3(G651), .ZN(new_n521));
  OAI211_X1 g096(.A(G543), .B(new_n512), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT69), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n511), .B1(new_n507), .B2(new_n509), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n525), .A2(KEYINPUT69), .A3(G543), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n519), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n525), .A2(G89), .A3(new_n502), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT7), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n531), .A2(KEYINPUT70), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(KEYINPUT70), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT70), .B(KEYINPUT7), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(new_n529), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n502), .A2(G63), .A3(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n528), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n527), .A2(new_n539), .ZN(G168));
  XNOR2_X1  g115(.A(KEYINPUT71), .B(G52), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n541), .B1(new_n524), .B2(new_n526), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n525), .A2(G90), .A3(new_n502), .ZN(new_n543));
  INV_X1    g118(.A(G64), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n544), .B1(new_n500), .B2(new_n501), .ZN(new_n545));
  AND2_X1   g120(.A1(G77), .A2(G543), .ZN(new_n546));
  OAI21_X1  g121(.A(G651), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n542), .A2(new_n548), .ZN(G171));
  INV_X1    g124(.A(G56), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n550), .B1(new_n500), .B2(new_n501), .ZN(new_n551));
  AND2_X1   g126(.A1(G68), .A2(G543), .ZN(new_n552));
  OAI21_X1  g127(.A(G651), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g128(.A(KEYINPUT72), .B(G81), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n510), .A2(new_n502), .A3(new_n512), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n524), .A2(new_n526), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n556), .B1(new_n557), .B2(G43), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  NAND3_X1  g138(.A1(new_n525), .A2(G53), .A3(G543), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(KEYINPUT9), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  AND2_X1   g143(.A1(KEYINPUT5), .A2(G543), .ZN(new_n569));
  NOR2_X1   g144(.A1(KEYINPUT5), .A2(G543), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n568), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G651), .ZN(new_n574));
  INV_X1    g149(.A(G91), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n510), .A2(new_n502), .A3(new_n512), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n567), .A2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  INV_X1    g155(.A(G168), .ZN(G286));
  NAND2_X1  g156(.A1(new_n517), .A2(KEYINPUT73), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT73), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n583), .B(new_n505), .C1(new_n515), .C2(new_n516), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n582), .A2(new_n584), .ZN(G303));
  NAND3_X1  g160(.A1(new_n525), .A2(G49), .A3(G543), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n525), .A2(G87), .A3(new_n502), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(KEYINPUT74), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT74), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G288));
  NAND4_X1  g170(.A1(new_n510), .A2(G86), .A3(new_n502), .A4(new_n512), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n510), .A2(G48), .A3(G543), .A4(new_n512), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(G73), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(G61), .B1(new_n569), .B2(new_n570), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT75), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI211_X1 g178(.A(KEYINPUT75), .B(G61), .C1(new_n569), .C2(new_n570), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n504), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT76), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n598), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(G61), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(new_n500), .B2(new_n501), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n599), .B1(new_n609), .B2(KEYINPUT75), .ZN(new_n610));
  INV_X1    g185(.A(new_n604), .ZN(new_n611));
  OAI21_X1  g186(.A(G651), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(KEYINPUT76), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n607), .A2(new_n613), .ZN(G305));
  NAND2_X1  g189(.A1(G72), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G60), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n571), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G651), .ZN(new_n618));
  INV_X1    g193(.A(G85), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n576), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(G47), .B2(new_n557), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(G290));
  NAND2_X1  g197(.A1(G301), .A2(G868), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT77), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n624), .A2(G66), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(G66), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n502), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(G79), .A2(G543), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n504), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT10), .ZN(new_n630));
  INV_X1    g205(.A(G92), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n576), .B2(new_n631), .ZN(new_n632));
  NAND4_X1  g207(.A1(new_n525), .A2(KEYINPUT10), .A3(G92), .A4(new_n502), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n629), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n557), .A2(G54), .ZN(new_n635));
  AND2_X1   g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n623), .B1(new_n636), .B2(G868), .ZN(G321));
  XOR2_X1   g212(.A(G321), .B(KEYINPUT78), .Z(G284));
  NAND2_X1  g213(.A1(G286), .A2(G868), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n577), .B1(new_n565), .B2(new_n566), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(G868), .B2(new_n640), .ZN(G297));
  OAI21_X1  g216(.A(new_n639), .B1(G868), .B2(new_n640), .ZN(G280));
  INV_X1    g217(.A(G559), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n636), .B1(new_n643), .B2(G860), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT79), .ZN(G148));
  NAND2_X1  g220(.A1(new_n636), .A2(new_n643), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(G868), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(G868), .B2(new_n558), .ZN(G323));
  XNOR2_X1  g223(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g224(.A1(new_n486), .A2(G123), .ZN(new_n650));
  OAI21_X1  g225(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n651));
  INV_X1    g226(.A(G111), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n651), .B1(new_n652), .B2(G2105), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n653), .B1(new_n479), .B2(G135), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n655), .A2(G2096), .ZN(new_n656));
  INV_X1    g231(.A(new_n491), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n469), .A2(G2104), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(KEYINPUT13), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n655), .A2(G2096), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n656), .A2(new_n663), .A3(new_n664), .ZN(G156));
  XOR2_X1   g240(.A(G2451), .B(G2454), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT16), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1341), .B(G1348), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT14), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2427), .B(G2438), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2430), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT15), .B(G2435), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n670), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(new_n673), .B2(new_n672), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n669), .B(new_n675), .Z(new_n676));
  XNOR2_X1  g251(.A(G2443), .B(G2446), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  AND3_X1   g254(.A1(new_n678), .A2(G14), .A3(new_n679), .ZN(G401));
  INV_X1    g255(.A(KEYINPUT18), .ZN(new_n681));
  XOR2_X1   g256(.A(G2084), .B(G2090), .Z(new_n682));
  XNOR2_X1  g257(.A(G2067), .B(G2678), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(KEYINPUT17), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n682), .A2(new_n683), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n681), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G2100), .ZN(new_n688));
  XOR2_X1   g263(.A(G2072), .B(G2078), .Z(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n684), .B2(KEYINPUT18), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G2096), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n688), .B(new_n691), .ZN(G227));
  XNOR2_X1  g267(.A(G1961), .B(G1966), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT81), .ZN(new_n694));
  XOR2_X1   g269(.A(G1956), .B(G2474), .Z(new_n695));
  OR2_X1    g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1971), .B(G1976), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT19), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n694), .A2(new_n695), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n696), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n698), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT20), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR3_X1   g278(.A1(new_n699), .A2(KEYINPUT20), .A3(new_n698), .ZN(new_n704));
  OAI221_X1 g279(.A(new_n700), .B1(new_n698), .B2(new_n696), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT82), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n705), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1991), .B(G1996), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1981), .B(G1986), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n710), .A2(new_n712), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(G229));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G33), .ZN(new_n717));
  NAND2_X1  g292(.A1(G115), .A2(G2104), .ZN(new_n718));
  INV_X1    g293(.A(G127), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n657), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n469), .B1(new_n720), .B2(KEYINPUT92), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(KEYINPUT92), .B2(new_n720), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT91), .B(KEYINPUT25), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G139), .B2(new_n479), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n717), .B1(new_n728), .B2(new_n716), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G2072), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT85), .B(G16), .Z(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n732), .A2(G19), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n558), .B2(new_n732), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G1341), .ZN(new_n735));
  INV_X1    g310(.A(G16), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G21), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G168), .B2(new_n736), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT94), .B(G1966), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n738), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n716), .A2(G27), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G164), .B2(new_n716), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2078), .ZN(new_n744));
  NOR4_X1   g319(.A1(new_n730), .A2(new_n735), .A3(new_n741), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n731), .A2(G20), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT98), .B(KEYINPUT23), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G299), .B2(G16), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT99), .B(G1956), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(G171), .A2(new_n736), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G5), .B2(new_n736), .ZN(new_n753));
  INV_X1    g328(.A(G1961), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT30), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT95), .ZN(new_n757));
  AND3_X1   g332(.A1(new_n757), .A2(new_n756), .A3(G28), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n757), .B1(new_n756), .B2(G28), .ZN(new_n759));
  OAI221_X1 g334(.A(new_n716), .B1(new_n756), .B2(G28), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT31), .B(G11), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT24), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n763), .A2(G34), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(G34), .ZN(new_n766));
  AOI21_X1  g341(.A(G29), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n474), .B2(G29), .ZN(new_n768));
  INV_X1    g343(.A(G2084), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n762), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n655), .ZN(new_n771));
  INV_X1    g346(.A(new_n768), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n771), .A2(G29), .B1(new_n772), .B2(G2084), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n755), .A2(new_n770), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n479), .A2(G141), .ZN(new_n775));
  NAND3_X1  g350(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT26), .Z(new_n777));
  INV_X1    g352(.A(G105), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n775), .B(new_n777), .C1(new_n778), .C2(new_n658), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT93), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n486), .A2(new_n780), .A3(G129), .ZN(new_n781));
  INV_X1    g356(.A(G129), .ZN(new_n782));
  OAI21_X1  g357(.A(KEYINPUT93), .B1(new_n485), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n779), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n784), .A2(new_n716), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n716), .B2(G32), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT27), .B(G1996), .ZN(new_n787));
  AOI211_X1 g362(.A(new_n751), .B(new_n774), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n716), .A2(G26), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT28), .Z(new_n790));
  NAND3_X1  g365(.A1(new_n482), .A2(G128), .A3(new_n484), .ZN(new_n791));
  OAI21_X1  g366(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n792));
  INV_X1    g367(.A(G116), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n792), .B1(new_n793), .B2(G2105), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n479), .B2(G140), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT89), .ZN(new_n796));
  AND3_X1   g371(.A1(new_n791), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n796), .B1(new_n791), .B2(new_n795), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n790), .B1(new_n800), .B2(G29), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT90), .B(G2067), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n745), .A2(new_n788), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(G4), .A2(G16), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n636), .B2(G16), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT88), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1348), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n753), .A2(new_n754), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT96), .ZN(new_n810));
  NOR2_X1   g385(.A1(G29), .A2(G35), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G162), .B2(G29), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(G2090), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n810), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n814), .A2(new_n815), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n786), .B2(new_n787), .ZN(new_n818));
  NOR4_X1   g393(.A1(new_n804), .A2(new_n808), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n732), .A2(G22), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G166), .B2(new_n732), .ZN(new_n821));
  INV_X1    g396(.A(G1971), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n736), .A2(G23), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n590), .B2(new_n736), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT33), .B(G1976), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT32), .B(G1981), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT86), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n606), .B(G651), .C1(new_n610), .C2(new_n611), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n596), .A2(new_n597), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n603), .A2(new_n604), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n606), .B1(new_n833), .B2(G651), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(G16), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(G6), .B2(G16), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n827), .B1(new_n829), .B2(new_n837), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n823), .B(new_n838), .C1(new_n829), .C2(new_n837), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n839), .A2(KEYINPUT34), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(KEYINPUT34), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n486), .A2(G119), .ZN(new_n842));
  OAI21_X1  g417(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n843));
  INV_X1    g418(.A(G107), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n843), .B1(new_n844), .B2(G2105), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(new_n479), .B2(G131), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(G29), .ZN(new_n848));
  INV_X1    g423(.A(G25), .ZN(new_n849));
  OR3_X1    g424(.A1(new_n849), .A2(KEYINPUT83), .A3(G29), .ZN(new_n850));
  OAI21_X1  g425(.A(KEYINPUT83), .B1(new_n849), .B2(G29), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n848), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(KEYINPUT35), .B(G1991), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT84), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n852), .B(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n732), .A2(G24), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(new_n621), .B2(new_n732), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(G1986), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n840), .A2(new_n841), .A3(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT36), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n860), .A2(KEYINPUT87), .A3(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(KEYINPUT87), .B(KEYINPUT36), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n840), .A2(new_n841), .A3(new_n859), .A4(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n819), .A2(new_n862), .A3(new_n864), .ZN(G150));
  INV_X1    g440(.A(G150), .ZN(G311));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n867));
  INV_X1    g442(.A(G55), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(new_n524), .B2(new_n526), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n525), .A2(G93), .A3(new_n502), .ZN(new_n870));
  INV_X1    g445(.A(G67), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n871), .B1(new_n500), .B2(new_n501), .ZN(new_n872));
  AND2_X1   g447(.A1(G80), .A2(G543), .ZN(new_n873));
  OAI21_X1  g448(.A(G651), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n867), .B1(new_n869), .B2(new_n875), .ZN(new_n876));
  AND4_X1   g451(.A1(KEYINPUT69), .A2(new_n510), .A3(G543), .A4(new_n512), .ZN(new_n877));
  AOI21_X1  g452(.A(KEYINPUT69), .B1(new_n525), .B2(G543), .ZN(new_n878));
  OAI21_X1  g453(.A(G55), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n870), .A2(new_n874), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(KEYINPUT100), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n876), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(G860), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(KEYINPUT37), .Z(new_n884));
  NAND2_X1  g459(.A1(new_n636), .A2(G559), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT102), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT38), .ZN(new_n887));
  OAI21_X1  g462(.A(G43), .B1(new_n877), .B2(new_n878), .ZN(new_n888));
  INV_X1    g463(.A(new_n556), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n876), .A2(new_n881), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n879), .A2(new_n880), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT101), .B1(new_n892), .B2(new_n558), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n876), .A2(new_n881), .A3(KEYINPUT101), .A4(new_n890), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n887), .B(new_n896), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n897), .A2(KEYINPUT39), .ZN(new_n898));
  INV_X1    g473(.A(G860), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n899), .B1(new_n897), .B2(KEYINPUT39), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n884), .B1(new_n898), .B2(new_n900), .ZN(G145));
  INV_X1    g476(.A(KEYINPUT40), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n479), .A2(G142), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n469), .A2(G118), .ZN(new_n904));
  OAI21_X1  g479(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n906), .B1(G130), .B2(new_n486), .ZN(new_n907));
  XOR2_X1   g482(.A(new_n847), .B(new_n907), .Z(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(new_n661), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(G164), .B1(new_n797), .B2(new_n798), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n791), .A2(new_n795), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT89), .ZN(new_n913));
  INV_X1    g488(.A(G164), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n791), .A2(new_n796), .A3(new_n795), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n911), .A2(new_n916), .A3(new_n784), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n784), .B1(new_n911), .B2(new_n916), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT103), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n781), .A2(new_n783), .ZN(new_n920));
  INV_X1    g495(.A(new_n779), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n797), .A2(new_n798), .A3(G164), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n914), .B1(new_n913), .B2(new_n915), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT103), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n911), .A2(new_n916), .A3(new_n784), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n728), .B1(new_n919), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n728), .B1(new_n917), .B2(new_n918), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT104), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  AOI211_X1 g507(.A(KEYINPUT104), .B(new_n728), .C1(new_n919), .C2(new_n928), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n910), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n655), .B(new_n474), .ZN(new_n935));
  XOR2_X1   g510(.A(new_n935), .B(G162), .Z(new_n936));
  NAND2_X1  g511(.A1(new_n919), .A2(new_n928), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(new_n938), .A3(new_n727), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n939), .B(new_n909), .C1(new_n929), .C2(new_n931), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n934), .A2(new_n936), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(G37), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n936), .B1(new_n934), .B2(new_n940), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n902), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n934), .A2(new_n940), .ZN(new_n946));
  INV_X1    g521(.A(new_n936), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n948), .A2(KEYINPUT40), .A3(new_n942), .A4(new_n941), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n945), .A2(new_n949), .ZN(G395));
  XNOR2_X1  g525(.A(G305), .B(new_n621), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n517), .B(new_n590), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n951), .B(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n953), .B1(KEYINPUT105), .B2(KEYINPUT42), .ZN(new_n954));
  OR2_X1    g529(.A1(KEYINPUT105), .A2(KEYINPUT42), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n954), .B(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n634), .A2(new_n635), .ZN(new_n957));
  NOR2_X1   g532(.A1(G299), .A2(new_n957), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n567), .A2(new_n578), .B1(new_n634), .B2(new_n635), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT41), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n636), .A2(new_n640), .ZN(new_n961));
  NAND2_X1  g536(.A1(G299), .A2(new_n957), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT41), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n960), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n958), .A2(new_n959), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n896), .B(new_n646), .ZN(new_n967));
  MUX2_X1   g542(.A(new_n965), .B(new_n966), .S(new_n967), .Z(new_n968));
  AND2_X1   g543(.A1(new_n956), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n956), .A2(new_n968), .ZN(new_n970));
  OAI21_X1  g545(.A(G868), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n882), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n971), .B1(G868), .B2(new_n972), .ZN(G295));
  OAI21_X1  g548(.A(new_n971), .B1(G868), .B2(new_n972), .ZN(G331));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n976));
  OAI22_X1  g551(.A1(new_n527), .A2(new_n539), .B1(new_n542), .B2(new_n548), .ZN(new_n977));
  OAI21_X1  g552(.A(G51), .B1(new_n877), .B2(new_n878), .ZN(new_n978));
  INV_X1    g553(.A(new_n541), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n877), .B2(new_n878), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n528), .A2(new_n537), .A3(new_n538), .ZN(new_n981));
  INV_X1    g556(.A(new_n548), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n978), .A2(new_n980), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n977), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n894), .A2(new_n895), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT106), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n984), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n896), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n894), .A2(KEYINPUT106), .A3(new_n984), .A4(new_n895), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n987), .A2(new_n989), .A3(new_n966), .A4(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n985), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n984), .B1(new_n894), .B2(new_n895), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n965), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n991), .A2(new_n953), .A3(new_n994), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n995), .A2(new_n942), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n987), .A2(new_n989), .A3(new_n990), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n960), .A2(KEYINPUT108), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT107), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n964), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n961), .A2(new_n962), .A3(KEYINPUT107), .A4(new_n963), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT108), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n1002), .B(KEYINPUT41), .C1(new_n958), .C2(new_n959), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n998), .A2(new_n1000), .A3(new_n1001), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n997), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n989), .A2(new_n966), .A3(new_n985), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n953), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT43), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n996), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n995), .A2(new_n942), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n953), .B1(new_n991), .B2(new_n994), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT43), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n976), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n953), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1016), .A2(new_n1012), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT109), .B1(new_n1017), .B2(new_n1010), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n975), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1020), .A2(KEYINPUT43), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n1016), .A2(new_n1012), .A3(new_n1010), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT44), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1019), .A2(new_n1023), .ZN(G397));
  INV_X1    g599(.A(new_n498), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n491), .A2(new_n492), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1384), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n466), .A2(new_n472), .A3(G40), .A4(new_n473), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n1029), .A2(KEYINPUT45), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G1996), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1032), .B1(new_n922), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n1033), .B2(new_n922), .ZN(new_n1035));
  INV_X1    g610(.A(G2067), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n799), .B(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT111), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1037), .A2(new_n1038), .A3(new_n1031), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1038), .B1(new_n1037), .B2(new_n1031), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1035), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT112), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g618(.A(KEYINPUT112), .B(new_n1035), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n847), .A2(new_n854), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n799), .A2(new_n1036), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1032), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT46), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1049), .B1(KEYINPUT127), .B2(new_n1050), .ZN(new_n1051));
  XOR2_X1   g626(.A(KEYINPUT127), .B(KEYINPUT46), .Z(new_n1052));
  AOI21_X1  g627(.A(new_n1051), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1031), .B1(new_n1037), .B2(new_n922), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g630(.A(new_n1055), .B(KEYINPUT47), .Z(new_n1056));
  INV_X1    g631(.A(G1986), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n621), .A2(new_n1057), .ZN(new_n1058));
  XOR2_X1   g633(.A(new_n1058), .B(KEYINPUT110), .Z(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n1031), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n1060), .B(KEYINPUT48), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n847), .A2(new_n854), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1031), .B1(new_n1062), .B2(new_n1045), .ZN(new_n1063));
  AND4_X1   g638(.A1(new_n1043), .A2(new_n1061), .A3(new_n1044), .A4(new_n1063), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1048), .A2(new_n1056), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n582), .A2(G8), .A3(new_n584), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n582), .A2(KEYINPUT55), .A3(G8), .A4(new_n584), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G1384), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(new_n493), .B2(new_n498), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT45), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1030), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g650(.A(KEYINPUT45), .B(new_n1072), .C1(new_n493), .C2(new_n498), .ZN(new_n1076));
  AOI21_X1  g651(.A(G1971), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT50), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1078), .B(new_n1072), .C1(new_n493), .C2(new_n498), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n1080));
  XNOR2_X1  g655(.A(new_n1079), .B(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1073), .A2(KEYINPUT50), .ZN(new_n1082));
  AND4_X1   g657(.A1(G40), .A2(new_n466), .A3(new_n472), .A4(new_n473), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT115), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1030), .B1(new_n1073), .B2(KEYINPUT50), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1081), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1077), .B1(new_n1089), .B2(new_n815), .ZN(new_n1090));
  INV_X1    g665(.A(G8), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1071), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G1976), .ZN(new_n1093));
  OAI221_X1 g668(.A(G8), .B1(new_n589), .B2(new_n1093), .C1(new_n1073), .C2(new_n1030), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT52), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n594), .B2(G1976), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1095), .B1(new_n1097), .B2(new_n1094), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT49), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n832), .A2(G1981), .A3(new_n834), .ZN(new_n1100));
  INV_X1    g675(.A(G1981), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1101), .B1(new_n607), .B2(new_n613), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1099), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT114), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(G1981), .B1(new_n832), .B2(new_n834), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n607), .A2(new_n1101), .A3(new_n613), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1108), .A2(KEYINPUT114), .A3(new_n1099), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1106), .A2(KEYINPUT49), .A3(new_n1107), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1091), .B1(new_n1029), .B2(new_n1083), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1098), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1086), .A2(new_n815), .A3(new_n1079), .ZN(new_n1115));
  OAI21_X1  g690(.A(G8), .B1(new_n1115), .B2(new_n1077), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n1070), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT117), .B(G2084), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1086), .A2(new_n1079), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n740), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1122), .A2(new_n1091), .A3(G286), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1092), .A2(new_n1114), .A3(new_n1118), .A4(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT63), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT114), .B1(new_n1108), .B2(new_n1099), .ZN(new_n1127));
  AOI211_X1 g702(.A(new_n1104), .B(KEYINPUT49), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1113), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1098), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1116), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(KEYINPUT118), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1118), .A2(new_n1123), .A3(KEYINPUT63), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT118), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1129), .A2(new_n1131), .A3(new_n1130), .A4(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1133), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1126), .A2(new_n1137), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1092), .A2(new_n1114), .A3(new_n1118), .ZN(new_n1139));
  INV_X1    g714(.A(G2078), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1075), .A2(new_n1140), .A3(new_n1076), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT53), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1086), .A2(new_n1079), .ZN(new_n1143));
  AOI22_X1  g718(.A1(new_n1141), .A2(new_n1142), .B1(new_n1143), .B2(new_n754), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1142), .A2(G2078), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1075), .A2(new_n1076), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(G301), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1122), .A2(G168), .ZN(new_n1148));
  OAI21_X1  g723(.A(G286), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1148), .A2(G8), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT51), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT62), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1091), .B1(new_n1122), .B2(G168), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT51), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1151), .A2(new_n1152), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1154), .B1(new_n1153), .B2(new_n1149), .ZN(new_n1157));
  AOI211_X1 g732(.A(KEYINPUT51), .B(new_n1091), .C1(new_n1122), .C2(G168), .ZN(new_n1158));
  OAI21_X1  g733(.A(KEYINPUT62), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1139), .A2(new_n1147), .A3(new_n1156), .A4(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1129), .A2(new_n1093), .A3(new_n594), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(new_n1107), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1118), .ZN(new_n1163));
  AOI22_X1  g738(.A1(new_n1162), .A2(new_n1112), .B1(new_n1114), .B2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1138), .A2(new_n1160), .A3(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1144), .A2(G301), .A3(new_n1146), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n1075), .A2(KEYINPUT125), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1075), .A2(KEYINPUT125), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1168), .A2(new_n1076), .A3(new_n1169), .A4(new_n1145), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n1144), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1167), .B1(new_n1171), .B2(G171), .ZN(new_n1172));
  AOI211_X1 g747(.A(KEYINPUT126), .B(G301), .C1(new_n1170), .C2(new_n1144), .ZN(new_n1173));
  OAI211_X1 g748(.A(KEYINPUT54), .B(new_n1166), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT54), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1171), .A2(G171), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1175), .B1(new_n1176), .B2(new_n1147), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1139), .A2(new_n1174), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1079), .B(KEYINPUT116), .ZN(new_n1181));
  AOI211_X1 g756(.A(KEYINPUT115), .B(new_n1030), .C1(KEYINPUT50), .C2(new_n1073), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1087), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(G1956), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g761(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n640), .B(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g763(.A(KEYINPUT56), .B(G2072), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1075), .A2(new_n1076), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT120), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1075), .A2(KEYINPUT120), .A3(new_n1076), .A4(new_n1189), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  AND3_X1   g769(.A1(new_n1186), .A2(new_n1188), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1188), .B1(new_n1186), .B2(new_n1194), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1180), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT121), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1029), .A2(new_n1083), .A3(new_n1198), .ZN(new_n1199));
  OAI21_X1  g774(.A(KEYINPUT121), .B1(new_n1073), .B2(new_n1030), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n1036), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT60), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT123), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1203), .B1(new_n636), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(G1348), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1143), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1202), .A2(new_n1205), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g783(.A(G2067), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1209));
  AOI21_X1  g784(.A(G1348), .B1(new_n1086), .B2(new_n1079), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1203), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n957), .A2(KEYINPUT123), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1208), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1214));
  NAND4_X1  g789(.A1(new_n1214), .A2(KEYINPUT123), .A3(KEYINPUT60), .A4(new_n957), .ZN(new_n1215));
  XOR2_X1   g790(.A(KEYINPUT58), .B(G1341), .Z(new_n1216));
  NAND3_X1  g791(.A1(new_n1199), .A2(new_n1200), .A3(new_n1216), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1075), .A2(new_n1033), .A3(new_n1076), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1219), .A2(new_n558), .ZN(new_n1220));
  INV_X1    g795(.A(KEYINPUT59), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g797(.A1(new_n1219), .A2(KEYINPUT59), .A3(new_n558), .ZN(new_n1223));
  AND4_X1   g798(.A1(new_n1213), .A2(new_n1215), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1194), .B1(new_n1089), .B2(G1956), .ZN(new_n1225));
  INV_X1    g800(.A(new_n1188), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g802(.A1(new_n1186), .A2(new_n1188), .A3(new_n1194), .ZN(new_n1228));
  NAND3_X1  g803(.A1(new_n1227), .A2(KEYINPUT61), .A3(new_n1228), .ZN(new_n1229));
  NAND3_X1  g804(.A1(new_n1197), .A2(new_n1224), .A3(new_n1229), .ZN(new_n1230));
  NOR2_X1   g805(.A1(new_n1214), .A2(new_n957), .ZN(new_n1231));
  OAI211_X1 g806(.A(KEYINPUT122), .B(new_n1228), .C1(new_n1196), .C2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g807(.A(new_n1228), .B1(new_n1196), .B2(new_n1231), .ZN(new_n1233));
  INV_X1    g808(.A(KEYINPUT122), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g810(.A1(new_n1230), .A2(new_n1232), .A3(new_n1235), .ZN(new_n1236));
  AOI21_X1  g811(.A(new_n1179), .B1(new_n1236), .B2(KEYINPUT124), .ZN(new_n1237));
  INV_X1    g812(.A(KEYINPUT124), .ZN(new_n1238));
  NAND4_X1  g813(.A1(new_n1230), .A2(new_n1232), .A3(new_n1235), .A4(new_n1238), .ZN(new_n1239));
  AOI21_X1  g814(.A(new_n1165), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1240));
  NOR2_X1   g815(.A1(new_n621), .A2(new_n1057), .ZN(new_n1241));
  OAI21_X1  g816(.A(new_n1031), .B1(new_n1059), .B2(new_n1241), .ZN(new_n1242));
  NAND4_X1  g817(.A1(new_n1043), .A2(new_n1044), .A3(new_n1063), .A4(new_n1242), .ZN(new_n1243));
  XNOR2_X1  g818(.A(new_n1243), .B(KEYINPUT113), .ZN(new_n1244));
  OAI21_X1  g819(.A(new_n1065), .B1(new_n1240), .B2(new_n1244), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g820(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1247));
  OR3_X1    g821(.A1(G401), .A2(new_n457), .A3(G227), .ZN(new_n1248));
  AOI21_X1  g822(.A(new_n1248), .B1(new_n713), .B2(new_n714), .ZN(new_n1249));
  OAI21_X1  g823(.A(new_n1249), .B1(new_n943), .B2(new_n944), .ZN(new_n1250));
  NOR2_X1   g824(.A1(new_n1247), .A2(new_n1250), .ZN(G308));
  OAI221_X1 g825(.A(new_n1249), .B1(new_n943), .B2(new_n944), .C1(new_n1015), .C2(new_n1018), .ZN(G225));
endmodule


