//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(G110), .B(G140), .Z(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G227), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n189), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT10), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT65), .B1(new_n195), .B2(G146), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n195), .A2(G146), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n202));
  AND4_X1   g016(.A1(new_n196), .A2(new_n199), .A3(new_n200), .A4(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT1), .B1(new_n195), .B2(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT79), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT79), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n206), .B(KEYINPUT1), .C1(new_n195), .C2(G146), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(G128), .A3(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n196), .A2(new_n199), .A3(new_n200), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n203), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G104), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT3), .B1(new_n211), .B2(G107), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT3), .ZN(new_n213));
  INV_X1    g027(.A(G107), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(G104), .ZN(new_n215));
  INV_X1    g029(.A(G101), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n211), .A2(G107), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n212), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n211), .A2(G107), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n214), .A2(G104), .ZN(new_n220));
  OAI21_X1  g034(.A(G101), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n194), .B1(new_n210), .B2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n212), .A2(new_n215), .A3(new_n217), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G101), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(KEYINPUT4), .A3(new_n218), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n196), .A2(new_n199), .A3(new_n200), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT64), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n228), .B(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n198), .A2(G143), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n232), .B1(new_n233), .B2(new_n200), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n227), .A2(new_n229), .B1(new_n231), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT4), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n224), .A2(new_n236), .A3(G101), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n226), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n233), .A2(new_n200), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT68), .B(G128), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n241), .B1(G143), .B2(new_n198), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n239), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n196), .A2(new_n199), .A3(new_n200), .A4(new_n202), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n194), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  AND2_X1   g059(.A1(new_n218), .A2(new_n221), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n245), .A2(KEYINPUT80), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(KEYINPUT80), .B1(new_n245), .B2(new_n246), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n223), .B(new_n238), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G131), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT11), .ZN(new_n252));
  INV_X1    g066(.A(G137), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n251), .A2(new_n252), .A3(new_n253), .A4(G134), .ZN(new_n254));
  INV_X1    g068(.A(G134), .ZN(new_n255));
  OAI22_X1  g069(.A1(new_n255), .A2(G137), .B1(KEYINPUT66), .B2(KEYINPUT11), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n255), .A2(G137), .B1(KEYINPUT66), .B2(KEYINPUT11), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n250), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n250), .A3(new_n258), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n193), .B1(new_n249), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n222), .A2(new_n243), .A3(new_n244), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n207), .A2(G128), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n206), .B1(new_n233), .B2(KEYINPUT1), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n209), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n222), .B1(new_n268), .B2(new_n244), .ZN(new_n269));
  OAI211_X1 g083(.A(KEYINPUT12), .B(new_n262), .C1(new_n265), .C2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n264), .B1(new_n210), .B2(new_n222), .ZN(new_n272));
  AOI21_X1  g086(.A(KEYINPUT12), .B1(new_n272), .B2(new_n262), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n263), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n249), .A2(new_n262), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n243), .A2(new_n244), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n246), .A2(new_n277), .A3(KEYINPUT10), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT80), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n245), .A2(KEYINPUT80), .A3(new_n246), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n262), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n282), .A2(new_n283), .A3(new_n223), .A4(new_n238), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n193), .B1(new_n276), .B2(new_n284), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n187), .B(new_n188), .C1(new_n275), .C2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n276), .A2(new_n284), .A3(new_n193), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n262), .B1(new_n265), .B2(new_n269), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT12), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n270), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n291), .A2(new_n284), .ZN(new_n292));
  OAI211_X1 g106(.A(G469), .B(new_n287), .C1(new_n292), .C2(new_n193), .ZN(new_n293));
  NAND2_X1  g107(.A1(G469), .A2(G902), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n286), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(KEYINPUT9), .B(G234), .ZN(new_n296));
  OAI21_X1  g110(.A(G221), .B1(new_n296), .B2(G902), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n295), .A2(KEYINPUT81), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(KEYINPUT81), .B1(new_n295), .B2(new_n297), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G214), .B1(G237), .B2(G902), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT6), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n226), .A2(new_n237), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT69), .ZN(new_n305));
  INV_X1    g119(.A(G116), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(G119), .ZN(new_n307));
  INV_X1    g121(.A(G119), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n308), .A2(G116), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n305), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT2), .B(G113), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(G116), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n306), .A2(G119), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n313), .A3(KEYINPUT69), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n310), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT70), .ZN(new_n316));
  XOR2_X1   g130(.A(KEYINPUT2), .B(G113), .Z(new_n317));
  INV_X1    g131(.A(KEYINPUT71), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n317), .A2(new_n318), .A3(new_n312), .A4(new_n313), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n312), .A2(new_n313), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT71), .B1(new_n320), .B2(new_n311), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT70), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n310), .A2(new_n323), .A3(new_n311), .A4(new_n314), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n316), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  AND3_X1   g139(.A1(new_n312), .A2(new_n313), .A3(KEYINPUT69), .ZN(new_n326));
  AOI21_X1  g140(.A(KEYINPUT69), .B1(new_n312), .B2(new_n313), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT5), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G113), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT5), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n329), .B1(new_n307), .B2(new_n330), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n328), .A2(new_n331), .B1(new_n319), .B2(new_n321), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n304), .A2(new_n325), .B1(new_n246), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(G110), .B(G122), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n303), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n334), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT82), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n336), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n304), .A2(new_n325), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n332), .A2(new_n246), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n339), .A2(new_n337), .A3(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n335), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT83), .ZN(new_n343));
  OR3_X1    g157(.A1(new_n338), .A2(new_n341), .A3(KEYINPUT6), .ZN(new_n344));
  MUX2_X1   g158(.A(new_n277), .B(new_n235), .S(G125), .Z(new_n345));
  NAND2_X1  g159(.A1(new_n190), .A2(G224), .ZN(new_n346));
  XOR2_X1   g160(.A(new_n346), .B(KEYINPUT84), .Z(new_n347));
  XOR2_X1   g161(.A(new_n345), .B(new_n347), .Z(new_n348));
  INV_X1    g162(.A(KEYINPUT83), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n349), .B(new_n335), .C1(new_n338), .C2(new_n341), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n343), .A2(new_n344), .A3(new_n348), .A4(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n328), .A2(new_n331), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n322), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT85), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(new_n222), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT85), .B1(new_n332), .B2(new_n246), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n331), .B1(new_n330), .B2(new_n320), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n322), .A2(new_n246), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n355), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n334), .B(KEYINPUT8), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT86), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT86), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n359), .A2(new_n363), .A3(new_n360), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n346), .A2(KEYINPUT7), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n345), .B(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n367), .B1(new_n333), .B2(new_n334), .ZN(new_n368));
  AOI21_X1  g182(.A(G902), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n351), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(G210), .B1(G237), .B2(G902), .ZN(new_n371));
  XOR2_X1   g185(.A(new_n371), .B(KEYINPUT87), .Z(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n351), .A2(new_n369), .A3(new_n371), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n302), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(G116), .B(G122), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n214), .ZN(new_n377));
  INV_X1    g191(.A(G122), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT14), .B1(new_n378), .B2(G116), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n379), .B1(new_n306), .B2(G122), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT95), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n306), .A2(G122), .ZN(new_n383));
  OAI21_X1  g197(.A(KEYINPUT95), .B1(new_n383), .B2(KEYINPUT14), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n382), .B(G107), .C1(new_n380), .C2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n201), .A2(KEYINPUT68), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT68), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G128), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n388), .A3(G143), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT93), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n240), .A2(KEYINPUT93), .A3(G143), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n201), .A2(G143), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n255), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  AOI211_X1 g210(.A(G134), .B(new_n394), .C1(new_n391), .C2(new_n392), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n377), .B(new_n385), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G217), .ZN(new_n399));
  NOR3_X1   g213(.A1(new_n296), .A2(new_n399), .A3(G953), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n394), .A2(KEYINPUT13), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n394), .A2(KEYINPUT13), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n403), .B1(new_n391), .B2(new_n392), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n402), .B1(new_n404), .B2(KEYINPUT94), .ZN(new_n405));
  INV_X1    g219(.A(new_n403), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT93), .B1(new_n240), .B2(G143), .ZN(new_n407));
  AND4_X1   g221(.A1(KEYINPUT93), .A2(new_n386), .A3(new_n388), .A4(G143), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT94), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n255), .B1(new_n405), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n393), .A2(new_n255), .A3(new_n395), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n376), .B(new_n214), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n398), .B(new_n400), .C1(new_n412), .C2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT96), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n398), .B1(new_n412), .B2(new_n415), .ZN(new_n419));
  INV_X1    g233(.A(new_n400), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(KEYINPUT94), .B(new_n406), .C1(new_n407), .C2(new_n408), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n401), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n404), .A2(KEYINPUT94), .ZN(new_n424));
  OAI21_X1  g238(.A(G134), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n415), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n427), .A2(KEYINPUT96), .A3(new_n398), .A4(new_n400), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n418), .A2(new_n421), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G478), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(KEYINPUT15), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n429), .A2(new_n188), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n432), .B1(new_n429), .B2(new_n188), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n378), .A2(G113), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n329), .A2(G122), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(new_n437), .A3(G104), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(G104), .B1(new_n436), .B2(new_n437), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(G237), .A2(G953), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n442), .A2(G143), .A3(G214), .ZN(new_n443));
  AOI21_X1  g257(.A(G143), .B1(new_n442), .B2(G214), .ZN(new_n444));
  OAI21_X1  g258(.A(G131), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n442), .A2(G214), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n195), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n442), .A2(G143), .A3(G214), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n250), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT88), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(G125), .B(G140), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT16), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT16), .ZN(new_n455));
  INV_X1    g269(.A(G140), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n456), .A3(G125), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n454), .A2(G146), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n445), .A2(new_n449), .A3(KEYINPUT88), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n456), .A2(G125), .ZN(new_n460));
  INV_X1    g274(.A(G125), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G140), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT19), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n460), .B(new_n462), .C1(KEYINPUT89), .C2(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n464), .B(new_n198), .C1(new_n453), .C2(new_n465), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n452), .A2(new_n458), .A3(new_n459), .A4(new_n466), .ZN(new_n467));
  OAI211_X1 g281(.A(KEYINPUT18), .B(G131), .C1(new_n443), .C2(new_n444), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n460), .A2(new_n462), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G146), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n453), .A2(new_n198), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(KEYINPUT18), .A2(G131), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n447), .A2(new_n448), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n468), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n441), .B1(new_n467), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT17), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n445), .A2(new_n449), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n457), .B1(new_n469), .B2(new_n455), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n198), .ZN(new_n480));
  OAI211_X1 g294(.A(KEYINPUT17), .B(G131), .C1(new_n443), .C2(new_n444), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n478), .A2(new_n480), .A3(new_n458), .A4(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT90), .ZN(new_n483));
  INV_X1    g297(.A(new_n440), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n483), .B1(new_n484), .B2(new_n438), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n439), .A2(new_n440), .A3(KEYINPUT90), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n482), .A2(new_n475), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n476), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(G475), .A2(G902), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(KEYINPUT91), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n475), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT88), .B1(new_n445), .B2(new_n449), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n466), .A2(new_n458), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n494), .B1(new_n497), .B2(new_n459), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n488), .B1(new_n498), .B2(new_n441), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT91), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n500), .A3(new_n491), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n493), .A2(KEYINPUT20), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT20), .ZN(new_n503));
  OAI211_X1 g317(.A(KEYINPUT91), .B(new_n503), .C1(new_n490), .C2(new_n492), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n480), .A2(new_n481), .A3(new_n458), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n445), .A2(new_n449), .A3(new_n477), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n475), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n441), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(G902), .B1(new_n509), .B2(new_n488), .ZN(new_n510));
  OR2_X1    g324(.A1(new_n510), .A2(KEYINPUT92), .ZN(new_n511));
  INV_X1    g325(.A(G475), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n512), .B1(new_n510), .B2(KEYINPUT92), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n502), .A2(new_n504), .A3(new_n514), .ZN(new_n515));
  AOI211_X1 g329(.A(new_n188), .B(new_n190), .C1(G234), .C2(G237), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT21), .B(G898), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n190), .A2(G952), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(G234), .B2(G237), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n435), .A2(new_n515), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n300), .A2(new_n375), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT67), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n255), .A2(G137), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n253), .A2(G134), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n525), .B(G131), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(G134), .B(G137), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT67), .B1(new_n529), .B2(new_n250), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n261), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n531), .A2(KEYINPUT72), .B1(new_n243), .B2(new_n244), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT72), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n261), .A2(new_n533), .A3(new_n528), .A4(new_n530), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n532), .A2(new_n534), .B1(new_n262), .B2(new_n235), .ZN(new_n535));
  INV_X1    g349(.A(new_n325), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n442), .A2(G210), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(KEYINPUT27), .ZN(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT26), .B(G101), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n539), .B(new_n540), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n257), .A2(new_n250), .A3(new_n258), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n235), .B1(new_n542), .B2(new_n259), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT30), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n277), .A2(new_n261), .A3(new_n528), .A4(new_n530), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n530), .A2(new_n528), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT72), .B1(new_n542), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n548), .A2(new_n277), .A3(new_n534), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n543), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n546), .B1(new_n550), .B2(KEYINPUT30), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n537), .B(new_n541), .C1(new_n551), .C2(new_n536), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT31), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n543), .A2(new_n545), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n325), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT28), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n556), .B1(new_n535), .B2(new_n536), .ZN(new_n557));
  AND4_X1   g371(.A1(new_n556), .A2(new_n549), .A3(new_n543), .A4(new_n536), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n555), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n541), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n544), .B1(new_n549), .B2(new_n543), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n325), .B1(new_n562), .B2(new_n546), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT31), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n563), .A2(new_n564), .A3(new_n537), .A4(new_n541), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n553), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(G472), .A2(G902), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  XOR2_X1   g382(.A(KEYINPUT73), .B(KEYINPUT32), .Z(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n566), .A2(KEYINPUT32), .A3(new_n567), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n559), .A2(new_n541), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n563), .A2(new_n537), .A3(new_n560), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT29), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI22_X1  g389(.A1(new_n557), .A2(new_n558), .B1(new_n536), .B2(new_n535), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n541), .A2(KEYINPUT29), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n188), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(G472), .B1(new_n575), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n571), .A2(new_n572), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(KEYINPUT76), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT22), .B(G137), .ZN(new_n583));
  XOR2_X1   g397(.A(new_n582), .B(new_n583), .Z(new_n584));
  NAND2_X1  g398(.A1(new_n240), .A2(G119), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n308), .A2(G128), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT24), .B(G110), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n479), .A2(new_n198), .ZN(new_n590));
  AOI21_X1  g404(.A(G146), .B1(new_n454), .B2(new_n457), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n240), .A2(KEYINPUT23), .A3(G119), .ZN(new_n593));
  AND2_X1   g407(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n594));
  NOR2_X1   g408(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n595));
  OAI22_X1  g409(.A1(new_n594), .A2(new_n595), .B1(new_n308), .B2(G128), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n593), .A2(new_n596), .A3(KEYINPUT75), .A4(new_n586), .ZN(new_n597));
  INV_X1    g411(.A(G110), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n593), .A2(new_n586), .A3(new_n596), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT75), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n592), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n593), .A2(new_n596), .A3(new_n598), .A4(new_n586), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n585), .A2(new_n586), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n603), .B1(new_n604), .B2(new_n588), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n605), .A2(new_n458), .A3(new_n471), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n584), .B1(new_n602), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n599), .A2(new_n600), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n608), .A2(G110), .A3(new_n597), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n480), .A2(new_n458), .B1(new_n604), .B2(new_n588), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n605), .A2(new_n458), .A3(new_n471), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n582), .B(new_n583), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n607), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n399), .B1(G234), .B2(new_n188), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n615), .A2(G902), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n616), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n607), .A2(new_n188), .A3(new_n614), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT77), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT25), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n618), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n619), .A2(KEYINPUT77), .A3(KEYINPUT25), .ZN(new_n623));
  AOI211_X1 g437(.A(KEYINPUT78), .B(new_n617), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT78), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n620), .A2(new_n621), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n626), .A2(new_n623), .A3(new_n616), .ZN(new_n627));
  INV_X1    g441(.A(new_n617), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n580), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n524), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(new_n216), .ZN(G3));
  INV_X1    g447(.A(new_n568), .ZN(new_n634));
  INV_X1    g448(.A(G472), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n566), .B2(new_n188), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n300), .A2(new_n630), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT97), .ZN(new_n639));
  INV_X1    g453(.A(new_n371), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n370), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT98), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n641), .A2(new_n642), .A3(new_n374), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT33), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n429), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n421), .A2(KEYINPUT33), .A3(new_n416), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n430), .A2(G902), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n429), .A2(new_n188), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n430), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n500), .B1(new_n499), .B2(new_n491), .ZN(new_n652));
  AOI22_X1  g466(.A1(new_n511), .A2(new_n513), .B1(new_n652), .B2(new_n503), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n502), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n351), .A2(KEYINPUT98), .A3(new_n369), .A4(new_n371), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n657), .A2(new_n301), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n643), .A2(new_n656), .A3(new_n658), .A4(new_n522), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n639), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT34), .B(G104), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G6));
  OAI211_X1 g477(.A(new_n515), .B(new_n522), .C1(new_n434), .C2(new_n433), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT99), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n435), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n667), .A2(KEYINPUT99), .A3(new_n515), .A4(new_n522), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n666), .A2(new_n668), .A3(new_n643), .A4(new_n658), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n639), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT35), .B(G107), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  NAND2_X1  g487(.A1(new_n611), .A2(new_n612), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n584), .A2(KEYINPUT36), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n676), .A2(new_n188), .A3(new_n618), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(new_n622), .B2(new_n623), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n634), .A2(new_n636), .A3(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n679), .A2(new_n300), .A3(new_n375), .A4(new_n523), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT37), .B(G110), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G12));
  INV_X1    g496(.A(new_n678), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n300), .A2(new_n580), .A3(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(G900), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n520), .B1(new_n516), .B2(new_n685), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n435), .A2(new_n654), .A3(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n643), .A2(new_n658), .A3(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n201), .ZN(G30));
  NAND2_X1  g504(.A1(new_n537), .A2(new_n560), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n535), .A2(new_n536), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n188), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n560), .B1(new_n563), .B2(new_n537), .ZN(new_n694));
  OAI21_X1  g508(.A(G472), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(KEYINPUT100), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT100), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n697), .B(G472), .C1(new_n693), .C2(new_n694), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n571), .A2(new_n572), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT101), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  XOR2_X1   g516(.A(new_n686), .B(KEYINPUT39), .Z(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n298), .A2(new_n299), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT40), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n435), .A2(new_n515), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n301), .A3(new_n678), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n373), .A2(new_n374), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n709), .A2(KEYINPUT38), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(KEYINPUT38), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n708), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n702), .A2(new_n706), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G143), .ZN(G45));
  AND3_X1   g528(.A1(new_n300), .A2(new_n580), .A3(new_n683), .ZN(new_n715));
  AOI221_X4 g529(.A(new_n686), .B1(new_n653), .B2(new_n502), .C1(new_n648), .C2(new_n650), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n643), .A2(new_n716), .A3(new_n658), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G146), .ZN(G48));
  OAI21_X1  g534(.A(new_n188), .B1(new_n275), .B2(new_n285), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(G469), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n286), .ZN(new_n723));
  INV_X1    g537(.A(new_n297), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n580), .A2(new_n630), .A3(new_n725), .ZN(new_n726));
  OR2_X1    g540(.A1(new_n659), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT41), .B(G113), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G15));
  OR2_X1    g543(.A1(new_n669), .A2(new_n726), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G116), .ZN(G18));
  NAND3_X1  g545(.A1(new_n580), .A2(new_n523), .A3(new_n683), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n643), .A2(new_n658), .A3(new_n725), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n308), .ZN(G21));
  NAND3_X1  g549(.A1(new_n643), .A2(new_n658), .A3(new_n707), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n566), .A2(new_n188), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n576), .A2(new_n560), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n553), .A2(new_n738), .A3(new_n565), .ZN(new_n739));
  AOI22_X1  g553(.A1(new_n737), .A2(G472), .B1(new_n567), .B2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n627), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n617), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n740), .A2(new_n742), .A3(new_n522), .A4(new_n725), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n736), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n378), .ZN(G24));
  NAND3_X1  g559(.A1(new_n716), .A2(new_n683), .A3(new_n740), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n733), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n461), .ZN(G27));
  NAND2_X1  g562(.A1(new_n295), .A2(new_n297), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n750), .A2(new_n373), .A3(new_n374), .A4(new_n301), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT32), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n568), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n572), .A3(new_n579), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n752), .A2(new_n742), .A3(new_n716), .A4(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n631), .A2(new_n751), .ZN(new_n757));
  INV_X1    g571(.A(new_n686), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n651), .A2(new_n654), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(KEYINPUT42), .ZN(new_n760));
  AOI22_X1  g574(.A1(new_n756), .A2(KEYINPUT42), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G131), .ZN(G33));
  INV_X1    g576(.A(new_n631), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n687), .A3(new_n752), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  INV_X1    g579(.A(KEYINPUT104), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT43), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n648), .A2(new_n650), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n654), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT103), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n767), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI211_X1 g585(.A(KEYINPUT103), .B(KEYINPUT43), .C1(new_n768), .C2(new_n654), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n766), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n771), .A2(new_n766), .A3(new_n772), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n637), .A2(new_n678), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n774), .A2(KEYINPUT44), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n775), .A2(new_n776), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n778), .B1(new_n779), .B2(new_n773), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n287), .B1(new_n292), .B2(new_n193), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n187), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n783), .B1(new_n782), .B2(new_n781), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n294), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT46), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n784), .A2(KEYINPUT46), .A3(new_n294), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(new_n286), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n297), .ZN(new_n790));
  OAI21_X1  g604(.A(KEYINPUT102), .B1(new_n790), .B2(new_n704), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT102), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n789), .A2(new_n792), .A3(new_n297), .A4(new_n703), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n373), .A2(new_n374), .A3(new_n301), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n777), .A2(new_n780), .A3(new_n794), .A4(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G137), .ZN(G39));
  INV_X1    g612(.A(KEYINPUT47), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n790), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n789), .A2(KEYINPUT47), .A3(new_n297), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR4_X1   g616(.A1(new_n580), .A2(new_n630), .A3(new_n795), .A4(new_n759), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G140), .ZN(G42));
  INV_X1    g619(.A(KEYINPUT50), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n710), .A2(new_n711), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(new_n302), .A3(new_n725), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n740), .A2(new_n742), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n771), .A2(new_n809), .A3(new_n520), .A4(new_n772), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n806), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n771), .ZN(new_n812));
  INV_X1    g626(.A(new_n772), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n812), .A2(new_n521), .A3(new_n813), .ZN(new_n814));
  AND4_X1   g628(.A1(new_n302), .A2(new_n710), .A3(new_n711), .A4(new_n725), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n814), .A2(new_n815), .A3(KEYINPUT50), .A4(new_n809), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n722), .A2(new_n724), .A3(new_n286), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n800), .A2(new_n801), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n810), .A2(new_n795), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n818), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n739), .A2(new_n567), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n823), .A2(new_n636), .A3(new_n678), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n795), .A2(new_n724), .A3(new_n723), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n814), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n825), .A2(new_n630), .A3(new_n520), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(new_n515), .A3(new_n768), .A4(new_n701), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n826), .A2(KEYINPUT112), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT112), .B1(new_n826), .B2(new_n828), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n817), .B(new_n822), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n827), .A2(new_n656), .A3(new_n701), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n810), .A2(new_n733), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n519), .B(KEYINPUT113), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT114), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n814), .A2(new_n825), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n755), .A2(new_n742), .ZN(new_n839));
  OR3_X1    g653(.A1(new_n838), .A2(KEYINPUT48), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT48), .B1(new_n838), .B2(new_n839), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n831), .A2(new_n837), .A3(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n819), .B(KEYINPUT110), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n821), .B1(new_n802), .B2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n817), .A2(new_n826), .A3(new_n828), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n818), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT111), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n846), .A2(KEYINPUT111), .A3(new_n818), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n843), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  XNOR2_X1  g665(.A(KEYINPUT109), .B(KEYINPUT53), .ZN(new_n852));
  INV_X1    g666(.A(new_n688), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n643), .A2(new_n658), .A3(new_n725), .ZN(new_n854));
  NOR4_X1   g668(.A1(new_n759), .A2(new_n823), .A3(new_n636), .A4(new_n678), .ZN(new_n855));
  AOI22_X1  g669(.A1(new_n715), .A2(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n643), .A2(new_n658), .A3(new_n707), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n678), .A2(new_n297), .A3(new_n295), .A4(new_n758), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n568), .A2(new_n570), .B1(new_n696), .B2(new_n698), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n858), .B1(new_n859), .B2(new_n572), .ZN(new_n860));
  AOI22_X1  g674(.A1(new_n715), .A2(new_n718), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT52), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n856), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT108), .ZN(new_n864));
  INV_X1    g678(.A(new_n858), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n700), .A2(new_n865), .ZN(new_n866));
  OAI22_X1  g680(.A1(new_n684), .A2(new_n717), .B1(new_n866), .B2(new_n736), .ZN(new_n867));
  OAI22_X1  g681(.A1(new_n684), .A2(new_n688), .B1(new_n733), .B2(new_n746), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT52), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n863), .A2(new_n864), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n864), .B1(new_n863), .B2(new_n869), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n855), .A2(new_n752), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n764), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n435), .A2(new_n515), .A3(new_n758), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT105), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n435), .A2(new_n515), .A3(KEYINPUT105), .A4(new_n758), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n796), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(new_n684), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT106), .B1(new_n874), .B2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n880), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT106), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n882), .A2(new_n883), .A3(new_n764), .A4(new_n873), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n726), .B1(new_n669), .B2(new_n659), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n680), .B1(new_n524), .B2(new_n631), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI22_X1  g702(.A1(new_n732), .A2(new_n733), .B1(new_n736), .B2(new_n743), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n655), .B1(new_n435), .B2(new_n654), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n890), .A2(new_n630), .A3(new_n522), .A4(new_n637), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n300), .A2(new_n375), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n888), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n885), .A2(new_n761), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n852), .B1(new_n872), .B2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n862), .B1(new_n856), .B2(new_n861), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n867), .A2(new_n868), .A3(KEYINPUT52), .ZN(new_n900));
  OAI21_X1  g714(.A(KEYINPUT107), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT107), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n863), .A2(new_n902), .A3(new_n869), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n888), .A2(new_n894), .A3(new_n761), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n884), .B2(new_n881), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n904), .A2(new_n906), .A3(KEYINPUT53), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n897), .A2(new_n898), .A3(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n872), .A2(new_n896), .ZN(new_n909));
  INV_X1    g723(.A(new_n852), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n904), .A2(new_n906), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT53), .ZN(new_n912));
  AOI22_X1  g726(.A1(new_n909), .A2(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n851), .B(new_n908), .C1(new_n898), .C2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(KEYINPUT115), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n913), .A2(new_n898), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT115), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n916), .A2(new_n917), .A3(new_n908), .A4(new_n851), .ZN(new_n918));
  OR2_X1    g732(.A1(G952), .A2(G953), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n915), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NOR4_X1   g734(.A1(new_n741), .A2(new_n617), .A3(new_n724), .A4(new_n302), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n723), .A2(KEYINPUT49), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n723), .A2(KEYINPUT49), .ZN(new_n923));
  AND4_X1   g737(.A1(new_n769), .A2(new_n921), .A3(new_n922), .A4(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n807), .A2(new_n701), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n920), .A2(new_n925), .ZN(G75));
  NAND3_X1  g740(.A1(new_n343), .A2(new_n344), .A3(new_n350), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(new_n348), .ZN(new_n928));
  XNOR2_X1  g742(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n928), .B(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n930), .A2(KEYINPUT56), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n897), .A2(new_n907), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(G902), .ZN(new_n933));
  INV_X1    g747(.A(new_n372), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n190), .A2(G952), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n933), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT117), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n939), .A2(new_n940), .A3(G210), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT56), .ZN(new_n942));
  INV_X1    g756(.A(G210), .ZN(new_n943));
  OAI21_X1  g757(.A(KEYINPUT117), .B1(new_n933), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n941), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n938), .B1(new_n945), .B2(new_n930), .ZN(G51));
  XOR2_X1   g760(.A(new_n294), .B(KEYINPUT57), .Z(new_n947));
  AND3_X1   g761(.A1(new_n904), .A2(KEYINPUT53), .A3(new_n906), .ZN(new_n948));
  OAI21_X1  g762(.A(KEYINPUT108), .B1(new_n899), .B2(new_n900), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n863), .A2(new_n864), .A3(new_n869), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n910), .B1(new_n951), .B2(new_n906), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n948), .A2(new_n952), .A3(KEYINPUT54), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n898), .B1(new_n897), .B2(new_n907), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n947), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(KEYINPUT118), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n275), .A2(new_n285), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT118), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n958), .B(new_n947), .C1(new_n953), .C2(new_n954), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n956), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n933), .A2(new_n784), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n936), .B1(new_n960), .B2(new_n961), .ZN(G54));
  NAND2_X1  g776(.A1(KEYINPUT58), .A2(G475), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT119), .Z(new_n964));
  AND3_X1   g778(.A1(new_n939), .A2(new_n499), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n499), .B1(new_n939), .B2(new_n964), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n965), .A2(new_n966), .A3(new_n936), .ZN(G60));
  NOR2_X1   g781(.A1(new_n953), .A2(new_n954), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n645), .A2(new_n646), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(G478), .A2(G902), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT59), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n937), .B1(new_n968), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n908), .B1(new_n913), .B2(new_n898), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n970), .B1(new_n975), .B2(new_n972), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n974), .A2(new_n976), .ZN(G63));
  NAND2_X1  g791(.A1(G217), .A2(G902), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT60), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n932), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n936), .B1(new_n981), .B2(new_n615), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n979), .B1(new_n897), .B2(new_n907), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT120), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n983), .A2(new_n984), .A3(new_n676), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n984), .B1(new_n983), .B2(new_n676), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n982), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT61), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n982), .B(KEYINPUT61), .C1(new_n985), .C2(new_n986), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(G66));
  INV_X1    g805(.A(G224), .ZN(new_n992));
  OAI21_X1  g806(.A(G953), .B1(new_n517), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n993), .B1(new_n895), .B2(G953), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n927), .B1(G898), .B2(new_n190), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n994), .B(new_n995), .ZN(G69));
  AND2_X1   g810(.A1(new_n797), .A2(new_n804), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n761), .A2(new_n764), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT123), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n761), .A2(KEYINPUT123), .A3(new_n764), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n856), .A2(new_n719), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n839), .A2(new_n736), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1003), .B1(new_n794), .B2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n997), .A2(KEYINPUT124), .A3(new_n1002), .A4(new_n1005), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n1002), .A2(new_n797), .A3(new_n804), .A4(new_n1005), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT124), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1006), .A2(new_n1009), .A3(new_n190), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n464), .B1(new_n453), .B2(new_n465), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT121), .Z(new_n1012));
  XNOR2_X1  g826(.A(new_n551), .B(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1013), .B1(G900), .B2(G953), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n713), .A2(new_n719), .A3(new_n856), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT62), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1016), .B(new_n1017), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n763), .A2(new_n705), .A3(new_n796), .A4(new_n890), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1019), .B(KEYINPUT122), .ZN(new_n1020));
  AND3_X1   g834(.A1(new_n1018), .A2(new_n997), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1013), .B1(new_n1021), .B2(G953), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1015), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1023), .B(new_n1024), .ZN(G72));
  NAND2_X1  g839(.A1(G472), .A2(G902), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(KEYINPUT63), .Z(new_n1027));
  NAND2_X1  g841(.A1(new_n574), .A2(new_n1027), .ZN(new_n1028));
  NOR3_X1   g842(.A1(new_n913), .A2(new_n694), .A3(new_n1028), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n1018), .A2(new_n997), .A3(new_n895), .A4(new_n1020), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1030), .A2(new_n1027), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1031), .A2(new_n694), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1032), .A2(KEYINPUT125), .ZN(new_n1033));
  INV_X1    g847(.A(KEYINPUT125), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1031), .A2(new_n1034), .A3(new_n694), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1029), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n1006), .A2(new_n1009), .A3(new_n895), .ZN(new_n1037));
  AND2_X1   g851(.A1(new_n1037), .A2(new_n1027), .ZN(new_n1038));
  OAI211_X1 g852(.A(KEYINPUT126), .B(new_n937), .C1(new_n1038), .C2(new_n574), .ZN(new_n1039));
  INV_X1    g853(.A(KEYINPUT126), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n574), .B1(new_n1037), .B2(new_n1027), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n1040), .B1(new_n1041), .B2(new_n936), .ZN(new_n1042));
  AND3_X1   g856(.A1(new_n1036), .A2(new_n1039), .A3(new_n1042), .ZN(G57));
endmodule


