

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593;

  XNOR2_X1 U321 ( .A(n423), .B(n422), .ZN(n551) );
  AND2_X1 U322 ( .A1(n425), .A2(n424), .ZN(n289) );
  XNOR2_X1 U323 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U324 ( .A(n339), .B(n338), .ZN(n342) );
  XNOR2_X1 U325 ( .A(n376), .B(KEYINPUT47), .ZN(n377) );
  XNOR2_X1 U326 ( .A(n378), .B(n377), .ZN(n386) );
  INV_X1 U327 ( .A(n551), .ZN(n424) );
  XNOR2_X1 U328 ( .A(n372), .B(n371), .ZN(n588) );
  INV_X1 U329 ( .A(n588), .ZN(n562) );
  XOR2_X1 U330 ( .A(n311), .B(n310), .Z(n555) );
  XOR2_X1 U331 ( .A(KEYINPUT28), .B(n476), .Z(n532) );
  XNOR2_X1 U332 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U333 ( .A(n466), .B(n465), .ZN(G1351GAT) );
  XOR2_X1 U334 ( .A(KEYINPUT67), .B(KEYINPUT65), .Z(n291) );
  XNOR2_X1 U335 ( .A(G197GAT), .B(G8GAT), .ZN(n290) );
  XNOR2_X1 U336 ( .A(n291), .B(n290), .ZN(n311) );
  INV_X1 U337 ( .A(G141GAT), .ZN(n292) );
  NAND2_X1 U338 ( .A1(G22GAT), .A2(n292), .ZN(n295) );
  INV_X1 U339 ( .A(G22GAT), .ZN(n293) );
  NAND2_X1 U340 ( .A1(n293), .A2(G141GAT), .ZN(n294) );
  NAND2_X1 U341 ( .A1(n295), .A2(n294), .ZN(n297) );
  XNOR2_X1 U342 ( .A(G36GAT), .B(G50GAT), .ZN(n296) );
  XNOR2_X1 U343 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U344 ( .A(n298), .B(G113GAT), .Z(n300) );
  XOR2_X1 U345 ( .A(G15GAT), .B(G1GAT), .Z(n359) );
  XNOR2_X1 U346 ( .A(G169GAT), .B(n359), .ZN(n299) );
  XNOR2_X1 U347 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U348 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n302) );
  NAND2_X1 U349 ( .A1(G229GAT), .A2(G233GAT), .ZN(n301) );
  XOR2_X1 U350 ( .A(n302), .B(n301), .Z(n303) );
  XNOR2_X1 U351 ( .A(n304), .B(n303), .ZN(n309) );
  XOR2_X1 U352 ( .A(KEYINPUT68), .B(KEYINPUT7), .Z(n306) );
  XNOR2_X1 U353 ( .A(G43GAT), .B(G29GAT), .ZN(n305) );
  XNOR2_X1 U354 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U355 ( .A(KEYINPUT8), .B(n307), .Z(n324) );
  XNOR2_X1 U356 ( .A(n324), .B(KEYINPUT29), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n310) );
  INV_X1 U358 ( .A(n555), .ZN(n579) );
  XOR2_X1 U359 ( .A(G85GAT), .B(KEYINPUT73), .Z(n313) );
  XNOR2_X1 U360 ( .A(G99GAT), .B(G92GAT), .ZN(n312) );
  XNOR2_X1 U361 ( .A(n313), .B(n312), .ZN(n340) );
  XOR2_X1 U362 ( .A(n340), .B(KEYINPUT10), .Z(n315) );
  XOR2_X1 U363 ( .A(G36GAT), .B(G190GAT), .Z(n396) );
  XNOR2_X1 U364 ( .A(G218GAT), .B(n396), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n315), .B(n314), .ZN(n320) );
  XNOR2_X1 U366 ( .A(G50GAT), .B(KEYINPUT76), .ZN(n316) );
  XOR2_X1 U367 ( .A(n316), .B(G162GAT), .Z(n426) );
  XNOR2_X1 U368 ( .A(G106GAT), .B(n426), .ZN(n318) );
  NAND2_X1 U369 ( .A1(G232GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n326) );
  XOR2_X1 U372 ( .A(KEYINPUT9), .B(KEYINPUT77), .Z(n322) );
  XNOR2_X1 U373 ( .A(G134GAT), .B(KEYINPUT11), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U376 ( .A(n326), .B(n325), .ZN(n482) );
  INV_X1 U377 ( .A(n482), .ZN(n565) );
  XOR2_X1 U378 ( .A(G78GAT), .B(G148GAT), .Z(n328) );
  XNOR2_X1 U379 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n432) );
  XOR2_X1 U381 ( .A(G64GAT), .B(KEYINPUT75), .Z(n330) );
  XNOR2_X1 U382 ( .A(G176GAT), .B(G204GAT), .ZN(n329) );
  XNOR2_X1 U383 ( .A(n330), .B(n329), .ZN(n397) );
  XNOR2_X1 U384 ( .A(n432), .B(n397), .ZN(n352) );
  XNOR2_X1 U385 ( .A(G57GAT), .B(KEYINPUT69), .ZN(n331) );
  XNOR2_X1 U386 ( .A(n331), .B(KEYINPUT13), .ZN(n354) );
  INV_X1 U387 ( .A(n354), .ZN(n333) );
  XOR2_X1 U388 ( .A(G120GAT), .B(G71GAT), .Z(n442) );
  INV_X1 U389 ( .A(n442), .ZN(n332) );
  NAND2_X1 U390 ( .A1(n333), .A2(n332), .ZN(n335) );
  NAND2_X1 U391 ( .A1(n354), .A2(n442), .ZN(n334) );
  NAND2_X1 U392 ( .A1(n335), .A2(n334), .ZN(n339) );
  AND2_X1 U393 ( .A1(G230GAT), .A2(G233GAT), .ZN(n337) );
  INV_X1 U394 ( .A(KEYINPUT71), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n340), .B(KEYINPUT33), .ZN(n341) );
  XNOR2_X1 U396 ( .A(n342), .B(n341), .ZN(n345) );
  XOR2_X1 U397 ( .A(KEYINPUT31), .B(KEYINPUT74), .Z(n344) );
  XNOR2_X1 U398 ( .A(KEYINPUT32), .B(KEYINPUT70), .ZN(n343) );
  XOR2_X1 U399 ( .A(n344), .B(n343), .Z(n346) );
  NAND2_X1 U400 ( .A1(n345), .A2(n346), .ZN(n350) );
  INV_X1 U401 ( .A(n345), .ZN(n348) );
  INV_X1 U402 ( .A(n346), .ZN(n347) );
  NAND2_X1 U403 ( .A1(n348), .A2(n347), .ZN(n349) );
  NAND2_X1 U404 ( .A1(n350), .A2(n349), .ZN(n351) );
  XOR2_X1 U405 ( .A(n352), .B(n351), .Z(n379) );
  XNOR2_X1 U406 ( .A(n379), .B(KEYINPUT41), .ZN(n513) );
  NAND2_X1 U407 ( .A1(n513), .A2(n555), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n353), .B(KEYINPUT46), .ZN(n373) );
  XOR2_X1 U409 ( .A(G22GAT), .B(G155GAT), .Z(n435) );
  XOR2_X1 U410 ( .A(G8GAT), .B(G183GAT), .Z(n394) );
  XNOR2_X1 U411 ( .A(n435), .B(n394), .ZN(n355) );
  XNOR2_X1 U412 ( .A(n355), .B(n333), .ZN(n363) );
  XNOR2_X1 U413 ( .A(G78GAT), .B(G211GAT), .ZN(n356) );
  XNOR2_X1 U414 ( .A(n356), .B(G71GAT), .ZN(n358) );
  XOR2_X1 U415 ( .A(KEYINPUT14), .B(G64GAT), .Z(n357) );
  XNOR2_X1 U416 ( .A(n358), .B(n357), .ZN(n361) );
  XOR2_X1 U417 ( .A(n359), .B(G127GAT), .Z(n360) );
  XNOR2_X1 U418 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U419 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U420 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n365) );
  NAND2_X1 U421 ( .A1(G231GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U422 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U423 ( .A(n367), .B(n366), .Z(n372) );
  XOR2_X1 U424 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n369) );
  XNOR2_X1 U425 ( .A(KEYINPUT78), .B(KEYINPUT79), .ZN(n368) );
  XNOR2_X1 U426 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U427 ( .A(n370), .B(KEYINPUT80), .ZN(n371) );
  NAND2_X1 U428 ( .A1(n373), .A2(n588), .ZN(n374) );
  XOR2_X1 U429 ( .A(n374), .B(KEYINPUT109), .Z(n375) );
  NOR2_X1 U430 ( .A1(n565), .A2(n375), .ZN(n378) );
  INV_X1 U431 ( .A(KEYINPUT110), .ZN(n376) );
  INV_X1 U432 ( .A(n379), .ZN(n469) );
  XNOR2_X1 U433 ( .A(n482), .B(KEYINPUT36), .ZN(n591) );
  NOR2_X1 U434 ( .A1(n588), .A2(n591), .ZN(n380) );
  XOR2_X1 U435 ( .A(KEYINPUT45), .B(n380), .Z(n381) );
  NOR2_X1 U436 ( .A1(n469), .A2(n381), .ZN(n382) );
  XNOR2_X1 U437 ( .A(n382), .B(KEYINPUT111), .ZN(n383) );
  NOR2_X1 U438 ( .A1(n383), .A2(n555), .ZN(n384) );
  XNOR2_X1 U439 ( .A(n384), .B(KEYINPUT112), .ZN(n385) );
  NOR2_X1 U440 ( .A1(n386), .A2(n385), .ZN(n387) );
  XOR2_X1 U441 ( .A(KEYINPUT48), .B(n387), .Z(n552) );
  XOR2_X1 U442 ( .A(G211GAT), .B(KEYINPUT21), .Z(n389) );
  XNOR2_X1 U443 ( .A(G197GAT), .B(G218GAT), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n389), .B(n388), .ZN(n431) );
  XOR2_X1 U445 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n391) );
  XNOR2_X1 U446 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n390) );
  XNOR2_X1 U447 ( .A(n391), .B(n390), .ZN(n443) );
  XOR2_X1 U448 ( .A(G92GAT), .B(n443), .Z(n393) );
  NAND2_X1 U449 ( .A1(G226GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U450 ( .A(n393), .B(n392), .ZN(n395) );
  XOR2_X1 U451 ( .A(n395), .B(n394), .Z(n399) );
  XNOR2_X1 U452 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U453 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U454 ( .A(n431), .B(n400), .ZN(n529) );
  NAND2_X1 U455 ( .A1(n552), .A2(n529), .ZN(n401) );
  XNOR2_X1 U456 ( .A(n401), .B(KEYINPUT54), .ZN(n402) );
  XNOR2_X1 U457 ( .A(n402), .B(KEYINPUT119), .ZN(n425) );
  XOR2_X1 U458 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n404) );
  XNOR2_X1 U459 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n403) );
  XNOR2_X1 U460 ( .A(n404), .B(n403), .ZN(n423) );
  XOR2_X1 U461 ( .A(G127GAT), .B(KEYINPUT0), .Z(n406) );
  XNOR2_X1 U462 ( .A(G113GAT), .B(G134GAT), .ZN(n405) );
  XNOR2_X1 U463 ( .A(n406), .B(n405), .ZN(n446) );
  XOR2_X1 U464 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n408) );
  XNOR2_X1 U465 ( .A(G141GAT), .B(KEYINPUT87), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n427) );
  XNOR2_X1 U467 ( .A(n446), .B(n427), .ZN(n421) );
  XOR2_X1 U468 ( .A(G85GAT), .B(G162GAT), .Z(n410) );
  XNOR2_X1 U469 ( .A(G29GAT), .B(G120GAT), .ZN(n409) );
  XNOR2_X1 U470 ( .A(n410), .B(n409), .ZN(n414) );
  XOR2_X1 U471 ( .A(G57GAT), .B(G155GAT), .Z(n412) );
  XNOR2_X1 U472 ( .A(G1GAT), .B(G148GAT), .ZN(n411) );
  XNOR2_X1 U473 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U474 ( .A(n414), .B(n413), .Z(n419) );
  XOR2_X1 U475 ( .A(KEYINPUT89), .B(KEYINPUT4), .Z(n416) );
  NAND2_X1 U476 ( .A1(G225GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U477 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U478 ( .A(KEYINPUT5), .B(n417), .ZN(n418) );
  XNOR2_X1 U479 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U480 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n427), .B(n426), .ZN(n440) );
  XOR2_X1 U482 ( .A(G204GAT), .B(KEYINPUT88), .Z(n429) );
  NAND2_X1 U483 ( .A1(G228GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U484 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U485 ( .A(n430), .B(KEYINPUT23), .Z(n434) );
  XNOR2_X1 U486 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n436) );
  XOR2_X1 U488 ( .A(n436), .B(n435), .Z(n438) );
  XNOR2_X1 U489 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n437) );
  XNOR2_X1 U490 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U491 ( .A(n440), .B(n439), .ZN(n476) );
  NAND2_X1 U492 ( .A1(n289), .A2(n476), .ZN(n441) );
  XNOR2_X1 U493 ( .A(n441), .B(KEYINPUT55), .ZN(n459) );
  XOR2_X1 U494 ( .A(n443), .B(n442), .Z(n445) );
  XNOR2_X1 U495 ( .A(G43GAT), .B(G190GAT), .ZN(n444) );
  XNOR2_X1 U496 ( .A(n445), .B(n444), .ZN(n450) );
  XOR2_X1 U497 ( .A(G15GAT), .B(n446), .Z(n448) );
  NAND2_X1 U498 ( .A1(G227GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U499 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U500 ( .A(n450), .B(n449), .Z(n458) );
  XOR2_X1 U501 ( .A(KEYINPUT20), .B(KEYINPUT85), .Z(n452) );
  XNOR2_X1 U502 ( .A(G99GAT), .B(KEYINPUT84), .ZN(n451) );
  XNOR2_X1 U503 ( .A(n452), .B(n451), .ZN(n456) );
  XOR2_X1 U504 ( .A(G176GAT), .B(G183GAT), .Z(n454) );
  XNOR2_X1 U505 ( .A(KEYINPUT86), .B(KEYINPUT64), .ZN(n453) );
  XNOR2_X1 U506 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U507 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U508 ( .A(n458), .B(n457), .ZN(n538) );
  NAND2_X1 U509 ( .A1(n459), .A2(n538), .ZN(n575) );
  NOR2_X1 U510 ( .A1(n579), .A2(n575), .ZN(n462) );
  INV_X1 U511 ( .A(G169GAT), .ZN(n460) );
  XNOR2_X1 U512 ( .A(n460), .B(KEYINPUT120), .ZN(n461) );
  XNOR2_X1 U513 ( .A(n462), .B(n461), .ZN(G1348GAT) );
  NOR2_X1 U514 ( .A1(n575), .A2(n482), .ZN(n466) );
  XNOR2_X1 U515 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n464) );
  INV_X1 U516 ( .A(G190GAT), .ZN(n463) );
  XNOR2_X1 U517 ( .A(G1GAT), .B(KEYINPUT94), .ZN(n467) );
  XNOR2_X1 U518 ( .A(n467), .B(KEYINPUT93), .ZN(n468) );
  XOR2_X1 U519 ( .A(KEYINPUT34), .B(n468), .Z(n487) );
  NAND2_X1 U520 ( .A1(n379), .A2(n555), .ZN(n499) );
  NAND2_X1 U521 ( .A1(n538), .A2(n529), .ZN(n470) );
  NAND2_X1 U522 ( .A1(n476), .A2(n470), .ZN(n471) );
  XNOR2_X1 U523 ( .A(KEYINPUT25), .B(n471), .ZN(n474) );
  XNOR2_X1 U524 ( .A(KEYINPUT27), .B(n529), .ZN(n477) );
  NOR2_X1 U525 ( .A1(n476), .A2(n538), .ZN(n472) );
  XNOR2_X1 U526 ( .A(n472), .B(KEYINPUT26), .ZN(n578) );
  NAND2_X1 U527 ( .A1(n477), .A2(n578), .ZN(n554) );
  XOR2_X1 U528 ( .A(KEYINPUT92), .B(n554), .Z(n473) );
  NOR2_X1 U529 ( .A1(n474), .A2(n473), .ZN(n475) );
  NOR2_X1 U530 ( .A1(n475), .A2(n551), .ZN(n481) );
  INV_X1 U531 ( .A(n477), .ZN(n478) );
  NOR2_X1 U532 ( .A1(n532), .A2(n478), .ZN(n479) );
  NAND2_X1 U533 ( .A1(n479), .A2(n551), .ZN(n540) );
  NOR2_X1 U534 ( .A1(n538), .A2(n540), .ZN(n480) );
  NOR2_X1 U535 ( .A1(n481), .A2(n480), .ZN(n495) );
  XOR2_X1 U536 ( .A(KEYINPUT16), .B(KEYINPUT83), .Z(n484) );
  NAND2_X1 U537 ( .A1(n562), .A2(n482), .ZN(n483) );
  XNOR2_X1 U538 ( .A(n484), .B(n483), .ZN(n485) );
  OR2_X1 U539 ( .A1(n495), .A2(n485), .ZN(n515) );
  NOR2_X1 U540 ( .A1(n499), .A2(n515), .ZN(n493) );
  NAND2_X1 U541 ( .A1(n493), .A2(n551), .ZN(n486) );
  XNOR2_X1 U542 ( .A(n487), .B(n486), .ZN(G1324GAT) );
  XOR2_X1 U543 ( .A(G8GAT), .B(KEYINPUT95), .Z(n489) );
  NAND2_X1 U544 ( .A1(n493), .A2(n529), .ZN(n488) );
  XNOR2_X1 U545 ( .A(n489), .B(n488), .ZN(G1325GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT35), .B(KEYINPUT96), .Z(n491) );
  NAND2_X1 U547 ( .A1(n493), .A2(n538), .ZN(n490) );
  XNOR2_X1 U548 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U549 ( .A(G15GAT), .B(n492), .ZN(G1326GAT) );
  NAND2_X1 U550 ( .A1(n532), .A2(n493), .ZN(n494) );
  XNOR2_X1 U551 ( .A(n494), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U552 ( .A1(n591), .A2(n495), .ZN(n496) );
  NAND2_X1 U553 ( .A1(n588), .A2(n496), .ZN(n497) );
  XNOR2_X1 U554 ( .A(KEYINPUT37), .B(n497), .ZN(n498) );
  XOR2_X1 U555 ( .A(KEYINPUT98), .B(n498), .Z(n525) );
  NOR2_X1 U556 ( .A1(n499), .A2(n525), .ZN(n500) );
  XNOR2_X1 U557 ( .A(n500), .B(KEYINPUT38), .ZN(n511) );
  NAND2_X1 U558 ( .A1(n511), .A2(n551), .ZN(n503) );
  XNOR2_X1 U559 ( .A(G29GAT), .B(KEYINPUT97), .ZN(n501) );
  XNOR2_X1 U560 ( .A(n501), .B(KEYINPUT39), .ZN(n502) );
  XNOR2_X1 U561 ( .A(n503), .B(n502), .ZN(G1328GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n505) );
  NAND2_X1 U563 ( .A1(n511), .A2(n529), .ZN(n504) );
  XNOR2_X1 U564 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U565 ( .A(G36GAT), .B(n506), .ZN(G1329GAT) );
  XNOR2_X1 U566 ( .A(G43GAT), .B(KEYINPUT101), .ZN(n510) );
  XOR2_X1 U567 ( .A(KEYINPUT40), .B(KEYINPUT102), .Z(n508) );
  NAND2_X1 U568 ( .A1(n538), .A2(n511), .ZN(n507) );
  XNOR2_X1 U569 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U570 ( .A(n510), .B(n509), .ZN(G1330GAT) );
  NAND2_X1 U571 ( .A1(n511), .A2(n532), .ZN(n512) );
  XNOR2_X1 U572 ( .A(n512), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n518) );
  INV_X1 U574 ( .A(n513), .ZN(n569) );
  NOR2_X1 U575 ( .A1(n569), .A2(n555), .ZN(n514) );
  XNOR2_X1 U576 ( .A(n514), .B(KEYINPUT103), .ZN(n526) );
  NOR2_X1 U577 ( .A1(n526), .A2(n515), .ZN(n516) );
  XNOR2_X1 U578 ( .A(KEYINPUT104), .B(n516), .ZN(n522) );
  NAND2_X1 U579 ( .A1(n551), .A2(n522), .ZN(n517) );
  XNOR2_X1 U580 ( .A(n518), .B(n517), .ZN(G1332GAT) );
  XOR2_X1 U581 ( .A(G64GAT), .B(KEYINPUT105), .Z(n520) );
  NAND2_X1 U582 ( .A1(n522), .A2(n529), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n520), .B(n519), .ZN(G1333GAT) );
  NAND2_X1 U584 ( .A1(n522), .A2(n538), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n521), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U586 ( .A(G78GAT), .B(KEYINPUT43), .Z(n524) );
  NAND2_X1 U587 ( .A1(n522), .A2(n532), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n524), .B(n523), .ZN(G1335GAT) );
  NOR2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U590 ( .A(n527), .B(KEYINPUT106), .ZN(n533) );
  NAND2_X1 U591 ( .A1(n533), .A2(n551), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n528), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U593 ( .A1(n533), .A2(n529), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n530), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U595 ( .A1(n533), .A2(n538), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n531), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n537) );
  XOR2_X1 U598 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n535) );
  NAND2_X1 U599 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n537), .B(n536), .ZN(G1339GAT) );
  NAND2_X1 U602 ( .A1(n538), .A2(n552), .ZN(n539) );
  NOR2_X1 U603 ( .A1(n540), .A2(n539), .ZN(n547) );
  NAND2_X1 U604 ( .A1(n555), .A2(n547), .ZN(n541) );
  XNOR2_X1 U605 ( .A(G113GAT), .B(n541), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT49), .Z(n543) );
  NAND2_X1 U607 ( .A1(n547), .A2(n513), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(G1341GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n545) );
  NAND2_X1 U610 ( .A1(n547), .A2(n562), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT51), .B(KEYINPUT114), .Z(n549) );
  NAND2_X1 U614 ( .A1(n547), .A2(n565), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U616 ( .A(G134GAT), .B(n550), .ZN(G1343GAT) );
  XOR2_X1 U617 ( .A(G141GAT), .B(KEYINPUT115), .Z(n557) );
  NAND2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U619 ( .A1(n554), .A2(n553), .ZN(n566) );
  NAND2_X1 U620 ( .A1(n566), .A2(n555), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n557), .B(n556), .ZN(G1344GAT) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n561) );
  XOR2_X1 U623 ( .A(KEYINPUT52), .B(KEYINPUT116), .Z(n559) );
  NAND2_X1 U624 ( .A1(n566), .A2(n513), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(G1345GAT) );
  XOR2_X1 U627 ( .A(G155GAT), .B(KEYINPUT117), .Z(n564) );
  NAND2_X1 U628 ( .A1(n566), .A2(n562), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(G1346GAT) );
  NAND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U631 ( .A(n567), .B(KEYINPUT118), .ZN(n568) );
  XNOR2_X1 U632 ( .A(G162GAT), .B(n568), .ZN(G1347GAT) );
  NOR2_X1 U633 ( .A1(n569), .A2(n575), .ZN(n574) );
  XOR2_X1 U634 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n571) );
  XNOR2_X1 U635 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(KEYINPUT56), .B(n572), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(G1349GAT) );
  NOR2_X1 U639 ( .A1(n588), .A2(n575), .ZN(n577) );
  XNOR2_X1 U640 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(G1350GAT) );
  NAND2_X1 U642 ( .A1(n289), .A2(n578), .ZN(n590) );
  NOR2_X1 U643 ( .A1(n579), .A2(n590), .ZN(n583) );
  XOR2_X1 U644 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n581) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(G1352GAT) );
  NOR2_X1 U648 ( .A1(n590), .A2(n379), .ZN(n587) );
  XOR2_X1 U649 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n585) );
  XNOR2_X1 U650 ( .A(G204GAT), .B(KEYINPUT127), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1353GAT) );
  NOR2_X1 U653 ( .A1(n588), .A2(n590), .ZN(n589) );
  XOR2_X1 U654 ( .A(G211GAT), .B(n589), .Z(G1354GAT) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U656 ( .A(KEYINPUT62), .B(n592), .Z(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

