//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978;
  INV_X1    g000(.A(KEYINPUT96), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT67), .B(G116), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G122), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G122), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT81), .B(G107), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G134), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G143), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT13), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n194), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G128), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(new_n196), .ZN(new_n201));
  XNOR2_X1  g015(.A(new_n198), .B(new_n201), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n193), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT93), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT14), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n206), .B1(new_n190), .B2(G122), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n205), .B1(new_n189), .B2(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n189), .A2(KEYINPUT14), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n189), .A2(new_n205), .A3(new_n207), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G107), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n189), .B(new_n192), .C1(new_n190), .C2(G122), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n200), .A2(new_n196), .A3(G134), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n201), .A2(new_n194), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(KEYINPUT94), .B1(new_n213), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G107), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n220), .B1(new_n210), .B2(new_n211), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT94), .ZN(new_n222));
  NOR3_X1   g036(.A1(new_n221), .A2(new_n222), .A3(new_n217), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n204), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT9), .B(G234), .ZN(new_n225));
  INV_X1    g039(.A(G217), .ZN(new_n226));
  NOR3_X1   g040(.A1(new_n225), .A2(new_n226), .A3(G953), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G902), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n213), .A2(KEYINPUT94), .A3(new_n218), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n222), .B1(new_n221), .B2(new_n217), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n203), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n227), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n228), .A2(new_n229), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G478), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(KEYINPUT15), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n237), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n228), .A2(new_n234), .A3(new_n229), .A4(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G952), .ZN(new_n241));
  AOI211_X1 g055(.A(G953), .B(new_n241), .C1(G234), .C2(G237), .ZN(new_n242));
  INV_X1    g056(.A(G953), .ZN(new_n243));
  AOI211_X1 g057(.A(new_n229), .B(new_n243), .C1(G234), .C2(G237), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT21), .B(G898), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n242), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n238), .A2(new_n240), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(G113), .B(G122), .ZN(new_n249));
  INV_X1    g063(.A(G104), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n249), .B(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G237), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(new_n243), .A3(G214), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n254), .B(new_n199), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G131), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n254), .B(G143), .ZN(new_n257));
  INV_X1    g071(.A(G131), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT17), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n256), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n257), .A2(new_n258), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT17), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G125), .ZN(new_n265));
  NOR3_X1   g079(.A1(new_n265), .A2(KEYINPUT16), .A3(G140), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT74), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(G125), .B(G140), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT74), .B1(new_n269), .B2(KEYINPUT16), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n268), .B1(new_n270), .B2(new_n266), .ZN(new_n271));
  INV_X1    g085(.A(G146), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT75), .ZN(new_n274));
  OAI211_X1 g088(.A(G146), .B(new_n268), .C1(new_n270), .C2(new_n266), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n271), .A2(KEYINPUT75), .A3(new_n272), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n264), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT91), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n262), .A2(new_n279), .A3(KEYINPUT18), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n269), .B(new_n272), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n279), .A2(KEYINPUT18), .A3(G131), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n257), .A2(new_n282), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n280), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n252), .B1(new_n278), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n276), .A2(new_n277), .ZN(new_n286));
  INV_X1    g100(.A(new_n264), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n280), .A2(new_n281), .A3(new_n283), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n251), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(G902), .B1(new_n285), .B2(new_n290), .ZN(new_n291));
  OR2_X1    g105(.A1(new_n291), .A2(KEYINPUT92), .ZN(new_n292));
  INV_X1    g106(.A(G475), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n293), .B1(new_n291), .B2(KEYINPUT92), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n256), .A2(new_n259), .ZN(new_n295));
  XOR2_X1   g109(.A(new_n269), .B(KEYINPUT19), .Z(new_n296));
  OAI211_X1 g110(.A(new_n295), .B(new_n275), .C1(G146), .C2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n251), .B1(new_n297), .B2(new_n289), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n284), .B1(new_n286), .B2(new_n287), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n298), .B1(new_n299), .B2(new_n251), .ZN(new_n300));
  NOR2_X1   g114(.A1(G475), .A2(G902), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(KEYINPUT20), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT20), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n278), .A2(new_n252), .A3(new_n284), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n304), .B(new_n301), .C1(new_n305), .C2(new_n298), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n292), .A2(new_n294), .B1(new_n303), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n248), .A2(KEYINPUT95), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT95), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n303), .A2(new_n306), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n285), .A2(new_n290), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(KEYINPUT92), .A3(new_n229), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G475), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n291), .A2(KEYINPUT92), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n310), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n238), .A2(new_n240), .A3(new_n247), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n309), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n308), .A2(new_n317), .ZN(new_n318));
  AND2_X1   g132(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n319));
  NOR2_X1   g133(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(G143), .B(G146), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(G128), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n272), .A2(G143), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n199), .A2(G146), .ZN(new_n325));
  AOI21_X1  g139(.A(G128), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n199), .A2(KEYINPUT1), .A3(G146), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n323), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n220), .A2(KEYINPUT81), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT81), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G107), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n220), .A2(G104), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT3), .ZN(new_n336));
  AOI21_X1  g150(.A(G101), .B1(new_n250), .B2(G107), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n334), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n335), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n331), .A2(new_n333), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n339), .B1(new_n340), .B2(new_n250), .ZN(new_n341));
  INV_X1    g155(.A(G101), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n338), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT82), .B1(new_n329), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n323), .A2(new_n327), .A3(new_n328), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n335), .B1(new_n192), .B2(G104), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G101), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT82), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n345), .A2(new_n347), .A3(new_n348), .A4(new_n338), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT10), .B1(new_n344), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n324), .A2(new_n325), .ZN(new_n351));
  NAND2_X1  g165(.A1(KEYINPUT0), .A2(G128), .ZN(new_n352));
  OR2_X1    g166(.A1(KEYINPUT0), .A2(G128), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n322), .A2(KEYINPUT0), .A3(G128), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n250), .A2(G107), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n334), .A2(new_n336), .A3(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n342), .A2(KEYINPUT4), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n356), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(G101), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(KEYINPUT4), .A3(new_n338), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n192), .A2(new_n330), .B1(KEYINPUT3), .B2(new_n335), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n364), .A2(new_n337), .B1(new_n346), .B2(G101), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n199), .B(G146), .C1(new_n319), .C2(new_n320), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n323), .A2(new_n327), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n365), .A2(KEYINPUT10), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT11), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n370), .B1(new_n194), .B2(G137), .ZN(new_n371));
  INV_X1    g185(.A(G137), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(KEYINPUT11), .A3(G134), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n194), .A2(G137), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n371), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G131), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n371), .A2(new_n373), .A3(new_n258), .A4(new_n374), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n378), .B(KEYINPUT83), .ZN(new_n379));
  NOR3_X1   g193(.A1(new_n350), .A2(new_n369), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n243), .A2(G227), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(KEYINPUT80), .ZN(new_n382));
  XNOR2_X1  g196(.A(G110), .B(G140), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n382), .B(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n365), .A2(new_n367), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n387), .B1(new_n349), .B2(new_n344), .ZN(new_n388));
  INV_X1    g202(.A(new_n378), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT84), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT12), .B1(new_n378), .B2(new_n390), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n388), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n391), .ZN(new_n393));
  INV_X1    g207(.A(new_n388), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n393), .B1(new_n394), .B2(new_n378), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n386), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n378), .B1(new_n350), .B2(new_n369), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT86), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI211_X1 g213(.A(KEYINPUT86), .B(new_n378), .C1(new_n350), .C2(new_n369), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n380), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n396), .B1(new_n401), .B2(new_n384), .ZN(new_n402));
  INV_X1    g216(.A(G469), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(new_n229), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n403), .A2(new_n229), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  OR3_X1    g220(.A1(new_n350), .A2(new_n369), .A3(new_n379), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(KEYINPUT85), .A3(new_n384), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n399), .A2(new_n400), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT85), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n410), .B1(new_n380), .B2(new_n385), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n407), .B1(new_n395), .B2(new_n392), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n385), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n414), .A3(G469), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n404), .A2(new_n406), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n190), .A2(KEYINPUT67), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT67), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G116), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(new_n420), .A3(G119), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n190), .A2(G119), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(KEYINPUT2), .A2(G113), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT66), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT66), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(KEYINPUT2), .A3(G113), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT2), .ZN(new_n430));
  INV_X1    g244(.A(G113), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n424), .A2(new_n433), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n426), .A2(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(new_n423), .A3(new_n421), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n434), .A2(new_n436), .B1(new_n358), .B2(new_n359), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n421), .A2(KEYINPUT5), .A3(new_n423), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT5), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n431), .B1(new_n422), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n422), .B1(new_n188), .B2(G119), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n438), .A2(new_n440), .B1(new_n441), .B2(new_n435), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n437), .A2(new_n362), .B1(new_n365), .B2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(G110), .B(G122), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n417), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n444), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT87), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n446), .B1(new_n443), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n437), .A2(new_n362), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n365), .A2(new_n442), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n449), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n445), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n361), .A2(KEYINPUT4), .A3(new_n338), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n358), .A2(new_n359), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n424), .A2(new_n433), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n423), .A2(new_n421), .B1(new_n429), .B2(new_n432), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n450), .B1(new_n453), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT87), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n443), .A2(new_n447), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n459), .A2(new_n460), .A3(new_n417), .A4(new_n446), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n452), .A2(KEYINPUT88), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT88), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n463), .B(new_n445), .C1(new_n448), .C2(new_n451), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n324), .A2(new_n325), .A3(G128), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n326), .B1(new_n466), .B2(new_n321), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(new_n265), .A3(new_n366), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n356), .A2(G125), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n243), .A2(G224), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n470), .B(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n465), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(G210), .B1(G237), .B2(G902), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT7), .A4(new_n471), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT7), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(KEYINPUT89), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT89), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n471), .B1(new_n479), .B2(KEYINPUT7), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n470), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT90), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n442), .B(new_n343), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n444), .B(KEYINPUT8), .Z(new_n484));
  OAI221_X1 g298(.A(new_n476), .B1(new_n481), .B2(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n481), .A2(new_n482), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n486), .B1(new_n458), .B2(new_n446), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n229), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n474), .A2(new_n475), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n475), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n472), .B1(new_n462), .B2(new_n464), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n491), .B1(new_n492), .B2(new_n488), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(G214), .B1(G237), .B2(G902), .ZN(new_n495));
  OAI21_X1  g309(.A(G221), .B1(new_n225), .B2(G902), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n416), .A2(new_n494), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n187), .B1(new_n318), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n226), .B1(G234), .B2(new_n229), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n229), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(KEYINPUT79), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT22), .B(G137), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n243), .A2(G221), .A3(G234), .ZN(new_n505));
  XOR2_X1   g319(.A(new_n504), .B(new_n505), .Z(new_n506));
  INV_X1    g320(.A(G119), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT73), .B1(new_n507), .B2(G128), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n508), .A2(KEYINPUT23), .B1(new_n507), .B2(G128), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n509), .B1(KEYINPUT23), .B2(new_n508), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(G110), .ZN(new_n511));
  XOR2_X1   g325(.A(KEYINPUT24), .B(G110), .Z(new_n512));
  XNOR2_X1  g326(.A(G119), .B(G128), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(KEYINPUT72), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n276), .A2(new_n277), .A3(new_n511), .A4(new_n515), .ZN(new_n516));
  XOR2_X1   g330(.A(KEYINPUT76), .B(G110), .Z(new_n517));
  OAI22_X1  g331(.A1(new_n510), .A2(new_n517), .B1(new_n513), .B2(new_n512), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n269), .A2(new_n272), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(new_n275), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n506), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n516), .A2(new_n520), .A3(new_n506), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n524), .A2(KEYINPUT78), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(KEYINPUT78), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n503), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n528), .B1(new_n524), .B2(G902), .ZN(new_n529));
  INV_X1    g343(.A(new_n528), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n522), .A2(new_n229), .A3(new_n523), .A4(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n500), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  OR2_X1    g346(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(G472), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n378), .A2(new_n355), .A3(new_n354), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n194), .A2(G137), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n372), .A2(G134), .ZN(new_n537));
  OAI21_X1  g351(.A(G131), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n377), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n367), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n455), .A2(new_n456), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(new_n535), .A3(new_n540), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(KEYINPUT70), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT70), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n541), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n546), .A2(KEYINPUT28), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n253), .A2(new_n243), .A3(G210), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(KEYINPUT27), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT26), .B(G101), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n551), .B(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT28), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n545), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n549), .A2(KEYINPUT29), .A3(new_n553), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n229), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n356), .B1(new_n377), .B2(new_n376), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n377), .A2(new_n538), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n559), .B1(new_n467), .B2(new_n366), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT30), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(KEYINPUT64), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT64), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n377), .A2(new_n538), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n562), .A2(new_n367), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT30), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n566), .A3(new_n535), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n543), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n545), .ZN(new_n570));
  INV_X1    g384(.A(new_n553), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(KEYINPUT68), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT68), .ZN(new_n573));
  INV_X1    g387(.A(new_n545), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n574), .B1(new_n568), .B2(new_n543), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n573), .B1(new_n575), .B2(new_n553), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n565), .A2(new_n535), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n543), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n542), .A2(new_n535), .A3(KEYINPUT28), .A4(new_n540), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n555), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT29), .B1(new_n580), .B2(new_n553), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n572), .A2(new_n576), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n557), .B1(new_n582), .B2(KEYINPUT69), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT69), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n572), .A2(new_n581), .A3(new_n576), .A4(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n534), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT31), .B1(new_n575), .B2(new_n553), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n542), .B1(new_n561), .B2(new_n567), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT31), .ZN(new_n589));
  NOR4_X1   g403(.A1(new_n588), .A2(new_n589), .A3(new_n571), .A4(new_n574), .ZN(new_n590));
  OAI22_X1  g404(.A1(new_n587), .A2(new_n590), .B1(new_n553), .B2(new_n580), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT32), .ZN(new_n592));
  NOR2_X1   g406(.A1(G472), .A2(G902), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n592), .B1(new_n591), .B2(new_n593), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n586), .A2(KEYINPUT71), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT71), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n583), .A2(new_n585), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n598), .B1(new_n599), .B2(new_n534), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n533), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n494), .ZN(new_n602));
  INV_X1    g416(.A(new_n495), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n416), .A2(new_n496), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n308), .A2(new_n317), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n604), .A2(new_n605), .A3(new_n606), .A4(KEYINPUT96), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n498), .A2(new_n601), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G101), .ZN(G3));
  NAND2_X1  g423(.A1(new_n235), .A2(new_n236), .ZN(new_n610));
  OR3_X1    g424(.A1(new_n232), .A2(KEYINPUT100), .A3(new_n227), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n227), .B1(new_n232), .B2(KEYINPUT100), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(KEYINPUT33), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT99), .B(KEYINPUT33), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n228), .A2(new_n234), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n229), .A2(G478), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n610), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n315), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n619), .A2(new_n246), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT98), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n490), .A2(KEYINPUT97), .A3(new_n493), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n495), .B1(new_n490), .B2(KEYINPUT97), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n492), .A2(new_n491), .A3(new_n488), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT97), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n603), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n490), .A2(KEYINPUT97), .A3(new_n493), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(new_n628), .A3(KEYINPUT98), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n620), .A2(new_n624), .A3(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n416), .A2(new_n496), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n591), .A2(new_n229), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(G472), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n591), .A2(new_n593), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n632), .A2(new_n636), .A3(new_n533), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n631), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT34), .B(G104), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  AND3_X1   g454(.A1(new_n627), .A2(new_n628), .A3(KEYINPUT98), .ZN(new_n641));
  AOI21_X1  g455(.A(KEYINPUT98), .B1(new_n627), .B2(new_n628), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n246), .B1(new_n292), .B2(new_n294), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n238), .A2(new_n240), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n310), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n303), .A2(KEYINPUT101), .A3(new_n306), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n644), .A2(new_n645), .A3(new_n647), .A4(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n643), .A2(new_n637), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT35), .B(G107), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  NAND2_X1  g468(.A1(new_n516), .A2(new_n520), .ZN(new_n655));
  INV_X1    g469(.A(new_n506), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n656), .A2(KEYINPUT36), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n655), .B(new_n657), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n658), .A2(new_n502), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n532), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n636), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n498), .A2(new_n607), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT37), .B(G110), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G12));
  NAND2_X1  g478(.A1(new_n647), .A2(new_n648), .ZN(new_n665));
  INV_X1    g479(.A(new_n645), .ZN(new_n666));
  INV_X1    g480(.A(new_n242), .ZN(new_n667));
  INV_X1    g481(.A(new_n244), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT103), .B(G900), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT104), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n671), .B1(new_n313), .B2(new_n314), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n665), .A2(new_n666), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n660), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n605), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n597), .A2(new_n600), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n675), .A2(new_n643), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(new_n195), .ZN(G30));
  XOR2_X1   g492(.A(new_n494), .B(KEYINPUT38), .Z(new_n679));
  NOR4_X1   g493(.A1(new_n679), .A2(new_n307), .A3(new_n666), .A4(new_n603), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n570), .A2(new_n553), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n546), .A2(new_n548), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n229), .B1(new_n683), .B2(new_n553), .ZN(new_n684));
  OAI21_X1  g498(.A(G472), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n594), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n685), .B1(new_n686), .B2(new_n595), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n660), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n671), .B(KEYINPUT39), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n605), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n688), .B1(new_n690), .B2(KEYINPUT40), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n680), .B(new_n691), .C1(KEYINPUT40), .C2(new_n690), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G143), .ZN(G45));
  AND2_X1   g507(.A1(new_n643), .A2(new_n676), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n618), .A2(new_n315), .A3(new_n671), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n695), .A2(new_n632), .A3(new_n660), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G146), .ZN(G48));
  INV_X1    g512(.A(new_n402), .ZN(new_n699));
  OAI21_X1  g513(.A(G469), .B1(new_n699), .B2(G902), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(new_n496), .A3(new_n404), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT105), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n700), .A2(new_n703), .A3(new_n496), .A4(new_n404), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n631), .A2(new_n601), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT41), .B(G113), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G15));
  NAND4_X1  g522(.A1(new_n705), .A2(new_n601), .A3(new_n643), .A4(new_n651), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G116), .ZN(G18));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n711));
  INV_X1    g525(.A(new_n701), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n624), .A2(new_n712), .A3(new_n629), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT106), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT106), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n624), .A2(new_n712), .A3(new_n629), .A4(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n660), .B1(new_n308), .B2(new_n317), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n676), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n711), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  AOI211_X1 g535(.A(KEYINPUT107), .B(new_n719), .C1(new_n714), .C2(new_n716), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n507), .ZN(G21));
  XNOR2_X1  g538(.A(KEYINPUT108), .B(G472), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n633), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n587), .A2(new_n590), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n553), .B1(new_n549), .B2(new_n555), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n593), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n533), .A2(new_n246), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(new_n702), .A3(new_n704), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n666), .A2(new_n307), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n624), .A2(new_n629), .A3(new_n733), .ZN(new_n734));
  OR2_X1    g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  INV_X1    g550(.A(new_n730), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n674), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n738), .A2(new_n695), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n715), .B1(new_n643), .B2(new_n712), .ZN(new_n740));
  INV_X1    g554(.A(new_n716), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G125), .ZN(G27));
  NOR3_X1   g557(.A1(new_n632), .A2(new_n603), .A3(new_n494), .ZN(new_n744));
  INV_X1    g558(.A(new_n695), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n601), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT42), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n601), .A2(new_n744), .A3(KEYINPUT42), .A4(new_n745), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G131), .ZN(G33));
  NAND3_X1  g565(.A1(new_n601), .A2(new_n744), .A3(new_n673), .ZN(new_n752));
  XOR2_X1   g566(.A(KEYINPUT109), .B(G134), .Z(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(G36));
  NAND2_X1  g568(.A1(new_n674), .A2(new_n636), .ZN(new_n755));
  XOR2_X1   g569(.A(new_n755), .B(KEYINPUT111), .Z(new_n756));
  NAND2_X1  g570(.A1(new_n618), .A2(new_n307), .ZN(new_n757));
  XOR2_X1   g571(.A(new_n757), .B(KEYINPUT43), .Z(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n494), .A2(new_n603), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n412), .A2(KEYINPUT45), .A3(new_n414), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT45), .B1(new_n412), .B2(new_n414), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n764), .A2(new_n765), .A3(new_n403), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n405), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT110), .ZN(new_n768));
  OR3_X1    g582(.A1(new_n767), .A2(new_n768), .A3(KEYINPUT46), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n768), .B1(new_n767), .B2(KEYINPUT46), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n402), .A2(new_n403), .A3(new_n229), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n771), .B1(new_n767), .B2(KEYINPUT46), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(new_n496), .A3(new_n689), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n759), .A2(new_n760), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n763), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(new_n372), .ZN(G39));
  AND2_X1   g591(.A1(new_n773), .A2(new_n496), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n778), .A2(KEYINPUT47), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(KEYINPUT47), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n676), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n782), .A2(new_n533), .A3(new_n745), .A4(new_n762), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G140), .ZN(G42));
  INV_X1    g600(.A(new_n496), .ZN(new_n787));
  OR3_X1    g601(.A1(new_n533), .A2(new_n603), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n700), .A2(new_n404), .ZN(new_n789));
  AOI211_X1 g603(.A(new_n757), .B(new_n788), .C1(KEYINPUT49), .C2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n687), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n789), .A2(KEYINPUT49), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n790), .A2(new_n679), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n758), .A2(new_n242), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n701), .A2(new_n603), .A3(new_n494), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n601), .A3(new_n795), .ZN(new_n796));
  XOR2_X1   g610(.A(new_n796), .B(KEYINPUT48), .Z(new_n797));
  NOR2_X1   g611(.A1(new_n533), .A2(new_n730), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n794), .A2(new_n717), .A3(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n533), .A2(new_n687), .A3(new_n667), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g615(.A(new_n801), .B(KEYINPUT120), .Z(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  OAI211_X1 g617(.A(G952), .B(new_n243), .C1(new_n803), .C2(new_n619), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n797), .A2(new_n799), .A3(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n701), .A2(new_n495), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n794), .A2(new_n679), .A3(new_n798), .A4(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT50), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n807), .A2(new_n808), .A3(KEYINPUT50), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT118), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n794), .A2(new_n674), .A3(new_n737), .A4(new_n795), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT119), .ZN(new_n817));
  OR3_X1    g631(.A1(new_n803), .A2(new_n315), .A3(new_n618), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n815), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n794), .A2(new_n798), .A3(new_n762), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n820), .B(KEYINPUT114), .Z(new_n821));
  OR2_X1    g635(.A1(new_n789), .A2(KEYINPUT115), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n789), .A2(KEYINPUT115), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(new_n787), .A3(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(KEYINPUT116), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n779), .A2(new_n780), .A3(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n821), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n813), .B1(new_n814), .B2(new_n828), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n819), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  AND4_X1   g644(.A1(new_n812), .A2(new_n818), .A3(new_n811), .A4(new_n817), .ZN(new_n831));
  INV_X1    g645(.A(new_n824), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n821), .B1(new_n781), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n828), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n805), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n706), .A2(new_n709), .A3(new_n735), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n717), .A2(new_n720), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT107), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n717), .A2(new_n711), .A3(new_n720), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n694), .A2(new_n675), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n415), .A2(new_n406), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n496), .B(new_n671), .C1(new_n771), .C2(new_n843), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n688), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n842), .B1(new_n734), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n688), .A2(new_n844), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n643), .A2(KEYINPUT112), .A3(new_n733), .A4(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n742), .A2(new_n841), .A3(new_n697), .A4(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT52), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n677), .B1(new_n717), .B2(new_n739), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT52), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n852), .A2(new_n853), .A3(new_n697), .A4(new_n849), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n748), .A2(new_n749), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n619), .B1(new_n315), .B2(new_n666), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n637), .A2(new_n247), .A3(new_n604), .A4(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n608), .A2(new_n662), .A3(new_n857), .ZN(new_n858));
  NOR4_X1   g672(.A1(new_n660), .A2(new_n665), .A3(new_n672), .A4(new_n645), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n739), .B1(new_n676), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n744), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n752), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n855), .A2(new_n858), .A3(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n840), .A2(new_n851), .A3(new_n854), .A4(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n852), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT53), .B1(new_n867), .B2(KEYINPUT52), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n866), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(KEYINPUT54), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n601), .A2(new_n702), .A3(new_n704), .ZN(new_n871));
  OAI22_X1  g685(.A1(new_n871), .A2(new_n630), .B1(new_n734), .B2(new_n732), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n643), .A2(new_n651), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n873), .A2(new_n871), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n875), .B1(new_n721), .B2(new_n722), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n608), .A2(new_n662), .A3(new_n857), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n860), .A2(new_n861), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n877), .A2(new_n878), .A3(new_n750), .A4(new_n752), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n865), .B1(new_n867), .B2(KEYINPUT52), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n880), .A2(new_n854), .A3(new_n851), .A4(new_n881), .ZN(new_n882));
  XOR2_X1   g696(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n883));
  NAND3_X1  g697(.A1(new_n866), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n870), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n835), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(G952), .A2(G953), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n793), .B1(new_n886), .B2(new_n887), .ZN(G75));
  AOI21_X1  g702(.A(new_n229), .B1(new_n866), .B2(new_n882), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(G210), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT56), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n465), .A2(new_n473), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n492), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT55), .Z(new_n895));
  AND2_X1   g709(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n892), .A2(new_n895), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n243), .A2(G952), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(G51));
  AND2_X1   g713(.A1(new_n889), .A2(new_n766), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n866), .A2(new_n882), .ZN(new_n901));
  INV_X1    g715(.A(new_n883), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n884), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n405), .B(KEYINPUT57), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n699), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n900), .B1(new_n906), .B2(KEYINPUT121), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT121), .ZN(new_n908));
  INV_X1    g722(.A(new_n905), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n909), .B1(new_n903), .B2(new_n884), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n910), .B2(new_n699), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n898), .B1(new_n907), .B2(new_n911), .ZN(G54));
  NAND3_X1  g726(.A1(new_n889), .A2(KEYINPUT58), .A3(G475), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n913), .A2(new_n300), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n913), .A2(new_n300), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n914), .A2(new_n915), .A3(new_n898), .ZN(G60));
  INV_X1    g730(.A(new_n616), .ZN(new_n917));
  NAND2_X1  g731(.A1(G478), .A2(G902), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT59), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n917), .B1(new_n885), .B2(new_n919), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n904), .A2(new_n917), .A3(new_n919), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n920), .A2(new_n921), .A3(new_n898), .ZN(G63));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT122), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT60), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n901), .A2(new_n658), .A3(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n898), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT61), .B1(new_n928), .B2(KEYINPUT123), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n901), .A2(new_n925), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n930), .A2(new_n525), .A3(new_n526), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n931), .A2(new_n927), .A3(new_n926), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n929), .B(new_n932), .ZN(G66));
  INV_X1    g747(.A(new_n245), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n243), .B1(new_n934), .B2(G224), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n840), .A2(new_n877), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n935), .B1(new_n936), .B2(new_n243), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n462), .B(new_n464), .C1(G898), .C2(new_n243), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT124), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n937), .B(new_n939), .ZN(G69));
  XOR2_X1   g754(.A(new_n568), .B(new_n296), .Z(new_n941));
  NAND3_X1  g755(.A1(new_n643), .A2(new_n601), .A3(new_n733), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n752), .B1(new_n774), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n776), .A2(new_n943), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n852), .A2(new_n697), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n945), .A2(new_n750), .ZN(new_n946));
  AND4_X1   g760(.A1(new_n243), .A2(new_n944), .A3(new_n785), .A4(new_n946), .ZN(new_n947));
  AND2_X1   g761(.A1(G900), .A2(G953), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n941), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n945), .A2(new_n692), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n950), .A2(KEYINPUT62), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(KEYINPUT62), .ZN(new_n952));
  AND4_X1   g766(.A1(new_n601), .A2(new_n744), .A3(new_n689), .A4(new_n856), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n776), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n951), .A2(new_n785), .A3(new_n952), .A4(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n941), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n955), .A2(new_n243), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n949), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n243), .B1(G227), .B2(G900), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT125), .Z(new_n960));
  XNOR2_X1  g774(.A(new_n958), .B(new_n960), .ZN(G72));
  NAND2_X1  g775(.A1(G472), .A2(G902), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT63), .Z(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(new_n955), .B2(new_n936), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT126), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n964), .A2(new_n965), .A3(new_n682), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n965), .B1(new_n964), .B2(new_n682), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n936), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n969), .A2(new_n944), .A3(new_n785), .A4(new_n946), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT127), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n970), .A2(new_n971), .A3(new_n963), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n971), .B1(new_n970), .B2(new_n963), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n571), .B(new_n575), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n572), .B(new_n576), .C1(new_n571), .C2(new_n570), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n869), .A2(new_n963), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n975), .A2(new_n927), .A3(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n968), .A2(new_n978), .ZN(G57));
endmodule


