

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U553 ( .A1(G2105), .A2(G2104), .ZN(n519) );
  NAND2_X2 U554 ( .A1(n592), .A2(n722), .ZN(n648) );
  AND2_X2 U555 ( .A1(n523), .A2(G2104), .ZN(n848) );
  INV_X1 U556 ( .A(KEYINPUT105), .ZN(n682) );
  NOR2_X1 U557 ( .A1(G164), .A2(G1384), .ZN(n722) );
  AND2_X1 U558 ( .A1(n539), .A2(n538), .ZN(n518) );
  NOR2_X1 U559 ( .A1(n610), .A2(n609), .ZN(n624) );
  INV_X1 U560 ( .A(KEYINPUT31), .ZN(n655) );
  XNOR2_X1 U561 ( .A(n655), .B(KEYINPUT102), .ZN(n656) );
  XNOR2_X1 U562 ( .A(n657), .B(n656), .ZN(n658) );
  NOR2_X1 U563 ( .A1(n671), .A2(n673), .ZN(n674) );
  XNOR2_X1 U564 ( .A(n683), .B(n682), .ZN(n684) );
  NAND2_X1 U565 ( .A1(G8), .A2(n648), .ZN(n697) );
  NOR2_X2 U566 ( .A1(G2104), .A2(n523), .ZN(n873) );
  NOR2_X1 U567 ( .A1(G651), .A2(n548), .ZN(n786) );
  NOR2_X1 U568 ( .A1(n606), .A2(n605), .ZN(n967) );
  NOR2_X1 U569 ( .A1(n527), .A2(n526), .ZN(G160) );
  XOR2_X2 U570 ( .A(KEYINPUT17), .B(n519), .Z(n870) );
  NAND2_X1 U571 ( .A1(n870), .A2(G137), .ZN(n522) );
  INV_X1 U572 ( .A(G2105), .ZN(n523) );
  NAND2_X1 U573 ( .A1(G101), .A2(n848), .ZN(n520) );
  XOR2_X1 U574 ( .A(KEYINPUT23), .B(n520), .Z(n521) );
  NAND2_X1 U575 ( .A1(n522), .A2(n521), .ZN(n527) );
  NAND2_X1 U576 ( .A1(G125), .A2(n873), .ZN(n525) );
  AND2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n875) );
  NAND2_X1 U578 ( .A1(G113), .A2(n875), .ZN(n524) );
  NAND2_X1 U579 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X2 U580 ( .A1(G651), .A2(G543), .ZN(n780) );
  NAND2_X1 U581 ( .A1(G86), .A2(n780), .ZN(n530) );
  INV_X1 U582 ( .A(G651), .ZN(n531) );
  OR2_X1 U583 ( .A1(G543), .A2(n531), .ZN(n528) );
  XNOR2_X2 U584 ( .A(KEYINPUT1), .B(n528), .ZN(n784) );
  NAND2_X1 U585 ( .A1(G61), .A2(n784), .ZN(n529) );
  NAND2_X1 U586 ( .A1(n530), .A2(n529), .ZN(n534) );
  XOR2_X1 U587 ( .A(G543), .B(KEYINPUT0), .Z(n548) );
  NOR2_X1 U588 ( .A1(n548), .A2(n531), .ZN(n781) );
  NAND2_X1 U589 ( .A1(n781), .A2(G73), .ZN(n532) );
  XOR2_X1 U590 ( .A(KEYINPUT2), .B(n532), .Z(n533) );
  NOR2_X1 U591 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U592 ( .A(KEYINPUT79), .B(n535), .Z(n537) );
  NAND2_X1 U593 ( .A1(n786), .A2(G48), .ZN(n536) );
  NAND2_X1 U594 ( .A1(n537), .A2(n536), .ZN(G305) );
  NAND2_X1 U595 ( .A1(n870), .A2(G138), .ZN(n543) );
  NAND2_X1 U596 ( .A1(G126), .A2(n873), .ZN(n539) );
  NAND2_X1 U597 ( .A1(G114), .A2(n875), .ZN(n538) );
  NAND2_X1 U598 ( .A1(n848), .A2(G102), .ZN(n540) );
  XNOR2_X1 U599 ( .A(n540), .B(KEYINPUT88), .ZN(n541) );
  AND2_X1 U600 ( .A1(n518), .A2(n541), .ZN(n542) );
  AND2_X1 U601 ( .A1(n543), .A2(n542), .ZN(G164) );
  NAND2_X1 U602 ( .A1(G49), .A2(n786), .ZN(n545) );
  NAND2_X1 U603 ( .A1(G74), .A2(G651), .ZN(n544) );
  NAND2_X1 U604 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U605 ( .A(KEYINPUT78), .B(n546), .ZN(n547) );
  NOR2_X1 U606 ( .A1(n784), .A2(n547), .ZN(n550) );
  NAND2_X1 U607 ( .A1(n548), .A2(G87), .ZN(n549) );
  NAND2_X1 U608 ( .A1(n550), .A2(n549), .ZN(G288) );
  NAND2_X1 U609 ( .A1(G78), .A2(n781), .ZN(n551) );
  XOR2_X1 U610 ( .A(KEYINPUT66), .B(n551), .Z(n556) );
  NAND2_X1 U611 ( .A1(G53), .A2(n786), .ZN(n553) );
  NAND2_X1 U612 ( .A1(G65), .A2(n784), .ZN(n552) );
  NAND2_X1 U613 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U614 ( .A(KEYINPUT67), .B(n554), .Z(n555) );
  NOR2_X1 U615 ( .A1(n556), .A2(n555), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n780), .A2(G91), .ZN(n557) );
  NAND2_X1 U617 ( .A1(n558), .A2(n557), .ZN(G299) );
  NAND2_X1 U618 ( .A1(G52), .A2(n786), .ZN(n560) );
  NAND2_X1 U619 ( .A1(G64), .A2(n784), .ZN(n559) );
  NAND2_X1 U620 ( .A1(n560), .A2(n559), .ZN(n566) );
  NAND2_X1 U621 ( .A1(n781), .A2(G77), .ZN(n561) );
  XOR2_X1 U622 ( .A(KEYINPUT65), .B(n561), .Z(n563) );
  NAND2_X1 U623 ( .A1(n780), .A2(G90), .ZN(n562) );
  NAND2_X1 U624 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U625 ( .A(KEYINPUT9), .B(n564), .Z(n565) );
  NOR2_X1 U626 ( .A1(n566), .A2(n565), .ZN(G171) );
  XNOR2_X1 U627 ( .A(KEYINPUT7), .B(KEYINPUT74), .ZN(n578) );
  NAND2_X1 U628 ( .A1(n780), .A2(G89), .ZN(n567) );
  XNOR2_X1 U629 ( .A(n567), .B(KEYINPUT4), .ZN(n569) );
  NAND2_X1 U630 ( .A1(G76), .A2(n781), .ZN(n568) );
  NAND2_X1 U631 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U632 ( .A(KEYINPUT5), .B(n570), .ZN(n576) );
  NAND2_X1 U633 ( .A1(n784), .A2(G63), .ZN(n571) );
  XOR2_X1 U634 ( .A(KEYINPUT73), .B(n571), .Z(n573) );
  NAND2_X1 U635 ( .A1(n786), .A2(G51), .ZN(n572) );
  NAND2_X1 U636 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U637 ( .A(KEYINPUT6), .B(n574), .Z(n575) );
  NAND2_X1 U638 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U639 ( .A(n578), .B(n577), .ZN(G168) );
  XOR2_X1 U640 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U641 ( .A1(G88), .A2(n780), .ZN(n580) );
  NAND2_X1 U642 ( .A1(G75), .A2(n781), .ZN(n579) );
  NAND2_X1 U643 ( .A1(n580), .A2(n579), .ZN(n584) );
  NAND2_X1 U644 ( .A1(G50), .A2(n786), .ZN(n582) );
  NAND2_X1 U645 ( .A1(G62), .A2(n784), .ZN(n581) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U647 ( .A1(n584), .A2(n583), .ZN(G166) );
  XNOR2_X1 U648 ( .A(KEYINPUT89), .B(G166), .ZN(G303) );
  NAND2_X1 U649 ( .A1(G85), .A2(n780), .ZN(n586) );
  NAND2_X1 U650 ( .A1(G72), .A2(n781), .ZN(n585) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U652 ( .A1(G60), .A2(n784), .ZN(n587) );
  XOR2_X1 U653 ( .A(KEYINPUT64), .B(n587), .Z(n588) );
  NOR2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U655 ( .A1(n786), .A2(G47), .ZN(n590) );
  NAND2_X1 U656 ( .A1(n591), .A2(n590), .ZN(G290) );
  XOR2_X1 U657 ( .A(G1981), .B(G305), .Z(n982) );
  NAND2_X1 U658 ( .A1(G160), .A2(G40), .ZN(n721) );
  INV_X1 U659 ( .A(n721), .ZN(n592) );
  NOR2_X1 U660 ( .A1(G1976), .A2(G288), .ZN(n678) );
  NAND2_X1 U661 ( .A1(n678), .A2(KEYINPUT33), .ZN(n593) );
  NOR2_X1 U662 ( .A1(n697), .A2(n593), .ZN(n687) );
  INV_X1 U663 ( .A(n648), .ZN(n639) );
  NAND2_X1 U664 ( .A1(G1996), .A2(n639), .ZN(n594) );
  XNOR2_X1 U665 ( .A(KEYINPUT26), .B(n594), .ZN(n607) );
  NAND2_X1 U666 ( .A1(G56), .A2(n784), .ZN(n595) );
  XNOR2_X1 U667 ( .A(n595), .B(KEYINPUT14), .ZN(n598) );
  NAND2_X1 U668 ( .A1(G43), .A2(n786), .ZN(n596) );
  XNOR2_X1 U669 ( .A(n596), .B(KEYINPUT70), .ZN(n597) );
  NAND2_X1 U670 ( .A1(n598), .A2(n597), .ZN(n606) );
  XOR2_X1 U671 ( .A(KEYINPUT12), .B(KEYINPUT69), .Z(n600) );
  NAND2_X1 U672 ( .A1(G81), .A2(n780), .ZN(n599) );
  XNOR2_X1 U673 ( .A(n600), .B(n599), .ZN(n601) );
  XNOR2_X1 U674 ( .A(KEYINPUT68), .B(n601), .ZN(n603) );
  NAND2_X1 U675 ( .A1(n781), .A2(G68), .ZN(n602) );
  NAND2_X1 U676 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U677 ( .A(KEYINPUT13), .B(n604), .Z(n605) );
  NAND2_X1 U678 ( .A1(n607), .A2(n967), .ZN(n610) );
  NAND2_X1 U679 ( .A1(G1341), .A2(n648), .ZN(n608) );
  XNOR2_X1 U680 ( .A(KEYINPUT99), .B(n608), .ZN(n609) );
  NAND2_X1 U681 ( .A1(G54), .A2(n786), .ZN(n612) );
  NAND2_X1 U682 ( .A1(G66), .A2(n784), .ZN(n611) );
  NAND2_X1 U683 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U684 ( .A1(G92), .A2(n780), .ZN(n614) );
  NAND2_X1 U685 ( .A1(G79), .A2(n781), .ZN(n613) );
  NAND2_X1 U686 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U687 ( .A1(n616), .A2(n615), .ZN(n618) );
  XNOR2_X1 U688 ( .A(KEYINPUT72), .B(KEYINPUT15), .ZN(n617) );
  XNOR2_X1 U689 ( .A(n618), .B(n617), .ZN(n892) );
  INV_X1 U690 ( .A(n892), .ZN(n975) );
  NAND2_X1 U691 ( .A1(n624), .A2(n975), .ZN(n623) );
  XNOR2_X2 U692 ( .A(n648), .B(KEYINPUT97), .ZN(n641) );
  NAND2_X1 U693 ( .A1(G2067), .A2(n641), .ZN(n619) );
  XNOR2_X1 U694 ( .A(n619), .B(KEYINPUT100), .ZN(n621) );
  NAND2_X1 U695 ( .A1(G1348), .A2(n648), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U697 ( .A1(n623), .A2(n622), .ZN(n626) );
  OR2_X1 U698 ( .A1(n624), .A2(n975), .ZN(n625) );
  NAND2_X1 U699 ( .A1(n626), .A2(n625), .ZN(n631) );
  NAND2_X1 U700 ( .A1(n641), .A2(G2072), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n627), .B(KEYINPUT27), .ZN(n629) );
  INV_X1 U702 ( .A(G1956), .ZN(n997) );
  NOR2_X1 U703 ( .A1(n997), .A2(n641), .ZN(n628) );
  NOR2_X1 U704 ( .A1(n629), .A2(n628), .ZN(n632) );
  INV_X1 U705 ( .A(G299), .ZN(n798) );
  NAND2_X1 U706 ( .A1(n632), .A2(n798), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n636) );
  NOR2_X1 U708 ( .A1(n632), .A2(n798), .ZN(n633) );
  XNOR2_X1 U709 ( .A(n633), .B(KEYINPUT28), .ZN(n634) );
  INV_X1 U710 ( .A(n634), .ZN(n635) );
  NAND2_X1 U711 ( .A1(n636), .A2(n635), .ZN(n638) );
  XNOR2_X1 U712 ( .A(KEYINPUT29), .B(KEYINPUT101), .ZN(n637) );
  XNOR2_X1 U713 ( .A(n638), .B(n637), .ZN(n646) );
  NOR2_X1 U714 ( .A1(n639), .A2(G1961), .ZN(n640) );
  XOR2_X1 U715 ( .A(KEYINPUT96), .B(n640), .Z(n643) );
  XNOR2_X1 U716 ( .A(KEYINPUT25), .B(G2078), .ZN(n952) );
  NAND2_X1 U717 ( .A1(n641), .A2(n952), .ZN(n642) );
  NAND2_X1 U718 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U719 ( .A1(G171), .A2(n647), .ZN(n644) );
  XNOR2_X1 U720 ( .A(n644), .B(KEYINPUT98), .ZN(n645) );
  NAND2_X1 U721 ( .A1(n646), .A2(n645), .ZN(n659) );
  NOR2_X1 U722 ( .A1(G171), .A2(n647), .ZN(n654) );
  NOR2_X1 U723 ( .A1(G1966), .A2(n697), .ZN(n671) );
  NOR2_X1 U724 ( .A1(G2084), .A2(n648), .ZN(n669) );
  INV_X1 U725 ( .A(n669), .ZN(n649) );
  NAND2_X1 U726 ( .A1(G8), .A2(n649), .ZN(n650) );
  OR2_X1 U727 ( .A1(n671), .A2(n650), .ZN(n651) );
  XNOR2_X1 U728 ( .A(KEYINPUT30), .B(n651), .ZN(n652) );
  NOR2_X1 U729 ( .A1(n652), .A2(G168), .ZN(n653) );
  NOR2_X1 U730 ( .A1(n654), .A2(n653), .ZN(n657) );
  NAND2_X1 U731 ( .A1(n659), .A2(n658), .ZN(n672) );
  NAND2_X1 U732 ( .A1(n672), .A2(G286), .ZN(n666) );
  NOR2_X1 U733 ( .A1(G1971), .A2(n697), .ZN(n660) );
  XOR2_X1 U734 ( .A(KEYINPUT103), .B(n660), .Z(n662) );
  NOR2_X1 U735 ( .A1(G2090), .A2(n648), .ZN(n661) );
  NOR2_X1 U736 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U737 ( .A1(n663), .A2(G303), .ZN(n664) );
  XNOR2_X1 U738 ( .A(n664), .B(KEYINPUT104), .ZN(n665) );
  NAND2_X1 U739 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U740 ( .A1(n667), .A2(G8), .ZN(n668) );
  XNOR2_X1 U741 ( .A(n668), .B(KEYINPUT32), .ZN(n690) );
  NAND2_X1 U742 ( .A1(G8), .A2(n669), .ZN(n670) );
  XOR2_X1 U743 ( .A(KEYINPUT95), .B(n670), .Z(n675) );
  INV_X1 U744 ( .A(n672), .ZN(n673) );
  NAND2_X1 U745 ( .A1(n675), .A2(n674), .ZN(n689) );
  NAND2_X1 U746 ( .A1(G1976), .A2(G288), .ZN(n980) );
  AND2_X1 U747 ( .A1(n689), .A2(n980), .ZN(n676) );
  NAND2_X1 U748 ( .A1(n690), .A2(n676), .ZN(n681) );
  INV_X1 U749 ( .A(n980), .ZN(n679) );
  NOR2_X1 U750 ( .A1(G1971), .A2(G303), .ZN(n677) );
  NOR2_X1 U751 ( .A1(n678), .A2(n677), .ZN(n971) );
  OR2_X1 U752 ( .A1(n679), .A2(n971), .ZN(n680) );
  AND2_X1 U753 ( .A1(n681), .A2(n680), .ZN(n683) );
  NOR2_X1 U754 ( .A1(n697), .A2(n684), .ZN(n685) );
  NOR2_X1 U755 ( .A1(KEYINPUT33), .A2(n685), .ZN(n686) );
  NOR2_X1 U756 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U757 ( .A1(n982), .A2(n688), .ZN(n702) );
  NAND2_X1 U758 ( .A1(n690), .A2(n689), .ZN(n693) );
  NOR2_X1 U759 ( .A1(G2090), .A2(G303), .ZN(n691) );
  NAND2_X1 U760 ( .A1(G8), .A2(n691), .ZN(n692) );
  NAND2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n694) );
  AND2_X1 U762 ( .A1(n694), .A2(n697), .ZN(n700) );
  NOR2_X1 U763 ( .A1(G1981), .A2(G305), .ZN(n695) );
  XOR2_X1 U764 ( .A(n695), .B(KEYINPUT24), .Z(n696) );
  NOR2_X1 U765 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U766 ( .A(n698), .B(KEYINPUT94), .ZN(n699) );
  NOR2_X1 U767 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U768 ( .A1(n702), .A2(n701), .ZN(n736) );
  NAND2_X1 U769 ( .A1(G119), .A2(n873), .ZN(n704) );
  NAND2_X1 U770 ( .A1(G107), .A2(n875), .ZN(n703) );
  NAND2_X1 U771 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U772 ( .A(KEYINPUT91), .B(n705), .ZN(n709) );
  NAND2_X1 U773 ( .A1(n848), .A2(G95), .ZN(n707) );
  NAND2_X1 U774 ( .A1(G131), .A2(n870), .ZN(n706) );
  AND2_X1 U775 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U776 ( .A1(n709), .A2(n708), .ZN(n886) );
  AND2_X1 U777 ( .A1(n886), .A2(G1991), .ZN(n720) );
  NAND2_X1 U778 ( .A1(G129), .A2(n873), .ZN(n711) );
  NAND2_X1 U779 ( .A1(G117), .A2(n875), .ZN(n710) );
  NAND2_X1 U780 ( .A1(n711), .A2(n710), .ZN(n714) );
  NAND2_X1 U781 ( .A1(n848), .A2(G105), .ZN(n712) );
  XOR2_X1 U782 ( .A(KEYINPUT38), .B(n712), .Z(n713) );
  NOR2_X1 U783 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U784 ( .A(n715), .B(KEYINPUT92), .ZN(n717) );
  NAND2_X1 U785 ( .A1(G141), .A2(n870), .ZN(n716) );
  NAND2_X1 U786 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U787 ( .A(KEYINPUT93), .B(n718), .Z(n881) );
  AND2_X1 U788 ( .A1(G1996), .A2(n881), .ZN(n719) );
  NOR2_X1 U789 ( .A1(n720), .A2(n719), .ZN(n914) );
  NOR2_X1 U790 ( .A1(n722), .A2(n721), .ZN(n750) );
  INV_X1 U791 ( .A(n750), .ZN(n723) );
  NOR2_X1 U792 ( .A1(n914), .A2(n723), .ZN(n742) );
  INV_X1 U793 ( .A(n742), .ZN(n734) );
  NAND2_X1 U794 ( .A1(n870), .A2(G140), .ZN(n724) );
  XNOR2_X1 U795 ( .A(n724), .B(KEYINPUT90), .ZN(n726) );
  NAND2_X1 U796 ( .A1(G104), .A2(n848), .ZN(n725) );
  NAND2_X1 U797 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U798 ( .A(KEYINPUT34), .B(n727), .ZN(n732) );
  NAND2_X1 U799 ( .A1(G128), .A2(n873), .ZN(n729) );
  NAND2_X1 U800 ( .A1(G116), .A2(n875), .ZN(n728) );
  NAND2_X1 U801 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U802 ( .A(KEYINPUT35), .B(n730), .Z(n731) );
  NOR2_X1 U803 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U804 ( .A(KEYINPUT36), .B(n733), .ZN(n887) );
  XNOR2_X1 U805 ( .A(G2067), .B(KEYINPUT37), .ZN(n748) );
  NOR2_X1 U806 ( .A1(n887), .A2(n748), .ZN(n917) );
  NAND2_X1 U807 ( .A1(n750), .A2(n917), .ZN(n746) );
  NAND2_X1 U808 ( .A1(n734), .A2(n746), .ZN(n735) );
  NOR2_X2 U809 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U810 ( .A(KEYINPUT106), .B(n737), .ZN(n739) );
  XNOR2_X1 U811 ( .A(G1986), .B(G290), .ZN(n979) );
  NAND2_X1 U812 ( .A1(n979), .A2(n750), .ZN(n738) );
  NAND2_X1 U813 ( .A1(n739), .A2(n738), .ZN(n753) );
  XOR2_X1 U814 ( .A(KEYINPUT107), .B(KEYINPUT39), .Z(n745) );
  NOR2_X1 U815 ( .A1(G1996), .A2(n881), .ZN(n928) );
  NOR2_X1 U816 ( .A1(G1986), .A2(G290), .ZN(n740) );
  NOR2_X1 U817 ( .A1(G1991), .A2(n886), .ZN(n919) );
  NOR2_X1 U818 ( .A1(n740), .A2(n919), .ZN(n741) );
  NOR2_X1 U819 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U820 ( .A1(n928), .A2(n743), .ZN(n744) );
  XNOR2_X1 U821 ( .A(n745), .B(n744), .ZN(n747) );
  NAND2_X1 U822 ( .A1(n747), .A2(n746), .ZN(n749) );
  NAND2_X1 U823 ( .A1(n887), .A2(n748), .ZN(n932) );
  NAND2_X1 U824 ( .A1(n749), .A2(n932), .ZN(n751) );
  NAND2_X1 U825 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U826 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U827 ( .A(n754), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U828 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U829 ( .A(G120), .ZN(G236) );
  INV_X1 U830 ( .A(G69), .ZN(G235) );
  INV_X1 U831 ( .A(G108), .ZN(G238) );
  NAND2_X1 U832 ( .A1(G7), .A2(G661), .ZN(n755) );
  XNOR2_X1 U833 ( .A(n755), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U834 ( .A(G223), .ZN(n823) );
  NAND2_X1 U835 ( .A1(n823), .A2(G567), .ZN(n756) );
  XOR2_X1 U836 ( .A(KEYINPUT11), .B(n756), .Z(G234) );
  NAND2_X1 U837 ( .A1(n967), .A2(G860), .ZN(G153) );
  XNOR2_X1 U838 ( .A(G171), .B(KEYINPUT71), .ZN(G301) );
  NAND2_X1 U839 ( .A1(G868), .A2(G301), .ZN(n758) );
  INV_X1 U840 ( .A(G868), .ZN(n765) );
  NAND2_X1 U841 ( .A1(n892), .A2(n765), .ZN(n757) );
  NAND2_X1 U842 ( .A1(n758), .A2(n757), .ZN(G284) );
  NAND2_X1 U843 ( .A1(n798), .A2(n765), .ZN(n759) );
  XNOR2_X1 U844 ( .A(n759), .B(KEYINPUT75), .ZN(n761) );
  NOR2_X1 U845 ( .A1(G286), .A2(n765), .ZN(n760) );
  NOR2_X1 U846 ( .A1(n761), .A2(n760), .ZN(G297) );
  INV_X1 U847 ( .A(G860), .ZN(n779) );
  NAND2_X1 U848 ( .A1(n779), .A2(G559), .ZN(n762) );
  NAND2_X1 U849 ( .A1(n762), .A2(n975), .ZN(n763) );
  XNOR2_X1 U850 ( .A(n763), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U851 ( .A1(G868), .A2(n975), .ZN(n764) );
  NOR2_X1 U852 ( .A1(G559), .A2(n764), .ZN(n767) );
  AND2_X1 U853 ( .A1(n765), .A2(n967), .ZN(n766) );
  NOR2_X1 U854 ( .A1(n767), .A2(n766), .ZN(G282) );
  NAND2_X1 U855 ( .A1(G123), .A2(n873), .ZN(n768) );
  XNOR2_X1 U856 ( .A(n768), .B(KEYINPUT18), .ZN(n770) );
  NAND2_X1 U857 ( .A1(n848), .A2(G99), .ZN(n769) );
  NAND2_X1 U858 ( .A1(n770), .A2(n769), .ZN(n774) );
  NAND2_X1 U859 ( .A1(G135), .A2(n870), .ZN(n772) );
  NAND2_X1 U860 ( .A1(G111), .A2(n875), .ZN(n771) );
  NAND2_X1 U861 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U862 ( .A1(n774), .A2(n773), .ZN(n918) );
  XNOR2_X1 U863 ( .A(n918), .B(G2096), .ZN(n775) );
  XNOR2_X1 U864 ( .A(n775), .B(KEYINPUT76), .ZN(n777) );
  INV_X1 U865 ( .A(G2100), .ZN(n776) );
  NAND2_X1 U866 ( .A1(n777), .A2(n776), .ZN(G156) );
  NAND2_X1 U867 ( .A1(n975), .A2(G559), .ZN(n778) );
  XNOR2_X1 U868 ( .A(n778), .B(n967), .ZN(n801) );
  NAND2_X1 U869 ( .A1(n779), .A2(n801), .ZN(n791) );
  NAND2_X1 U870 ( .A1(G93), .A2(n780), .ZN(n783) );
  NAND2_X1 U871 ( .A1(G80), .A2(n781), .ZN(n782) );
  NAND2_X1 U872 ( .A1(n783), .A2(n782), .ZN(n790) );
  NAND2_X1 U873 ( .A1(G67), .A2(n784), .ZN(n785) );
  XOR2_X1 U874 ( .A(KEYINPUT77), .B(n785), .Z(n788) );
  NAND2_X1 U875 ( .A1(n786), .A2(G55), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U877 ( .A1(n790), .A2(n789), .ZN(n804) );
  XOR2_X1 U878 ( .A(n791), .B(n804), .Z(G145) );
  XNOR2_X1 U879 ( .A(KEYINPUT80), .B(KEYINPUT81), .ZN(n793) );
  XNOR2_X1 U880 ( .A(G288), .B(G166), .ZN(n792) );
  XNOR2_X1 U881 ( .A(n793), .B(n792), .ZN(n794) );
  XNOR2_X1 U882 ( .A(KEYINPUT19), .B(n794), .ZN(n796) );
  XNOR2_X1 U883 ( .A(G305), .B(KEYINPUT82), .ZN(n795) );
  XNOR2_X1 U884 ( .A(n796), .B(n795), .ZN(n797) );
  XNOR2_X1 U885 ( .A(n804), .B(n797), .ZN(n800) );
  XNOR2_X1 U886 ( .A(G290), .B(n798), .ZN(n799) );
  XNOR2_X1 U887 ( .A(n800), .B(n799), .ZN(n891) );
  XNOR2_X1 U888 ( .A(n891), .B(n801), .ZN(n802) );
  NAND2_X1 U889 ( .A1(n802), .A2(G868), .ZN(n803) );
  XOR2_X1 U890 ( .A(KEYINPUT83), .B(n803), .Z(n806) );
  OR2_X1 U891 ( .A1(n804), .A2(G868), .ZN(n805) );
  NAND2_X1 U892 ( .A1(n806), .A2(n805), .ZN(G295) );
  NAND2_X1 U893 ( .A1(G2084), .A2(G2078), .ZN(n807) );
  XOR2_X1 U894 ( .A(KEYINPUT20), .B(n807), .Z(n808) );
  NAND2_X1 U895 ( .A1(n808), .A2(G2090), .ZN(n809) );
  XNOR2_X1 U896 ( .A(n809), .B(KEYINPUT21), .ZN(n810) );
  XNOR2_X1 U897 ( .A(KEYINPUT84), .B(n810), .ZN(n811) );
  NAND2_X1 U898 ( .A1(G2072), .A2(n811), .ZN(G158) );
  XNOR2_X1 U899 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U900 ( .A1(G235), .A2(G236), .ZN(n812) );
  XOR2_X1 U901 ( .A(KEYINPUT86), .B(n812), .Z(n813) );
  NOR2_X1 U902 ( .A1(G238), .A2(n813), .ZN(n814) );
  NAND2_X1 U903 ( .A1(G57), .A2(n814), .ZN(n827) );
  NAND2_X1 U904 ( .A1(G567), .A2(n827), .ZN(n820) );
  XOR2_X1 U905 ( .A(KEYINPUT22), .B(KEYINPUT85), .Z(n816) );
  NAND2_X1 U906 ( .A1(G132), .A2(G82), .ZN(n815) );
  XNOR2_X1 U907 ( .A(n816), .B(n815), .ZN(n817) );
  NOR2_X1 U908 ( .A1(n817), .A2(G218), .ZN(n818) );
  NAND2_X1 U909 ( .A1(G96), .A2(n818), .ZN(n828) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n828), .ZN(n819) );
  NAND2_X1 U911 ( .A1(n820), .A2(n819), .ZN(n829) );
  NAND2_X1 U912 ( .A1(G483), .A2(G661), .ZN(n821) );
  NOR2_X1 U913 ( .A1(n829), .A2(n821), .ZN(n822) );
  XOR2_X1 U914 ( .A(KEYINPUT87), .B(n822), .Z(n826) );
  NAND2_X1 U915 ( .A1(n826), .A2(G36), .ZN(G176) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n823), .ZN(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n824) );
  NAND2_X1 U918 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n826), .A2(n825), .ZN(G188) );
  INV_X1 U922 ( .A(G132), .ZN(G219) );
  INV_X1 U923 ( .A(G96), .ZN(G221) );
  INV_X1 U924 ( .A(G82), .ZN(G220) );
  NOR2_X1 U925 ( .A1(n828), .A2(n827), .ZN(G325) );
  INV_X1 U926 ( .A(G325), .ZN(G261) );
  XOR2_X1 U927 ( .A(KEYINPUT108), .B(n829), .Z(G319) );
  XOR2_X1 U928 ( .A(KEYINPUT42), .B(G2090), .Z(n831) );
  XNOR2_X1 U929 ( .A(G2084), .B(G2072), .ZN(n830) );
  XNOR2_X1 U930 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U931 ( .A(n832), .B(G2100), .Z(n834) );
  XNOR2_X1 U932 ( .A(G2067), .B(G2078), .ZN(n833) );
  XNOR2_X1 U933 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U934 ( .A(G2096), .B(KEYINPUT43), .Z(n836) );
  XNOR2_X1 U935 ( .A(KEYINPUT109), .B(G2678), .ZN(n835) );
  XNOR2_X1 U936 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U937 ( .A(n838), .B(n837), .Z(G227) );
  XOR2_X1 U938 ( .A(G1966), .B(G1971), .Z(n840) );
  XNOR2_X1 U939 ( .A(G1981), .B(G1976), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U941 ( .A(n841), .B(KEYINPUT41), .Z(n843) );
  XNOR2_X1 U942 ( .A(G1996), .B(G1991), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U944 ( .A(G2474), .B(G1956), .Z(n845) );
  XNOR2_X1 U945 ( .A(G1986), .B(G1961), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(G229) );
  NAND2_X1 U948 ( .A1(n875), .A2(G112), .ZN(n855) );
  NAND2_X1 U949 ( .A1(G100), .A2(n848), .ZN(n850) );
  NAND2_X1 U950 ( .A1(G136), .A2(n870), .ZN(n849) );
  NAND2_X1 U951 ( .A1(n850), .A2(n849), .ZN(n853) );
  NAND2_X1 U952 ( .A1(n873), .A2(G124), .ZN(n851) );
  XOR2_X1 U953 ( .A(KEYINPUT44), .B(n851), .Z(n852) );
  NOR2_X1 U954 ( .A1(n853), .A2(n852), .ZN(n854) );
  NAND2_X1 U955 ( .A1(n855), .A2(n854), .ZN(n856) );
  XOR2_X1 U956 ( .A(KEYINPUT110), .B(n856), .Z(G162) );
  NAND2_X1 U957 ( .A1(G130), .A2(n873), .ZN(n858) );
  NAND2_X1 U958 ( .A1(G118), .A2(n875), .ZN(n857) );
  NAND2_X1 U959 ( .A1(n858), .A2(n857), .ZN(n864) );
  NAND2_X1 U960 ( .A1(G106), .A2(n848), .ZN(n860) );
  NAND2_X1 U961 ( .A1(G142), .A2(n870), .ZN(n859) );
  NAND2_X1 U962 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U963 ( .A(KEYINPUT111), .B(n861), .ZN(n862) );
  XNOR2_X1 U964 ( .A(KEYINPUT45), .B(n862), .ZN(n863) );
  NOR2_X1 U965 ( .A1(n864), .A2(n863), .ZN(n868) );
  XOR2_X1 U966 ( .A(KEYINPUT48), .B(KEYINPUT113), .Z(n866) );
  XNOR2_X1 U967 ( .A(G164), .B(KEYINPUT46), .ZN(n865) );
  XNOR2_X1 U968 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U969 ( .A(n868), .B(n867), .Z(n869) );
  XNOR2_X1 U970 ( .A(G162), .B(n869), .ZN(n885) );
  NAND2_X1 U971 ( .A1(G103), .A2(n848), .ZN(n872) );
  NAND2_X1 U972 ( .A1(G139), .A2(n870), .ZN(n871) );
  NAND2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n880) );
  NAND2_X1 U974 ( .A1(n873), .A2(G127), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n874), .B(KEYINPUT112), .ZN(n877) );
  NAND2_X1 U976 ( .A1(G115), .A2(n875), .ZN(n876) );
  NAND2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U978 ( .A(KEYINPUT47), .B(n878), .Z(n879) );
  NOR2_X1 U979 ( .A1(n880), .A2(n879), .ZN(n923) );
  XOR2_X1 U980 ( .A(n918), .B(n923), .Z(n883) );
  XOR2_X1 U981 ( .A(G160), .B(n881), .Z(n882) );
  XNOR2_X1 U982 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U983 ( .A(n885), .B(n884), .ZN(n889) );
  XOR2_X1 U984 ( .A(n887), .B(n886), .Z(n888) );
  XNOR2_X1 U985 ( .A(n889), .B(n888), .ZN(n890) );
  NOR2_X1 U986 ( .A1(G37), .A2(n890), .ZN(G395) );
  XOR2_X1 U987 ( .A(KEYINPUT114), .B(n891), .Z(n894) );
  XNOR2_X1 U988 ( .A(n892), .B(n967), .ZN(n893) );
  XNOR2_X1 U989 ( .A(n894), .B(n893), .ZN(n896) );
  XOR2_X1 U990 ( .A(G286), .B(G171), .Z(n895) );
  XNOR2_X1 U991 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U992 ( .A1(G37), .A2(n897), .ZN(G397) );
  XOR2_X1 U993 ( .A(G2451), .B(G2430), .Z(n899) );
  XNOR2_X1 U994 ( .A(G2438), .B(G2443), .ZN(n898) );
  XNOR2_X1 U995 ( .A(n899), .B(n898), .ZN(n905) );
  XOR2_X1 U996 ( .A(G2435), .B(G2454), .Z(n901) );
  XNOR2_X1 U997 ( .A(G1341), .B(G1348), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n903) );
  XOR2_X1 U999 ( .A(G2446), .B(G2427), .Z(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1001 ( .A(n905), .B(n904), .Z(n906) );
  NAND2_X1 U1002 ( .A1(G14), .A2(n906), .ZN(n913) );
  NAND2_X1 U1003 ( .A1(n913), .A2(G319), .ZN(n910) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n907) );
  XOR2_X1 U1005 ( .A(KEYINPUT115), .B(n907), .Z(n908) );
  XNOR2_X1 U1006 ( .A(n908), .B(KEYINPUT49), .ZN(n909) );
  NOR2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(n912) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(G57), .ZN(G237) );
  INV_X1 U1012 ( .A(n913), .ZN(G401) );
  XNOR2_X1 U1013 ( .A(KEYINPUT52), .B(KEYINPUT117), .ZN(n937) );
  XNOR2_X1 U1014 ( .A(G160), .B(G2084), .ZN(n915) );
  NAND2_X1 U1015 ( .A1(n915), .A2(n914), .ZN(n916) );
  NOR2_X1 U1016 ( .A1(n917), .A2(n916), .ZN(n921) );
  NOR2_X1 U1017 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1019 ( .A(KEYINPUT116), .B(n922), .ZN(n935) );
  XOR2_X1 U1020 ( .A(G2072), .B(n923), .Z(n925) );
  XOR2_X1 U1021 ( .A(G164), .B(G2078), .Z(n924) );
  NOR2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1023 ( .A(KEYINPUT50), .B(n926), .Z(n931) );
  XOR2_X1 U1024 ( .A(G2090), .B(G162), .Z(n927) );
  NOR2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(KEYINPUT51), .B(n929), .ZN(n930) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n933) );
  NAND2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1030 ( .A(n937), .B(n936), .ZN(n938) );
  NOR2_X1 U1031 ( .A1(KEYINPUT55), .A2(n938), .ZN(n939) );
  XOR2_X1 U1032 ( .A(KEYINPUT118), .B(n939), .Z(n940) );
  NAND2_X1 U1033 ( .A1(n940), .A2(G29), .ZN(n941) );
  XOR2_X1 U1034 ( .A(KEYINPUT119), .B(n941), .Z(n1021) );
  XOR2_X1 U1035 ( .A(KEYINPUT55), .B(KEYINPUT124), .Z(n963) );
  XNOR2_X1 U1036 ( .A(G2090), .B(G35), .ZN(n942) );
  XNOR2_X1 U1037 ( .A(n942), .B(KEYINPUT120), .ZN(n958) );
  XNOR2_X1 U1038 ( .A(KEYINPUT121), .B(G2067), .ZN(n943) );
  XNOR2_X1 U1039 ( .A(n943), .B(G26), .ZN(n951) );
  XNOR2_X1 U1040 ( .A(G1996), .B(G32), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(G1991), .B(G25), .ZN(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1043 ( .A1(G28), .A2(n946), .ZN(n949) );
  XNOR2_X1 U1044 ( .A(KEYINPUT122), .B(G2072), .ZN(n947) );
  XNOR2_X1 U1045 ( .A(G33), .B(n947), .ZN(n948) );
  NOR2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(G27), .B(n952), .ZN(n953) );
  XNOR2_X1 U1049 ( .A(KEYINPUT123), .B(n953), .ZN(n954) );
  NOR2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(n956), .B(KEYINPUT53), .ZN(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n961) );
  XOR2_X1 U1053 ( .A(G2084), .B(G34), .Z(n959) );
  XNOR2_X1 U1054 ( .A(KEYINPUT54), .B(n959), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(n963), .B(n962), .ZN(n965) );
  INV_X1 U1057 ( .A(G29), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1059 ( .A1(G11), .A2(n966), .ZN(n1019) );
  XNOR2_X1 U1060 ( .A(G16), .B(KEYINPUT56), .ZN(n990) );
  XOR2_X1 U1061 ( .A(n967), .B(G1341), .Z(n969) );
  XNOR2_X1 U1062 ( .A(G299), .B(G1956), .ZN(n968) );
  NOR2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n974) );
  XNOR2_X1 U1065 ( .A(G1961), .B(G171), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(KEYINPUT125), .B(n972), .ZN(n973) );
  NOR2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n988) );
  XNOR2_X1 U1068 ( .A(n975), .B(G1348), .ZN(n977) );
  NAND2_X1 U1069 ( .A1(G303), .A2(G1971), .ZN(n976) );
  NAND2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n981) );
  NAND2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n986) );
  XNOR2_X1 U1073 ( .A(G1966), .B(G168), .ZN(n983) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1075 ( .A(KEYINPUT57), .B(n984), .Z(n985) );
  NOR2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n1017) );
  INV_X1 U1079 ( .A(G16), .ZN(n1015) );
  XNOR2_X1 U1080 ( .A(KEYINPUT59), .B(G1348), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(n991), .B(G4), .ZN(n996) );
  XOR2_X1 U1082 ( .A(G1981), .B(KEYINPUT127), .Z(n992) );
  XNOR2_X1 U1083 ( .A(G6), .B(n992), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(G19), .B(G1341), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n1000) );
  XOR2_X1 U1087 ( .A(KEYINPUT126), .B(n997), .Z(n998) );
  XNOR2_X1 U1088 ( .A(G20), .B(n998), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(KEYINPUT60), .B(n1001), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(G1966), .B(G21), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(G1961), .B(G5), .ZN(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1012) );
  XNOR2_X1 U1095 ( .A(G1976), .B(G23), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(G1971), .B(G22), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  XOR2_X1 U1098 ( .A(G1986), .B(G24), .Z(n1008) );
  NAND2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(KEYINPUT58), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(KEYINPUT61), .B(n1013), .ZN(n1014) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1022), .Z(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

