//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n927, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960;
  INV_X1    g000(.A(G226gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT24), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT64), .A4(new_n210), .ZN(new_n214));
  AND2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT67), .ZN(new_n216));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT66), .B(KEYINPUT23), .ZN(new_n218));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(G176gat), .ZN(new_n222));
  OR2_X1    g021(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n216), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n221), .A2(KEYINPUT66), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT23), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n229), .A3(new_n219), .ZN(new_n230));
  INV_X1    g029(.A(new_n217), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n232), .A2(KEYINPUT67), .A3(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n215), .A2(new_n226), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT25), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(KEYINPUT68), .B(G183gat), .Z(new_n238));
  OAI211_X1 g037(.A(new_n208), .B(new_n210), .C1(new_n238), .C2(G190gat), .ZN(new_n239));
  INV_X1    g038(.A(G169gat), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n236), .B1(new_n222), .B2(new_n240), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n239), .A2(new_n232), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n237), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT28), .ZN(new_n245));
  NOR2_X1   g044(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n246), .B1(new_n238), .B2(KEYINPUT27), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n245), .B1(new_n247), .B2(G190gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT27), .B(G183gat), .ZN(new_n249));
  INV_X1    g048(.A(G190gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(KEYINPUT28), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n253));
  OR3_X1    g052(.A1(new_n253), .A2(new_n217), .A3(KEYINPUT69), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT69), .B1(new_n253), .B2(new_n217), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT26), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n217), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n254), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n252), .A2(new_n206), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n205), .B1(new_n244), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT29), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n242), .B1(new_n235), .B2(new_n236), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n258), .A2(new_n206), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n263), .B1(new_n248), .B2(new_n251), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n261), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n260), .B1(new_n205), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G197gat), .B(G204gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT22), .ZN(new_n268));
  INV_X1    g067(.A(G211gat), .ZN(new_n269));
  INV_X1    g068(.A(G218gat), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G211gat), .B(G218gat), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n272), .B(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT76), .B1(new_n266), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n265), .A2(new_n205), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT77), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n204), .B1(new_n262), .B2(new_n264), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT78), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI211_X1 g081(.A(KEYINPUT78), .B(new_n204), .C1(new_n262), .C2(new_n264), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n265), .A2(KEYINPUT77), .A3(new_n205), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n279), .A2(new_n284), .A3(new_n275), .A4(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT37), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n277), .A2(new_n280), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT76), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n272), .B(new_n273), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND4_X1  g090(.A1(new_n276), .A2(new_n286), .A3(new_n287), .A4(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT87), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n289), .B1(new_n288), .B2(new_n290), .ZN(new_n295));
  AOI211_X1 g094(.A(KEYINPUT76), .B(new_n275), .C1(new_n277), .C2(new_n280), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n297), .A2(KEYINPUT87), .A3(new_n287), .A4(new_n286), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G8gat), .B(G36gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(G64gat), .B(G92gat), .ZN(new_n301));
  XOR2_X1   g100(.A(new_n300), .B(new_n301), .Z(new_n302));
  NAND3_X1  g101(.A1(new_n276), .A2(new_n286), .A3(new_n291), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n302), .B1(new_n303), .B2(KEYINPUT37), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n299), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT38), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n279), .A2(new_n284), .A3(new_n290), .A4(new_n285), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n287), .B1(new_n288), .B2(new_n275), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n302), .A2(KEYINPUT38), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n299), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT88), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT5), .ZN(new_n316));
  XNOR2_X1  g115(.A(G141gat), .B(G148gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n317), .B1(KEYINPUT2), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G155gat), .ZN(new_n320));
  INV_X1    g119(.A(G162gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(new_n318), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n318), .B(new_n322), .C1(new_n317), .C2(KEYINPUT2), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G127gat), .B(G134gat), .ZN(new_n327));
  INV_X1    g126(.A(G113gat), .ZN(new_n328));
  INV_X1    g127(.A(G120gat), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT1), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  XOR2_X1   g129(.A(KEYINPUT70), .B(G113gat), .Z(new_n331));
  OAI211_X1 g130(.A(new_n327), .B(new_n330), .C1(new_n331), .C2(new_n329), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n330), .B1(new_n328), .B2(new_n329), .ZN(new_n333));
  INV_X1    g132(.A(new_n327), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n326), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT80), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT80), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(new_n326), .B2(new_n336), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n326), .A2(new_n336), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n338), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G225gat), .A2(G233gat), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n316), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT79), .B1(new_n326), .B2(KEYINPUT3), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT79), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT3), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n324), .A2(new_n347), .A3(new_n348), .A4(new_n325), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n336), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n351), .B1(KEYINPUT3), .B2(new_n326), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT4), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n354), .A3(new_n340), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n344), .B1(new_n337), .B2(KEYINPUT4), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n353), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n345), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n337), .A2(KEYINPUT4), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n359), .B1(new_n350), .B2(new_n352), .ZN(new_n360));
  INV_X1    g159(.A(new_n340), .ZN(new_n361));
  NOR3_X1   g160(.A1(new_n326), .A2(new_n336), .A3(new_n339), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT4), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n360), .A2(new_n363), .A3(new_n316), .A4(new_n343), .ZN(new_n364));
  XOR2_X1   g163(.A(G1gat), .B(G29gat), .Z(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G57gat), .B(G85gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n358), .A2(new_n364), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT6), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n358), .A2(new_n364), .ZN(new_n373));
  INV_X1    g172(.A(new_n369), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n372), .B(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n297), .A2(new_n286), .A3(new_n302), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n299), .A2(KEYINPUT88), .A3(new_n312), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n306), .A2(new_n315), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n302), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n303), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n383), .A2(new_n377), .A3(KEYINPUT30), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n343), .B1(new_n360), .B2(new_n363), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT39), .B1(new_n342), .B2(new_n344), .ZN(new_n386));
  OR2_X1    g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT39), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n374), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n387), .A2(KEYINPUT40), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n375), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT40), .B1(new_n387), .B2(new_n389), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OR3_X1    g192(.A1(new_n303), .A2(KEYINPUT30), .A3(new_n382), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n384), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n350), .A2(new_n261), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n290), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n290), .A2(KEYINPUT29), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n348), .B1(new_n398), .B2(KEYINPUT85), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n275), .A2(KEYINPUT85), .A3(new_n261), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n326), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n397), .A2(G228gat), .A3(G233gat), .A4(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(G228gat), .A2(G233gat), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n275), .B1(new_n350), .B2(new_n261), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n275), .A2(new_n261), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT3), .B1(new_n405), .B2(KEYINPUT84), .ZN(new_n406));
  OR3_X1    g205(.A1(new_n290), .A2(KEYINPUT84), .A3(KEYINPUT29), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n406), .A2(new_n407), .B1(new_n325), .B2(new_n324), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n403), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n402), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(G22gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT86), .B(G22gat), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n402), .A2(new_n412), .A3(new_n409), .ZN(new_n413));
  XNOR2_X1  g212(.A(G78gat), .B(G106gat), .ZN(new_n414));
  INV_X1    g213(.A(G50gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n411), .A2(new_n413), .A3(new_n418), .ZN(new_n419));
  XOR2_X1   g218(.A(new_n418), .B(KEYINPUT83), .Z(new_n420));
  INV_X1    g219(.A(new_n412), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n410), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n420), .B1(new_n422), .B2(new_n413), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n395), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n381), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n376), .B1(new_n384), .B2(new_n394), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n429), .A2(new_n425), .ZN(new_n430));
  XNOR2_X1  g229(.A(G15gat), .B(G43gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(G71gat), .B(G99gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n213), .A2(new_n214), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n223), .A2(new_n224), .ZN(new_n435));
  AOI22_X1  g234(.A1(new_n435), .A2(new_n222), .B1(new_n230), .B2(new_n231), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n434), .B1(KEYINPUT67), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT25), .B1(new_n437), .B2(new_n226), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n259), .B(new_n336), .C1(new_n438), .C2(new_n242), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n351), .B1(new_n262), .B2(new_n264), .ZN(new_n440));
  INV_X1    g239(.A(G227gat), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n441), .A2(new_n203), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n439), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT71), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n439), .A2(new_n440), .A3(KEYINPUT71), .A4(new_n442), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT32), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT33), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n433), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n433), .ZN(new_n451));
  OR2_X1    g250(.A1(new_n451), .A2(KEYINPUT72), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT33), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n453), .B1(new_n451), .B2(KEYINPUT72), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n448), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n456), .B1(new_n445), .B2(new_n446), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT75), .B1(new_n450), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n447), .A2(new_n455), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT75), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n445), .A2(new_n446), .B1(new_n448), .B2(KEYINPUT33), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n459), .B(new_n460), .C1(new_n461), .C2(new_n433), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n442), .B1(new_n439), .B2(new_n440), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n464), .A2(KEYINPUT34), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT74), .ZN(new_n466));
  XNOR2_X1  g265(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n466), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n467), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n463), .A2(KEYINPUT74), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n465), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n458), .A2(new_n462), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n450), .A2(new_n457), .ZN(new_n475));
  OAI22_X1  g274(.A1(new_n468), .A2(new_n471), .B1(KEYINPUT34), .B2(new_n464), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(new_n460), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n474), .A2(KEYINPUT36), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT36), .B1(new_n474), .B2(new_n477), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n430), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n424), .B1(new_n474), .B2(new_n477), .ZN(new_n482));
  NAND2_X1  g281(.A1(KEYINPUT89), .A2(KEYINPUT35), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(new_n429), .A3(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(KEYINPUT89), .A2(KEYINPUT35), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n482), .A2(new_n429), .A3(new_n485), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n428), .A2(new_n481), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G113gat), .B(G141gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(G197gat), .ZN(new_n491));
  XOR2_X1   g290(.A(KEYINPUT11), .B(G169gat), .Z(new_n492));
  XNOR2_X1  g291(.A(new_n491), .B(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(KEYINPUT12), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(G229gat), .A2(G233gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(G15gat), .B(G22gat), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n497), .A2(G1gat), .ZN(new_n498));
  INV_X1    g297(.A(G1gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT16), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n498), .B1(new_n500), .B2(new_n497), .ZN(new_n501));
  INV_X1    g300(.A(G8gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT17), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n415), .A2(G43gat), .ZN(new_n505));
  INV_X1    g304(.A(G43gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(G50gat), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(new_n507), .A3(KEYINPUT15), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(G29gat), .A2(G36gat), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n511));
  NOR3_X1   g310(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n511), .B1(new_n512), .B2(KEYINPUT90), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT14), .ZN(new_n514));
  INV_X1    g313(.A(G29gat), .ZN(new_n515));
  INV_X1    g314(.A(G36gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT90), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n510), .B1(new_n513), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n517), .A2(new_n511), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n521), .A2(new_n508), .A3(new_n510), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT15), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n506), .A2(KEYINPUT91), .A3(G50gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n505), .A2(new_n507), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n523), .B(new_n524), .C1(new_n525), .C2(KEYINPUT91), .ZN(new_n526));
  AOI22_X1  g325(.A1(new_n509), .A2(new_n520), .B1(new_n522), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT92), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n504), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n520), .A2(new_n509), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n522), .A2(new_n526), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n532), .A2(KEYINPUT92), .A3(KEYINPUT17), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n503), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT93), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n501), .B(G8gat), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n535), .B1(new_n536), .B2(new_n527), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  AOI211_X1 g337(.A(new_n535), .B(new_n503), .C1(new_n533), .C2(new_n529), .ZN(new_n539));
  OAI211_X1 g338(.A(KEYINPUT18), .B(new_n496), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n503), .B(new_n527), .ZN(new_n541));
  XOR2_X1   g340(.A(new_n496), .B(KEYINPUT13), .Z(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n534), .A2(KEYINPUT93), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n546), .B1(new_n534), .B2(new_n537), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT18), .B1(new_n547), .B2(new_n496), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n495), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n496), .B1(new_n538), .B2(new_n539), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT18), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n552), .A2(new_n494), .A3(new_n540), .A4(new_n544), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n549), .A2(KEYINPUT94), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT94), .B1(new_n549), .B2(new_n553), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G134gat), .B(G162gat), .Z(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n560));
  INV_X1    g359(.A(G85gat), .ZN(new_n561));
  INV_X1    g360(.A(G92gat), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G99gat), .A2(G106gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(new_n562), .ZN(new_n566));
  NAND4_X1  g365(.A1(KEYINPUT98), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n563), .A2(new_n565), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G99gat), .B(G106gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  AOI22_X1  g370(.A1(KEYINPUT8), .A2(new_n564), .B1(new_n561), .B2(new_n562), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n572), .A2(new_n569), .A3(new_n563), .A4(new_n567), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  AND2_X1   g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n532), .A2(new_n575), .B1(KEYINPUT41), .B2(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n529), .A2(new_n533), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n250), .B(new_n577), .C1(new_n578), .C2(new_n575), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n575), .B1(new_n529), .B2(new_n533), .ZN(new_n580));
  INV_X1    g379(.A(new_n577), .ZN(new_n581));
  OAI21_X1  g380(.A(G190gat), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT97), .B1(new_n583), .B2(new_n270), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n576), .A2(KEYINPUT41), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n579), .A2(G218gat), .A3(new_n582), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n586), .B1(new_n584), .B2(new_n587), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n559), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n584), .A2(new_n587), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n585), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n592), .A2(new_n558), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT9), .ZN(new_n596));
  INV_X1    g395(.A(G71gat), .ZN(new_n597));
  INV_X1    g396(.A(G78gat), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT95), .ZN(new_n600));
  XOR2_X1   g399(.A(G57gat), .B(G64gat), .Z(new_n601));
  XNOR2_X1  g400(.A(G71gat), .B(G78gat), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT95), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n603), .B(new_n596), .C1(new_n597), .C2(new_n598), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n600), .A2(new_n601), .A3(new_n602), .A4(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n602), .ZN(new_n606));
  XNOR2_X1  g405(.A(G57gat), .B(G64gat), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n606), .B1(new_n596), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n610), .A2(KEYINPUT21), .ZN(new_n611));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G127gat), .B(G155gat), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n614), .B(KEYINPUT20), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n613), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G183gat), .B(G211gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n503), .B1(KEYINPUT21), .B2(new_n610), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n618), .B(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n595), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G230gat), .A2(G233gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n574), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT10), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n605), .A2(new_n571), .A3(new_n608), .A4(new_n573), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n628), .A2(KEYINPUT99), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT99), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n625), .A2(new_n630), .A3(new_n626), .A4(new_n627), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n610), .A2(new_n575), .A3(KEYINPUT10), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n624), .B1(new_n629), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n625), .A2(new_n627), .ZN(new_n635));
  INV_X1    g434(.A(new_n624), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G120gat), .B(G148gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(G176gat), .B(G204gat), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n639), .B(new_n640), .Z(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n634), .A2(new_n637), .A3(new_n641), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n623), .A2(new_n646), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n489), .A2(new_n557), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n376), .B(KEYINPUT100), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT101), .B(G1gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(G1324gat));
  NAND2_X1  g451(.A1(new_n384), .A2(new_n394), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  XOR2_X1   g453(.A(KEYINPUT16), .B(G8gat), .Z(new_n655));
  NAND3_X1  g454(.A1(new_n648), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n648), .ZN(new_n657));
  OAI21_X1  g456(.A(G8gat), .B1(new_n657), .B2(new_n653), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n656), .ZN(new_n659));
  MUX2_X1   g458(.A(new_n656), .B(new_n659), .S(KEYINPUT42), .Z(G1325gat));
  NOR2_X1   g459(.A1(new_n479), .A2(new_n480), .ZN(new_n661));
  OAI21_X1  g460(.A(G15gat), .B1(new_n657), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n474), .A2(new_n477), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n664), .A2(G15gat), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n662), .B1(new_n657), .B2(new_n665), .ZN(G1326gat));
  NAND2_X1  g465(.A1(new_n648), .A2(new_n424), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT43), .B(G22gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670));
  INV_X1    g469(.A(new_n595), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n670), .B1(new_n489), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(KEYINPUT88), .B1(new_n299), .B2(new_n312), .ZN(new_n673));
  AOI211_X1 g472(.A(new_n314), .B(new_n311), .C1(new_n294), .C2(new_n298), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n378), .B1(new_n305), .B2(KEYINPUT38), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n426), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT36), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n678), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n679), .B(new_n478), .C1(new_n425), .C2(new_n429), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  AND3_X1   g480(.A1(new_n482), .A2(new_n429), .A3(new_n485), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n486), .B2(new_n484), .ZN(new_n683));
  OAI211_X1 g482(.A(KEYINPUT44), .B(new_n595), .C1(new_n681), .C2(new_n683), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n672), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n622), .A2(new_n646), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n549), .A2(new_n553), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n649), .ZN(new_n691));
  OAI21_X1  g490(.A(G29gat), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n489), .A2(new_n557), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n671), .A2(new_n686), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n649), .A2(new_n515), .ZN(new_n696));
  OR3_X1    g495(.A1(new_n695), .A2(KEYINPUT102), .A3(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n698));
  OAI21_X1  g497(.A(KEYINPUT102), .B1(new_n695), .B2(new_n696), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n698), .B1(new_n697), .B2(new_n699), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n692), .B1(new_n700), .B2(new_n701), .ZN(G1328gat));
  NOR3_X1   g501(.A1(new_n695), .A2(G36gat), .A3(new_n653), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT46), .ZN(new_n704));
  OAI21_X1  g503(.A(G36gat), .B1(new_n690), .B2(new_n653), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(G1329gat));
  OAI21_X1  g505(.A(G43gat), .B1(new_n690), .B2(new_n661), .ZN(new_n707));
  NAND2_X1  g506(.A1(KEYINPUT104), .A2(KEYINPUT47), .ZN(new_n708));
  NOR2_X1   g507(.A1(KEYINPUT104), .A2(KEYINPUT47), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n664), .A2(G43gat), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n693), .A2(new_n694), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT103), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT103), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n693), .A2(new_n713), .A3(new_n694), .A4(new_n710), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n709), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n707), .A2(new_n708), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n708), .B1(new_n707), .B2(new_n715), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(G1330gat));
  OAI21_X1  g517(.A(new_n415), .B1(new_n695), .B2(new_n425), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n424), .A2(G50gat), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n719), .B1(new_n690), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g521(.A1(new_n487), .A2(new_n488), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(new_n677), .B2(new_n680), .ZN(new_n724));
  AND4_X1   g523(.A1(new_n688), .A2(new_n724), .A3(new_n623), .A4(new_n645), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n649), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT105), .B(G57gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1332gat));
  AOI21_X1  g527(.A(new_n653), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT106), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n725), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n731), .B(new_n732), .Z(G1333gat));
  NAND3_X1  g532(.A1(new_n725), .A2(new_n597), .A3(new_n663), .ZN(new_n734));
  INV_X1    g533(.A(new_n661), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n725), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n736), .B2(new_n597), .ZN(new_n737));
  XNOR2_X1  g536(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1334gat));
  NAND2_X1  g538(.A1(new_n725), .A2(new_n424), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G78gat), .ZN(G1335gat));
  INV_X1    g540(.A(new_n622), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n687), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n595), .B(new_n743), .C1(new_n681), .C2(new_n683), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n724), .A2(KEYINPUT51), .A3(new_n595), .A4(new_n743), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n746), .A2(KEYINPUT108), .A3(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n744), .A2(new_n749), .A3(new_n745), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n691), .A2(G85gat), .A3(new_n646), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n748), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n742), .A2(new_n687), .A3(new_n646), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n672), .A2(new_n649), .A3(new_n684), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G85gat), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT109), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1336gat));
  NOR3_X1   g557(.A1(new_n653), .A2(G92gat), .A3(new_n646), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n748), .A2(new_n750), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT110), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n672), .A2(new_n654), .A3(new_n684), .A4(new_n753), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G92gat), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n761), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n760), .A2(KEYINPUT110), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n744), .A2(new_n745), .ZN(new_n767));
  INV_X1    g566(.A(new_n747), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n759), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n769), .A2(new_n764), .ZN(new_n770));
  OAI22_X1  g569(.A1(new_n765), .A2(new_n766), .B1(new_n762), .B2(new_n770), .ZN(G1337gat));
  NAND3_X1  g570(.A1(new_n685), .A2(new_n735), .A3(new_n753), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G99gat), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n664), .A2(G99gat), .A3(new_n646), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n748), .A2(new_n750), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(G1338gat));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n425), .A2(G106gat), .A3(new_n646), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n748), .A2(new_n750), .A3(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n672), .A2(new_n424), .A3(new_n684), .A4(new_n753), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT53), .B1(new_n780), .B2(G106gat), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n778), .B1(new_n767), .B2(new_n768), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n780), .A2(G106gat), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n777), .B1(new_n782), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n779), .A2(new_n781), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n784), .A2(new_n785), .ZN(new_n789));
  OAI211_X1 g588(.A(KEYINPUT111), .B(new_n788), .C1(new_n789), .C2(new_n783), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(G1339gat));
  NAND2_X1  g590(.A1(new_n628), .A2(KEYINPUT99), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n792), .A2(new_n636), .A3(new_n631), .A4(new_n632), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n634), .A2(KEYINPUT54), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT54), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n795), .B(new_n624), .C1(new_n629), .C2(new_n633), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n794), .A2(KEYINPUT55), .A3(new_n642), .A4(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT112), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n796), .A2(new_n642), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n800), .A2(KEYINPUT112), .A3(KEYINPUT55), .A4(new_n794), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n799), .A2(new_n644), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n634), .A2(KEYINPUT54), .A3(new_n793), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n796), .A2(new_n642), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT113), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n794), .A2(new_n642), .A3(new_n796), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT113), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n809), .A2(new_n810), .A3(new_n804), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n802), .A2(new_n803), .A3(new_n808), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n808), .A2(new_n811), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n799), .A2(new_n644), .A3(new_n801), .ZN(new_n814));
  OAI21_X1  g613(.A(KEYINPUT114), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n812), .A2(new_n815), .A3(new_n687), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n541), .A2(new_n543), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n817), .B1(new_n547), .B2(new_n496), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n493), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n553), .A2(new_n645), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n595), .B1(new_n816), .B2(new_n820), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n553), .A2(new_n819), .ZN(new_n822));
  AND4_X1   g621(.A1(new_n595), .A2(new_n815), .A3(new_n812), .A4(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n622), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n623), .A2(new_n688), .A3(new_n646), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n826), .A2(new_n482), .A3(new_n649), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n653), .ZN(new_n828));
  OAI21_X1  g627(.A(G113gat), .B1(new_n828), .B2(new_n557), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n687), .A2(new_n331), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n828), .B2(new_n830), .ZN(G1340gat));
  NOR2_X1   g630(.A1(new_n828), .A2(new_n646), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(new_n329), .ZN(G1341gat));
  NOR2_X1   g632(.A1(new_n828), .A2(new_n622), .ZN(new_n834));
  NOR2_X1   g633(.A1(KEYINPUT115), .A2(G127gat), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n834), .B(new_n835), .ZN(G1342gat));
  INV_X1    g635(.A(G134gat), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n595), .A2(new_n653), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT116), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n827), .A2(new_n837), .A3(new_n840), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n841), .B(KEYINPUT56), .Z(new_n842));
  NAND3_X1  g641(.A1(new_n827), .A2(new_n653), .A3(new_n595), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n843), .A2(KEYINPUT117), .A3(G134gat), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT117), .B1(new_n843), .B2(G134gat), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(G1343gat));
  NAND2_X1  g645(.A1(new_n826), .A2(new_n424), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(KEYINPUT57), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n661), .A2(new_n653), .A3(new_n649), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n801), .A2(new_n644), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n852));
  XNOR2_X1  g651(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n809), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n851), .A2(new_n852), .A3(new_n799), .A4(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n799), .A2(new_n854), .A3(new_n644), .A4(new_n801), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT120), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n855), .B(new_n857), .C1(new_n554), .C2(new_n555), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n820), .B(KEYINPUT118), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n595), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n622), .B1(new_n860), .B2(new_n823), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n425), .B1(new_n861), .B2(new_n825), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n850), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n848), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(G141gat), .B1(new_n865), .B2(new_n688), .ZN(new_n866));
  INV_X1    g665(.A(new_n826), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n867), .A2(new_n691), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n735), .A2(new_n425), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n557), .A2(G141gat), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n868), .A2(new_n653), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT58), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT58), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(G141gat), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n848), .A2(new_n864), .A3(new_n557), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n875), .B(KEYINPUT121), .C1(new_n876), .C2(new_n877), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n873), .A2(new_n880), .A3(new_n881), .ZN(G1344gat));
  NAND2_X1  g681(.A1(new_n868), .A2(new_n869), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n883), .A2(new_n654), .ZN(new_n884));
  INV_X1    g683(.A(G148gat), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n885), .A3(new_n645), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT124), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n858), .A2(new_n859), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n671), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n813), .A2(new_n814), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n595), .A2(new_n891), .A3(new_n822), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n742), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n647), .A2(new_n556), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n888), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n892), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n622), .B1(new_n860), .B2(new_n896), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n897), .B(KEYINPUT124), .C1(new_n556), .C2(new_n647), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n425), .A2(KEYINPUT57), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n895), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n847), .A2(KEYINPUT57), .ZN(new_n901));
  XOR2_X1   g700(.A(new_n849), .B(KEYINPUT123), .Z(new_n902));
  AND4_X1   g701(.A1(new_n645), .A2(new_n900), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n885), .B1(new_n903), .B2(KEYINPUT125), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n900), .A2(new_n901), .A3(new_n902), .A4(new_n645), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT125), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n887), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n885), .A2(KEYINPUT59), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n909), .B(new_n910), .C1(new_n865), .C2(new_n646), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n848), .A2(new_n864), .A3(new_n646), .ZN(new_n912));
  INV_X1    g711(.A(new_n910), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT122), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n886), .B1(new_n908), .B2(new_n915), .ZN(G1345gat));
  OAI21_X1  g715(.A(G155gat), .B1(new_n865), .B2(new_n622), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n884), .A2(new_n320), .A3(new_n742), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1346gat));
  OAI21_X1  g718(.A(G162gat), .B1(new_n865), .B2(new_n671), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n840), .A2(new_n321), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n883), .B2(new_n921), .ZN(G1347gat));
  NAND4_X1  g721(.A1(new_n826), .A2(new_n654), .A3(new_n482), .A4(new_n691), .ZN(new_n923));
  OAI21_X1  g722(.A(G169gat), .B1(new_n923), .B2(new_n557), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n687), .A2(new_n435), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n923), .B2(new_n925), .ZN(G1348gat));
  NOR2_X1   g725(.A1(new_n923), .A2(new_n646), .ZN(new_n927));
  XOR2_X1   g726(.A(new_n927), .B(G176gat), .Z(G1349gat));
  NOR2_X1   g727(.A1(new_n923), .A2(new_n622), .ZN(new_n929));
  MUX2_X1   g728(.A(new_n238), .B(new_n249), .S(new_n929), .Z(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT60), .ZN(G1350gat));
  NOR2_X1   g730(.A1(new_n923), .A2(new_n671), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n933));
  AOI211_X1 g732(.A(new_n250), .B(new_n932), .C1(new_n933), .C2(KEYINPUT61), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n934), .B1(new_n933), .B2(KEYINPUT61), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n936));
  OAI211_X1 g735(.A(KEYINPUT126), .B(new_n936), .C1(new_n932), .C2(new_n250), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n932), .A2(new_n250), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n935), .A2(new_n937), .A3(new_n938), .ZN(G1351gat));
  NOR3_X1   g738(.A1(new_n735), .A2(new_n653), .A3(new_n649), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n826), .A2(new_n940), .A3(new_n424), .ZN(new_n941));
  INV_X1    g740(.A(G197gat), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n941), .A2(new_n942), .A3(new_n687), .ZN(new_n943));
  XOR2_X1   g742(.A(new_n943), .B(KEYINPUT127), .Z(new_n944));
  AND2_X1   g743(.A1(new_n900), .A2(new_n901), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(new_n940), .ZN(new_n946));
  OAI21_X1  g745(.A(G197gat), .B1(new_n946), .B2(new_n557), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n944), .A2(new_n947), .ZN(G1352gat));
  INV_X1    g747(.A(G204gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n941), .A2(new_n949), .A3(new_n645), .ZN(new_n950));
  XOR2_X1   g749(.A(new_n950), .B(KEYINPUT62), .Z(new_n951));
  AND3_X1   g750(.A1(new_n945), .A2(new_n645), .A3(new_n940), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n949), .B2(new_n952), .ZN(G1353gat));
  NAND3_X1  g752(.A1(new_n941), .A2(new_n269), .A3(new_n742), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n945), .A2(new_n742), .A3(new_n940), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n955), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n956));
  AOI21_X1  g755(.A(KEYINPUT63), .B1(new_n955), .B2(G211gat), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(G1354gat));
  OAI21_X1  g757(.A(G218gat), .B1(new_n946), .B2(new_n671), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n941), .A2(new_n270), .A3(new_n595), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(G1355gat));
endmodule


