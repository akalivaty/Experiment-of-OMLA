//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 1 1 1 0 0 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n571, new_n573,
    new_n574, new_n575, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n625,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1180, new_n1181, new_n1182, new_n1183;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n458), .A2(KEYINPUT65), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n458), .A2(KEYINPUT65), .B1(G567), .B2(new_n454), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G125), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n467), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n472), .A2(KEYINPUT67), .A3(G125), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n466), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT68), .B1(new_n470), .B2(G2104), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n479), .A2(new_n468), .A3(KEYINPUT3), .ZN(new_n480));
  AND3_X1   g055(.A1(new_n478), .A2(new_n480), .A3(new_n471), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n481), .A2(G137), .A3(new_n466), .ZN(new_n482));
  INV_X1    g057(.A(G101), .ZN(new_n483));
  INV_X1    g058(.A(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2104), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n482), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n477), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT69), .ZN(G160));
  NAND3_X1  g063(.A1(new_n478), .A2(new_n480), .A3(new_n471), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT70), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(new_n484), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G136), .ZN(new_n493));
  INV_X1    g068(.A(new_n466), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G124), .ZN(new_n496));
  NOR2_X1   g071(.A1(G100), .A2(G2105), .ZN(new_n497));
  XNOR2_X1  g072(.A(new_n497), .B(KEYINPUT71), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n499));
  XNOR2_X1  g074(.A(new_n499), .B(KEYINPUT72), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n493), .A2(new_n496), .A3(new_n500), .ZN(new_n501));
  XOR2_X1   g076(.A(new_n501), .B(KEYINPUT73), .Z(G162));
  NAND3_X1  g077(.A1(new_n481), .A2(G126), .A3(G2105), .ZN(new_n503));
  OR2_X1    g078(.A1(G102), .A2(G2105), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n504), .B(G2104), .C1(G114), .C2(new_n484), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G138), .ZN(new_n507));
  NOR3_X1   g082(.A1(new_n464), .A2(new_n465), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(KEYINPUT4), .B1(new_n508), .B2(new_n472), .ZN(new_n509));
  OR2_X1    g084(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n510));
  NAND4_X1  g085(.A1(new_n510), .A2(KEYINPUT4), .A3(G138), .A4(new_n463), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n489), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(G164));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  OAI21_X1  g091(.A(KEYINPUT74), .B1(new_n516), .B2(G651), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT74), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n518), .A2(new_n519), .A3(KEYINPUT6), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n516), .A2(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OR2_X1    g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G88), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n526), .A2(G62), .ZN(new_n530));
  INV_X1    g105(.A(G75), .ZN(new_n531));
  INV_X1    g106(.A(G543), .ZN(new_n532));
  OAI21_X1  g107(.A(KEYINPUT75), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OR3_X1    g108(.A1(new_n531), .A2(new_n532), .A3(KEYINPUT75), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n530), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G651), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n517), .A2(new_n520), .B1(new_n516), .B2(G651), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n537), .A2(G50), .A3(G543), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n529), .A2(new_n536), .A3(new_n538), .ZN(G303));
  INV_X1    g114(.A(G303), .ZN(G166));
  INV_X1    g115(.A(KEYINPUT76), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n523), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n537), .A2(KEYINPUT76), .ZN(new_n543));
  AND3_X1   g118(.A1(new_n542), .A2(G543), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G51), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n528), .A2(G89), .ZN(new_n546));
  NAND3_X1  g121(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(KEYINPUT7), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(KEYINPUT7), .ZN(new_n549));
  AND2_X1   g124(.A1(G63), .A2(G651), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n548), .A2(new_n549), .B1(new_n526), .B2(new_n550), .ZN(new_n551));
  AND2_X1   g126(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n545), .A2(new_n552), .ZN(G286));
  INV_X1    g128(.A(G286), .ZN(G168));
  AOI22_X1  g129(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(new_n519), .ZN(new_n556));
  XOR2_X1   g131(.A(new_n556), .B(KEYINPUT77), .Z(new_n557));
  INV_X1    g132(.A(G90), .ZN(new_n558));
  INV_X1    g133(.A(new_n528), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AND2_X1   g135(.A1(new_n544), .A2(G52), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n560), .A2(new_n561), .ZN(G171));
  NAND2_X1  g137(.A1(new_n544), .A2(G43), .ZN(new_n563));
  NAND2_X1  g138(.A1(G68), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G56), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n527), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n528), .A2(G81), .B1(new_n566), .B2(G651), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(G153));
  AND3_X1   g145(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G36), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT78), .ZN(G188));
  INV_X1    g151(.A(G91), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n526), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n578));
  OAI22_X1  g153(.A1(new_n559), .A2(new_n577), .B1(new_n578), .B2(new_n519), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n542), .A2(G53), .A3(new_n543), .A4(G543), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(KEYINPUT9), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(KEYINPUT9), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n579), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G299));
  INV_X1    g159(.A(G171), .ZN(G301));
  NAND2_X1  g160(.A1(new_n544), .A2(G49), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n526), .A2(G74), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n528), .A2(G87), .B1(G651), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n586), .A2(new_n588), .ZN(G288));
  AOI22_X1  g164(.A1(new_n526), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(new_n523), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n526), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n592), .A2(new_n519), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n593), .ZN(G305));
  NAND2_X1  g169(.A1(new_n544), .A2(G47), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n528), .A2(G85), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  OAI211_X1 g172(.A(new_n595), .B(new_n596), .C1(new_n519), .C2(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n521), .A2(G92), .A3(new_n522), .A4(new_n526), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT80), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT79), .ZN(new_n604));
  NAND4_X1  g179(.A1(new_n537), .A2(KEYINPUT80), .A3(G92), .A4(new_n526), .ZN(new_n605));
  AND3_X1   g180(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n604), .B1(new_n603), .B2(new_n605), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n603), .A2(new_n605), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(KEYINPUT79), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n610), .A2(KEYINPUT10), .A3(new_n611), .ZN(new_n612));
  NAND4_X1  g187(.A1(new_n542), .A2(G54), .A3(new_n543), .A4(G543), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n526), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n614), .A2(new_n519), .ZN(new_n615));
  AND3_X1   g190(.A1(new_n613), .A2(KEYINPUT81), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g191(.A(KEYINPUT81), .B1(new_n613), .B2(new_n615), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n608), .B(new_n612), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n599), .B1(new_n619), .B2(G868), .ZN(G321));
  XNOR2_X1  g195(.A(G321), .B(KEYINPUT82), .ZN(G284));
  NAND2_X1  g196(.A1(G286), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(new_n583), .B2(G868), .ZN(G297));
  OAI21_X1  g198(.A(new_n622), .B1(new_n583), .B2(G868), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n619), .B1(new_n625), .B2(G860), .ZN(G148));
  NOR2_X1   g201(.A1(new_n569), .A2(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n619), .A2(new_n625), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G868), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT83), .Z(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g206(.A(new_n485), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n472), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT12), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2100), .ZN(new_n636));
  OAI221_X1 g211(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n466), .C2(G111), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n490), .A2(new_n494), .ZN(new_n638));
  INV_X1    g213(.A(G123), .ZN(new_n639));
  INV_X1    g214(.A(G135), .ZN(new_n640));
  OAI221_X1 g215(.A(new_n637), .B1(new_n638), .B2(new_n639), .C1(new_n640), .C2(new_n491), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(G2096), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(G2096), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n636), .A2(new_n642), .A3(new_n643), .ZN(G156));
  XOR2_X1   g219(.A(KEYINPUT15), .B(G2435), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2427), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT84), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n646), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(KEYINPUT14), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2451), .B(G2454), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n651), .B(new_n655), .Z(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(new_n659), .A3(G14), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT85), .ZN(G401));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g239(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  AOI21_X1  g241(.A(KEYINPUT18), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n664), .B2(KEYINPUT18), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n667), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2096), .B(G2100), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1971), .B(G1976), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1956), .B(G2474), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1961), .B(G1966), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n674), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n674), .A2(new_n677), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  AOI211_X1 g257(.A(new_n679), .B(new_n682), .C1(new_n674), .C2(new_n678), .ZN(new_n683));
  XOR2_X1   g258(.A(G1991), .B(G1996), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1981), .B(G1986), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT87), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n685), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G229));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G25), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT88), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n495), .A2(G119), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT89), .ZN(new_n696));
  OAI21_X1  g271(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n697));
  INV_X1    g272(.A(G107), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n697), .B1(new_n494), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n492), .B2(G131), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n694), .B1(new_n701), .B2(G29), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT90), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT35), .B(G1991), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G288), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n707), .B2(G23), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT33), .B(G1976), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  MUX2_X1   g286(.A(G6), .B(G305), .S(G16), .Z(new_n712));
  XOR2_X1   g287(.A(KEYINPUT32), .B(G1981), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n709), .A2(new_n710), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n707), .A2(G22), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G166), .B2(new_n707), .ZN(new_n717));
  INV_X1    g292(.A(G1971), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n711), .A2(new_n714), .A3(new_n715), .A4(new_n719), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n720), .A2(KEYINPUT34), .ZN(new_n721));
  NOR2_X1   g296(.A1(G16), .A2(G24), .ZN(new_n722));
  XNOR2_X1  g297(.A(G290), .B(KEYINPUT91), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(G16), .ZN(new_n724));
  INV_X1    g299(.A(G1986), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n720), .A2(KEYINPUT34), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n705), .A2(new_n721), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT36), .Z(new_n729));
  NAND2_X1  g304(.A1(G168), .A2(G16), .ZN(new_n730));
  NOR2_X1   g305(.A1(G16), .A2(G21), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(KEYINPUT95), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(KEYINPUT95), .B2(new_n730), .ZN(new_n733));
  INV_X1    g308(.A(G1966), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G2072), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT25), .Z(new_n738));
  AOI22_X1  g313(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n739));
  INV_X1    g314(.A(G139), .ZN(new_n740));
  OAI221_X1 g315(.A(new_n738), .B1(new_n466), .B2(new_n739), .C1(new_n491), .C2(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT94), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n742), .A2(new_n692), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n692), .B2(G33), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n735), .B1(new_n736), .B2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT96), .ZN(new_n746));
  NAND2_X1  g321(.A1(G160), .A2(G29), .ZN(new_n747));
  INV_X1    g322(.A(G34), .ZN(new_n748));
  AOI21_X1  g323(.A(G29), .B1(new_n748), .B2(KEYINPUT24), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(KEYINPUT24), .B2(new_n748), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G2084), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n707), .A2(G5), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G171), .B2(new_n707), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n692), .A2(G32), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n495), .A2(G129), .ZN(new_n757));
  NAND3_X1  g332(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT26), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n760), .A2(new_n761), .B1(G105), .B2(new_n632), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G141), .B2(new_n492), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n756), .B1(new_n764), .B2(new_n692), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT27), .B(G1996), .ZN(new_n767));
  OAI221_X1 g342(.A(new_n753), .B1(G1961), .B2(new_n755), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  OAI221_X1 g343(.A(new_n745), .B1(new_n746), .B2(new_n768), .C1(new_n736), .C2(new_n744), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n768), .A2(new_n746), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n707), .A2(G4), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n619), .B2(new_n707), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT92), .B(G1348), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n772), .B(new_n773), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n692), .A2(G26), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT28), .Z(new_n776));
  OAI221_X1 g351(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n466), .C2(G116), .ZN(new_n777));
  INV_X1    g352(.A(G128), .ZN(new_n778));
  INV_X1    g353(.A(G140), .ZN(new_n779));
  OAI221_X1 g354(.A(new_n777), .B1(new_n638), .B2(new_n778), .C1(new_n779), .C2(new_n491), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n776), .B1(new_n780), .B2(G29), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT93), .B(G2067), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n751), .A2(new_n752), .ZN(new_n784));
  AOI211_X1 g359(.A(new_n783), .B(new_n784), .C1(new_n766), .C2(new_n767), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT98), .B(KEYINPUT23), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n707), .A2(G20), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n583), .B2(new_n707), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(G1956), .Z(new_n790));
  NAND2_X1  g365(.A1(new_n707), .A2(G19), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n569), .B2(new_n707), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G1341), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n755), .B2(G1961), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n692), .A2(G27), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G164), .B2(new_n692), .ZN(new_n796));
  INV_X1    g371(.A(G2078), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT31), .B(G11), .Z(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT30), .B(G28), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n799), .B1(new_n692), .B2(new_n800), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n798), .B(new_n801), .C1(new_n692), .C2(new_n641), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n782), .B2(new_n781), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n785), .A2(new_n790), .A3(new_n794), .A4(new_n803), .ZN(new_n804));
  NOR4_X1   g379(.A1(new_n769), .A2(new_n770), .A3(new_n774), .A4(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(G29), .A2(G35), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G162), .B2(G29), .ZN(new_n807));
  INV_X1    g382(.A(G2090), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT97), .B(KEYINPUT29), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n805), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n729), .A2(new_n812), .ZN(G311));
  OR2_X1    g388(.A1(new_n729), .A2(new_n812), .ZN(G150));
  XNOR2_X1  g389(.A(KEYINPUT100), .B(G55), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n544), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(G80), .A2(G543), .ZN(new_n817));
  INV_X1    g392(.A(G67), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n527), .B2(new_n818), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n528), .A2(G93), .B1(new_n819), .B2(G651), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G860), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT37), .Z(new_n823));
  NOR2_X1   g398(.A1(new_n618), .A2(new_n625), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n568), .A2(new_n821), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n568), .A2(new_n821), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n826), .B(new_n830), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n831), .A2(KEYINPUT39), .ZN(new_n832));
  INV_X1    g407(.A(G860), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n831), .B2(KEYINPUT39), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n823), .B1(new_n832), .B2(new_n834), .ZN(G145));
  INV_X1    g410(.A(KEYINPUT103), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n701), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n492), .A2(G142), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n495), .A2(G130), .ZN(new_n839));
  OAI221_X1 g414(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n466), .C2(G118), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n837), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n701), .B(KEYINPUT103), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(new_n841), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n634), .B(KEYINPUT102), .Z(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n843), .A2(new_n845), .A3(new_n847), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n503), .A2(new_n505), .ZN(new_n852));
  OAI21_X1  g427(.A(KEYINPUT101), .B1(new_n509), .B2(new_n512), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT4), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n510), .A2(G138), .A3(new_n463), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n469), .A2(new_n471), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT101), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n857), .B(new_n858), .C1(new_n489), .C2(new_n511), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n852), .B1(new_n853), .B2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n780), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n764), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(new_n741), .ZN(new_n863));
  INV_X1    g438(.A(new_n742), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n851), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(G160), .B(new_n641), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(G162), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n865), .A2(new_n863), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n849), .A2(new_n869), .A3(new_n850), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n866), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n868), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n849), .A2(new_n869), .A3(new_n850), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n869), .B1(new_n849), .B2(new_n850), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(G37), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n871), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g453(.A(KEYINPUT104), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n618), .A2(new_n879), .A3(new_n583), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n879), .B1(new_n618), .B2(new_n583), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n618), .A2(new_n583), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT41), .ZN(new_n883));
  NOR4_X1   g458(.A1(new_n880), .A2(new_n881), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(KEYINPUT105), .B1(new_n880), .B2(new_n881), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n608), .A2(new_n612), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n616), .A2(new_n617), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n583), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(KEYINPUT104), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT105), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n618), .A2(new_n879), .A3(new_n583), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n882), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n885), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n884), .B1(new_n894), .B2(new_n883), .ZN(new_n895));
  XOR2_X1   g470(.A(new_n628), .B(new_n830), .Z(new_n896));
  OR2_X1    g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n889), .A2(new_n891), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n898), .A2(new_n882), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(G290), .B(G305), .ZN(new_n902));
  XNOR2_X1  g477(.A(G288), .B(G166), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n902), .B(new_n903), .ZN(new_n904));
  XOR2_X1   g479(.A(new_n904), .B(KEYINPUT42), .Z(new_n905));
  NAND3_X1  g480(.A1(new_n897), .A2(new_n901), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n905), .B1(new_n897), .B2(new_n901), .ZN(new_n908));
  OAI21_X1  g483(.A(G868), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n821), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n909), .B1(G868), .B2(new_n910), .ZN(G295));
  OAI21_X1  g486(.A(new_n909), .B1(G868), .B2(new_n910), .ZN(G331));
  INV_X1    g487(.A(new_n829), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n913), .A2(G286), .A3(new_n827), .ZN(new_n914));
  OAI21_X1  g489(.A(G168), .B1(new_n828), .B2(new_n829), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(G301), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n914), .A2(new_n915), .A3(G171), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n900), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(new_n895), .B2(new_n919), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n904), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n923));
  INV_X1    g498(.A(new_n904), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n924), .B(new_n920), .C1(new_n895), .C2(new_n919), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n922), .A2(new_n923), .A3(new_n876), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT108), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n925), .A2(new_n876), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n928), .A2(new_n929), .A3(new_n923), .A4(new_n922), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n917), .A2(new_n918), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n932), .A2(KEYINPUT41), .A3(new_n894), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n899), .B1(new_n919), .B2(new_n883), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(new_n904), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n935), .A2(new_n925), .A3(new_n876), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT109), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(new_n937), .A3(KEYINPUT43), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n939), .B1(new_n940), .B2(KEYINPUT109), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n931), .A2(new_n938), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n882), .B1(new_n898), .B2(KEYINPUT105), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT41), .B1(new_n943), .B2(new_n892), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n932), .B1(new_n944), .B2(new_n884), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n924), .B1(new_n945), .B2(new_n920), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n925), .A2(new_n876), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT43), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT106), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n922), .A2(new_n876), .A3(new_n925), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT106), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n951), .A3(KEYINPUT43), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n953), .B1(new_n936), .B2(KEYINPUT43), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n928), .A2(KEYINPUT107), .A3(new_n923), .A4(new_n935), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n949), .A2(new_n952), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n942), .B1(new_n956), .B2(KEYINPUT44), .ZN(G397));
  XOR2_X1   g532(.A(new_n780), .B(G2067), .Z(new_n958));
  XNOR2_X1  g533(.A(new_n764), .B(G1996), .ZN(new_n959));
  OR2_X1    g534(.A1(new_n701), .A2(new_n704), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n701), .A2(new_n704), .ZN(new_n961));
  AND4_X1   g536(.A1(new_n958), .A2(new_n959), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  XOR2_X1   g537(.A(KEYINPUT110), .B(G1384), .Z(new_n963));
  NOR2_X1   g538(.A1(new_n860), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n964), .A2(KEYINPUT45), .ZN(new_n965));
  INV_X1    g540(.A(G40), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n477), .A2(new_n966), .A3(new_n486), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  OR2_X1    g543(.A1(new_n962), .A2(new_n968), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n968), .A2(G1986), .A3(G290), .ZN(new_n970));
  XOR2_X1   g545(.A(new_n970), .B(KEYINPUT48), .Z(new_n971));
  INV_X1    g546(.A(new_n968), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n959), .A2(new_n958), .ZN(new_n973));
  OAI22_X1  g548(.A1(new_n973), .A2(new_n960), .B1(G2067), .B2(new_n780), .ZN(new_n974));
  AOI22_X1  g549(.A1(new_n969), .A2(new_n971), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n968), .B1(new_n958), .B2(new_n764), .ZN(new_n976));
  INV_X1    g551(.A(G1996), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT46), .B1(new_n972), .B2(new_n977), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n972), .A2(KEYINPUT46), .A3(new_n977), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n976), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n980), .B(new_n981), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n975), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n984));
  INV_X1    g559(.A(G8), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n509), .A2(new_n512), .A3(KEYINPUT101), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n480), .A2(new_n471), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n987), .A2(new_n508), .A3(KEYINPUT4), .A4(new_n478), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n858), .B1(new_n988), .B2(new_n857), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n506), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G1384), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(KEYINPUT112), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(new_n860), .B2(G1384), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n992), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n514), .A2(KEYINPUT45), .A3(new_n991), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n997), .A2(new_n967), .ZN(new_n998));
  AOI21_X1  g573(.A(G1966), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(KEYINPUT117), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT117), .ZN(new_n1001));
  AOI211_X1 g576(.A(new_n1001), .B(G1966), .C1(new_n996), .C2(new_n998), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT50), .B1(new_n992), .B2(new_n994), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1384), .B1(new_n506), .B2(new_n513), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n967), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n1003), .A2(G2084), .A3(new_n1006), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n1000), .A2(new_n1002), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n985), .B1(new_n1008), .B2(G168), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n992), .A2(new_n994), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1006), .B1(new_n1010), .B2(new_n1004), .ZN(new_n1011));
  AOI22_X1  g586(.A1(new_n999), .A2(KEYINPUT117), .B1(new_n1011), .B2(new_n752), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n996), .A2(new_n998), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n734), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n1001), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(G286), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n984), .B1(new_n1009), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(G8), .B1(new_n1016), .B2(G286), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1019), .A2(KEYINPUT51), .ZN(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT62), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1008), .A2(G168), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT51), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT62), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1009), .A2(new_n984), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(G303), .A2(G8), .ZN(new_n1027));
  XNOR2_X1  g602(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n1028));
  XOR2_X1   g603(.A(new_n1027), .B(new_n1028), .Z(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1005), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n995), .ZN(new_n1032));
  INV_X1    g607(.A(new_n963), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n990), .A2(KEYINPUT45), .A3(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1034), .A2(KEYINPUT111), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT111), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1036), .B1(new_n964), .B2(KEYINPUT45), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n967), .B(new_n1032), .C1(new_n1035), .C2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n967), .B1(new_n1031), .B2(KEYINPUT50), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n992), .A2(new_n994), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1039), .B1(new_n1040), .B2(KEYINPUT50), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n718), .A2(new_n1038), .B1(new_n1041), .B2(new_n808), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1030), .B1(new_n1042), .B2(new_n985), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n985), .B1(new_n1010), .B2(new_n967), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n1046));
  NAND2_X1  g621(.A1(G305), .A2(G1981), .ZN(new_n1047));
  INV_X1    g622(.A(G1981), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n591), .A2(new_n593), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1046), .B1(new_n1050), .B2(KEYINPUT115), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT49), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT115), .B1(new_n1046), .B2(KEYINPUT49), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1051), .A2(new_n1052), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1045), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT114), .B1(new_n706), .B2(G1976), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1044), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n706), .A2(G1976), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1044), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1044), .B(new_n1057), .C1(KEYINPUT52), .C2(new_n1059), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1056), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1011), .A2(new_n808), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n487), .A2(G40), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1034), .A2(KEYINPUT111), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n964), .A2(new_n1036), .A3(KEYINPUT45), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(G1971), .B1(new_n1070), .B2(new_n1032), .ZN(new_n1071));
  OAI211_X1 g646(.A(G8), .B(new_n1029), .C1(new_n1066), .C2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1043), .A2(new_n1064), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1961), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1074), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1076), .A2(G2078), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n996), .A2(new_n1077), .A3(new_n998), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT123), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT123), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1075), .A2(new_n1081), .A3(new_n1078), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1070), .A2(new_n797), .A3(new_n1032), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1080), .A2(new_n1082), .B1(new_n1076), .B2(new_n1083), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1073), .A2(G301), .A3(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1021), .A2(new_n1026), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1038), .A2(new_n718), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n985), .B1(new_n1087), .B2(new_n1065), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1064), .A2(new_n1029), .A3(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(G288), .A2(G1976), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n1055), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1049), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1044), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1089), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT63), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT118), .ZN(new_n1096));
  NOR2_X1   g671(.A1(G286), .A2(new_n985), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1096), .B1(new_n1016), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1097), .ZN(new_n1099));
  AOI211_X1 g674(.A(KEYINPUT118), .B(new_n1099), .C1(new_n1012), .C2(new_n1015), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1095), .B1(new_n1101), .B2(new_n1073), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1064), .A2(new_n1072), .ZN(new_n1103));
  OAI21_X1  g678(.A(KEYINPUT63), .B1(new_n1088), .B2(new_n1029), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT118), .B1(new_n1008), .B2(new_n1099), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1016), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1094), .B1(new_n1102), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1086), .A2(new_n1110), .ZN(new_n1111));
  OR2_X1    g686(.A1(new_n1041), .A2(G1956), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n583), .B(KEYINPUT57), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT56), .B(G2072), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1070), .A2(new_n1032), .A3(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1112), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n1117), .A2(KEYINPUT122), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n1117), .B2(KEYINPUT122), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1113), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1121));
  OR2_X1    g696(.A1(new_n1121), .A2(KEYINPUT120), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(KEYINPUT120), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1118), .A2(new_n1120), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1010), .A2(new_n967), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT58), .B(G1341), .Z(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n1038), .B2(G1996), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n569), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1129), .B(KEYINPUT59), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1125), .A2(G2067), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1011), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1131), .B1(new_n773), .B2(new_n1132), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1133), .A2(new_n618), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1133), .A2(new_n618), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT60), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT60), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1133), .A2(new_n1137), .A3(new_n619), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1130), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1119), .B1(new_n1117), .B2(new_n1121), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1140), .A2(KEYINPUT121), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1140), .A2(KEYINPUT121), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1124), .B(new_n1139), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT119), .B1(new_n1133), .B2(new_n618), .ZN(new_n1144));
  OR3_X1    g719(.A1(new_n1133), .A2(KEYINPUT119), .A3(new_n618), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1122), .A2(new_n1123), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n1116), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1083), .A2(new_n1076), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1070), .B(new_n1077), .C1(KEYINPUT45), .C2(new_n964), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1150), .A2(G301), .A3(new_n1075), .A4(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1152), .B1(new_n1084), .B2(G301), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT54), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1073), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1149), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1150), .A2(new_n1075), .A3(new_n1151), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1154), .B1(new_n1157), .B2(G171), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1082), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1081), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1160));
  OAI211_X1 g735(.A(G301), .B(new_n1150), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1161), .A2(KEYINPUT124), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1161), .A2(KEYINPUT124), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1158), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(KEYINPUT125), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1166), .B(new_n1158), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1156), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1111), .B1(new_n1148), .B2(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(G290), .B(new_n725), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n968), .B1(new_n962), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n983), .B1(new_n1169), .B2(new_n1171), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g747(.A1(new_n461), .A2(G227), .ZN(new_n1174));
  NOR2_X1   g748(.A1(new_n1174), .A2(KEYINPUT127), .ZN(new_n1175));
  AND2_X1   g749(.A1(new_n1174), .A2(KEYINPUT127), .ZN(new_n1176));
  NOR4_X1   g750(.A1(G229), .A2(G401), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  NAND2_X1  g751(.A1(new_n877), .A2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g752(.A1(new_n956), .A2(new_n1178), .ZN(G308));
  NAND2_X1  g753(.A1(new_n955), .A2(new_n954), .ZN(new_n1180));
  INV_X1    g754(.A(new_n952), .ZN(new_n1181));
  AOI21_X1  g755(.A(new_n951), .B1(new_n950), .B2(KEYINPUT43), .ZN(new_n1182));
  OAI21_X1  g756(.A(new_n1180), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g757(.A1(new_n1183), .A2(new_n877), .A3(new_n1177), .ZN(G225));
endmodule


