//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 1 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0 1 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n557,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n576, new_n577, new_n578, new_n579, new_n580, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1187, new_n1188, new_n1189;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G69), .Z(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  NAND2_X1  g033(.A1(G113), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(G101), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  OR2_X1    g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n475), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G124), .ZN(new_n479));
  INV_X1    g054(.A(G136), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n477), .A2(new_n471), .ZN(new_n481));
  OAI221_X1 g056(.A(new_n476), .B1(new_n478), .B2(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  NOR2_X1   g058(.A1(new_n460), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G102), .ZN(new_n485));
  NAND2_X1  g060(.A1(G114), .A2(G2104), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n487), .B1(new_n477), .B2(G126), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n485), .B1(new_n488), .B2(new_n471), .ZN(new_n489));
  AND2_X1   g064(.A1(KEYINPUT67), .A2(G138), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n461), .A2(new_n463), .A3(new_n490), .A4(new_n471), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n477), .A2(KEYINPUT4), .A3(new_n471), .A4(new_n490), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n489), .A2(new_n495), .ZN(G164));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(KEYINPUT68), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(KEYINPUT5), .A3(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AND3_X1   g077(.A1(new_n502), .A2(KEYINPUT69), .A3(G62), .ZN(new_n503));
  AOI21_X1  g078(.A(KEYINPUT69), .B1(new_n502), .B2(G62), .ZN(new_n504));
  NAND2_X1  g079(.A1(G75), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  NOR3_X1   g081(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(new_n508), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n502), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n507), .A2(new_n508), .B1(new_n513), .B2(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  NAND3_X1  g091(.A1(new_n502), .A2(G89), .A3(new_n512), .ZN(new_n517));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT7), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n517), .A2(KEYINPUT72), .A3(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g096(.A(KEYINPUT72), .B1(new_n517), .B2(new_n519), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  INV_X1    g099(.A(new_n511), .ZN(new_n525));
  NOR2_X1   g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  OAI21_X1  g101(.A(KEYINPUT70), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n510), .A2(new_n528), .A3(new_n511), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n527), .A2(G543), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT71), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT71), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n527), .A2(new_n529), .A3(new_n532), .A4(G543), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n524), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n502), .A2(G63), .A3(G651), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  NOR3_X1   g111(.A1(new_n523), .A2(new_n534), .A3(new_n536), .ZN(G168));
  XNOR2_X1  g112(.A(KEYINPUT73), .B(G52), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n538), .B1(new_n531), .B2(new_n533), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n502), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n502), .A2(new_n512), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n540), .A2(new_n508), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n539), .A2(new_n543), .ZN(G171));
  AOI22_X1  g119(.A1(new_n502), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n546), .A2(KEYINPUT74), .A3(G651), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT74), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n548), .B1(new_n545), .B2(new_n508), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n551), .B1(new_n531), .B2(new_n533), .ZN(new_n552));
  INV_X1    g127(.A(new_n542), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n553), .A2(G81), .ZN(new_n554));
  NOR3_X1   g129(.A1(new_n550), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  NAND4_X1  g136(.A1(new_n527), .A2(new_n529), .A3(G53), .A4(G543), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT9), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(new_n499), .B2(new_n501), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT75), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n566), .B(new_n567), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT76), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n571));
  OAI211_X1 g146(.A(new_n571), .B(G651), .C1(new_n565), .C2(new_n568), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n553), .A2(G91), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n563), .A2(new_n573), .A3(new_n574), .ZN(G299));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n576), .B1(new_n539), .B2(new_n543), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NOR3_X1   g153(.A1(new_n539), .A2(new_n576), .A3(new_n543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G301));
  NAND2_X1  g156(.A1(new_n531), .A2(new_n533), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G51), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n583), .B(new_n535), .C1(new_n522), .C2(new_n521), .ZN(G286));
  NAND3_X1  g159(.A1(new_n502), .A2(G87), .A3(new_n512), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT78), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT80), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g164(.A(KEYINPUT80), .B(G651), .C1(new_n502), .C2(G74), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n527), .A2(new_n529), .A3(G49), .A4(G543), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n592), .A2(KEYINPUT79), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n592), .A2(KEYINPUT79), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n586), .B(new_n591), .C1(new_n593), .C2(new_n594), .ZN(G288));
  AND3_X1   g170(.A1(new_n512), .A2(G48), .A3(G543), .ZN(new_n596));
  INV_X1    g171(.A(G61), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n597), .B1(new_n499), .B2(new_n501), .ZN(new_n598));
  AND2_X1   g173(.A1(G73), .A2(G543), .ZN(new_n599));
  OAI21_X1  g174(.A(G651), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT81), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g177(.A(KEYINPUT81), .B(G651), .C1(new_n598), .C2(new_n599), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n596), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n553), .A2(G86), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(G305));
  AOI22_X1  g181(.A1(new_n582), .A2(G47), .B1(G85), .B2(new_n553), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n608), .A2(new_n508), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n607), .A2(new_n609), .ZN(G290));
  AOI22_X1  g185(.A1(new_n502), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n611), .A2(new_n508), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(new_n582), .B2(G54), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n502), .A2(G92), .A3(new_n512), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT10), .Z(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(new_n580), .B2(new_n617), .ZN(G284));
  OAI21_X1  g194(.A(new_n618), .B1(new_n580), .B2(new_n617), .ZN(G321));
  NAND2_X1  g195(.A1(G299), .A2(new_n617), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n617), .B2(G168), .ZN(G297));
  OAI21_X1  g197(.A(new_n621), .B1(new_n617), .B2(G168), .ZN(G280));
  INV_X1    g198(.A(new_n616), .ZN(new_n624));
  XOR2_X1   g199(.A(KEYINPUT82), .B(G559), .Z(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(G860), .B2(new_n625), .ZN(G148));
  NOR2_X1   g201(.A1(new_n555), .A2(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n624), .A2(new_n625), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT83), .Z(new_n629));
  AOI21_X1  g204(.A(new_n627), .B1(new_n629), .B2(G868), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT84), .Z(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g207(.A1(new_n477), .A2(new_n484), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT12), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  INV_X1    g210(.A(KEYINPUT85), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G2100), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n635), .B(new_n637), .Z(new_n638));
  INV_X1    g213(.A(new_n478), .ZN(new_n639));
  INV_X1    g214(.A(new_n481), .ZN(new_n640));
  AOI22_X1  g215(.A1(G123), .A2(new_n639), .B1(new_n640), .B2(G135), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n471), .A2(G111), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT86), .Z(new_n644));
  OAI21_X1  g219(.A(new_n641), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(G2096), .Z(new_n646));
  OAI211_X1 g221(.A(new_n638), .B(new_n646), .C1(new_n636), .C2(G2100), .ZN(G156));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2435), .ZN(new_n649));
  XOR2_X1   g224(.A(G2427), .B(G2438), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT14), .ZN(new_n652));
  XOR2_X1   g227(.A(G2451), .B(G2454), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1341), .B(G1348), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT87), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n654), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n658), .B(new_n659), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(G14), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G401));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2067), .B(G2678), .Z(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT88), .B(KEYINPUT18), .Z(new_n668));
  AOI21_X1  g243(.A(new_n663), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2096), .B(G2100), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT89), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n669), .B(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT17), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n665), .B2(new_n666), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n668), .B1(new_n667), .B2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n672), .B(new_n675), .Z(G227));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n677), .A2(new_n678), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n683), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n680), .A2(new_n682), .A3(new_n684), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n687), .B(new_n688), .C1(new_n686), .C2(new_n685), .ZN(new_n689));
  XOR2_X1   g264(.A(G1981), .B(G1986), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1991), .B(G1996), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT90), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n693), .B(new_n695), .ZN(G229));
  NAND2_X1  g271(.A1(G168), .A2(G16), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G16), .B2(G21), .ZN(new_n698));
  INV_X1    g273(.A(G1966), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G35), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G162), .B2(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT100), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT29), .ZN(new_n706));
  INV_X1    g281(.A(G2090), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n706), .A2(KEYINPUT101), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(G5), .A2(G16), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G171), .B2(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G1961), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n701), .A2(G26), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n639), .A2(G128), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n640), .A2(G140), .ZN(new_n714));
  OR2_X1    g289(.A1(G104), .A2(G2105), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n715), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n713), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n712), .B1(new_n718), .B2(new_n701), .ZN(new_n719));
  MUX2_X1   g294(.A(new_n712), .B(new_n719), .S(KEYINPUT28), .Z(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT93), .B(G2067), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  AND4_X1   g297(.A1(new_n700), .A2(new_n708), .A3(new_n711), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT95), .B(KEYINPUT24), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G34), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(new_n701), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n473), .B2(new_n701), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G2084), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n701), .A2(G32), .ZN(new_n729));
  AOI22_X1  g304(.A1(G129), .A2(new_n639), .B1(new_n640), .B2(G141), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n484), .A2(G105), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT96), .B(KEYINPUT26), .ZN(new_n733));
  NAND3_X1  g308(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n729), .B1(new_n737), .B2(new_n701), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT27), .B(G1996), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G27), .ZN(new_n741));
  OAI21_X1  g316(.A(KEYINPUT99), .B1(new_n741), .B2(G29), .ZN(new_n742));
  OR3_X1    g317(.A1(new_n741), .A2(KEYINPUT99), .A3(G29), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n742), .B(new_n743), .C1(G164), .C2(new_n701), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G2078), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n624), .A2(G16), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G4), .B2(G16), .ZN(new_n747));
  INV_X1    g322(.A(G1348), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n749), .A2(new_n471), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT94), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n640), .A2(G139), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n484), .A2(G103), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT25), .Z(new_n754));
  NAND3_X1  g329(.A1(new_n751), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G29), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G29), .B2(G33), .ZN(new_n758));
  INV_X1    g333(.A(G2072), .ZN(new_n759));
  OAI221_X1 g334(.A(new_n745), .B1(new_n747), .B2(new_n748), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(G299), .A2(G16), .ZN(new_n761));
  INV_X1    g336(.A(G16), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n762), .A2(KEYINPUT23), .A3(G20), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT23), .ZN(new_n764));
  INV_X1    g339(.A(G20), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(G16), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n761), .A2(new_n763), .A3(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1956), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n760), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n723), .A2(new_n728), .A3(new_n740), .A4(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(KEYINPUT101), .B1(new_n706), .B2(new_n707), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT97), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n698), .A2(new_n699), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n747), .A2(new_n748), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n762), .A2(G19), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n555), .B2(new_n762), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1341), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n710), .A2(G1961), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT30), .B(G28), .ZN(new_n780));
  OR2_X1    g355(.A1(KEYINPUT31), .A2(G11), .ZN(new_n781));
  NAND2_X1  g356(.A1(KEYINPUT31), .A2(G11), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n780), .A2(new_n701), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n645), .B2(new_n701), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT98), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n778), .A2(new_n779), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n744), .A2(G2078), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n758), .B2(new_n759), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n774), .A2(new_n775), .A3(new_n786), .A4(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n770), .A2(new_n789), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n706), .A2(new_n707), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT36), .ZN(new_n792));
  NAND2_X1  g367(.A1(G166), .A2(G16), .ZN(new_n793));
  NOR2_X1   g368(.A1(G16), .A2(G22), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(G1971), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(G1971), .ZN(new_n797));
  AOI211_X1 g372(.A(new_n797), .B(new_n794), .C1(G166), .C2(G16), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n762), .A2(G23), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G288), .B2(G16), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT33), .B(G1976), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n762), .A2(G6), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G305), .B2(G16), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT32), .B(G1981), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT34), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n799), .A2(new_n803), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n762), .A2(G24), .ZN(new_n810));
  INV_X1    g385(.A(G290), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(new_n762), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n812), .A2(G1986), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(G1986), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n701), .A2(G25), .ZN(new_n815));
  OR2_X1    g390(.A1(G95), .A2(G2105), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n816), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n817));
  INV_X1    g392(.A(G119), .ZN(new_n818));
  INV_X1    g393(.A(G131), .ZN(new_n819));
  OAI221_X1 g394(.A(new_n817), .B1(new_n478), .B2(new_n818), .C1(new_n819), .C2(new_n481), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n815), .B1(new_n821), .B2(new_n701), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT91), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT35), .B(G1991), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n809), .A2(new_n813), .A3(new_n814), .A4(new_n825), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n826), .A2(KEYINPUT92), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(KEYINPUT92), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n799), .A2(new_n803), .A3(new_n807), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT34), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n792), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n831), .ZN(new_n833));
  AOI211_X1 g408(.A(KEYINPUT36), .B(new_n833), .C1(new_n827), .C2(new_n828), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n790), .B(new_n791), .C1(new_n832), .C2(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n773), .A2(new_n772), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(G311));
  OR2_X1    g412(.A1(new_n832), .A2(new_n834), .ZN(new_n838));
  INV_X1    g413(.A(new_n836), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n838), .A2(new_n839), .A3(new_n791), .A4(new_n790), .ZN(G150));
  AOI22_X1  g415(.A1(new_n502), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n841));
  INV_X1    g416(.A(G93), .ZN(new_n842));
  OAI22_X1  g417(.A1(new_n841), .A2(new_n508), .B1(new_n842), .B2(new_n542), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT102), .B(G55), .Z(new_n844));
  AOI21_X1  g419(.A(new_n843), .B1(new_n582), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(G860), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT37), .Z(new_n848));
  NAND2_X1  g423(.A1(new_n555), .A2(new_n846), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n552), .A2(new_n554), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n845), .B1(new_n850), .B2(new_n550), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  XOR2_X1   g427(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n624), .A2(G559), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n854), .B(new_n855), .Z(new_n856));
  OAI21_X1  g431(.A(new_n848), .B1(new_n856), .B2(G860), .ZN(G145));
  XNOR2_X1  g432(.A(new_n645), .B(new_n473), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(G162), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n820), .ZN(new_n860));
  XNOR2_X1  g435(.A(G164), .B(new_n717), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n736), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT104), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n755), .B2(KEYINPUT103), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n863), .B2(new_n755), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n862), .B(new_n863), .C1(KEYINPUT103), .C2(new_n755), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n639), .A2(G130), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n640), .A2(G142), .ZN(new_n869));
  NOR2_X1   g444(.A1(G106), .A2(G2105), .ZN(new_n870));
  OAI21_X1  g445(.A(G2104), .B1(new_n471), .B2(G118), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n868), .B(new_n869), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n634), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n866), .A2(new_n867), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n874), .B1(new_n866), .B2(new_n867), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n860), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n866), .A2(new_n867), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(new_n873), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n859), .B(new_n821), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n866), .A2(new_n867), .A3(new_n874), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(G37), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n877), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g460(.A1(new_n846), .A2(new_n617), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n629), .B(new_n852), .ZN(new_n887));
  XNOR2_X1  g462(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n616), .A2(G299), .ZN(new_n889));
  AOI22_X1  g464(.A1(new_n570), .A2(new_n572), .B1(G91), .B2(new_n553), .ZN(new_n890));
  AOI22_X1  g465(.A1(new_n613), .A2(new_n615), .B1(new_n890), .B2(new_n563), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n888), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n616), .A2(G299), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT41), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n613), .A2(new_n890), .A3(new_n563), .A4(new_n615), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n887), .A2(new_n892), .A3(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n889), .A2(new_n891), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n897), .B1(new_n887), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(G288), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(G290), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n900), .A2(G290), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT106), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(G305), .B(G303), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n811), .A2(G288), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(new_n908), .A3(new_n901), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n904), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n905), .B(KEYINPUT106), .C1(new_n902), .C2(new_n903), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n914), .B(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n899), .B(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n886), .B1(new_n917), .B2(new_n617), .ZN(G295));
  OAI21_X1  g493(.A(new_n886), .B1(new_n917), .B2(new_n617), .ZN(G331));
  NAND2_X1  g494(.A1(G171), .A2(KEYINPUT77), .ZN(new_n920));
  AOI21_X1  g495(.A(G286), .B1(new_n577), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G171), .ZN(new_n922));
  NOR2_X1   g497(.A1(G168), .A2(new_n922), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n849), .B(new_n851), .C1(new_n921), .C2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(G168), .B1(new_n578), .B2(new_n579), .ZN(new_n925));
  NAND2_X1  g500(.A1(G286), .A2(G171), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n555), .A2(new_n846), .ZN(new_n927));
  NOR3_X1   g502(.A1(new_n850), .A2(new_n550), .A3(new_n845), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n925), .B(new_n926), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n898), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n892), .A2(new_n896), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n932), .A2(new_n924), .A3(new_n929), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n883), .B1(new_n934), .B2(new_n912), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n931), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n898), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n894), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n898), .A2(new_n888), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n939), .A2(new_n924), .A3(new_n929), .A4(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n938), .B1(new_n924), .B2(new_n929), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT109), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n937), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n935), .B1(new_n912), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT111), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n944), .A2(new_n912), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n932), .A2(new_n924), .A3(new_n929), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n949), .A2(new_n942), .ZN(new_n950));
  INV_X1    g525(.A(new_n912), .ZN(new_n951));
  AOI21_X1  g526(.A(G37), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n948), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT111), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(new_n954), .A3(KEYINPUT43), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT108), .B1(new_n949), .B2(new_n942), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n931), .A2(new_n957), .A3(new_n933), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n958), .A3(new_n912), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(new_n952), .A3(new_n946), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n947), .A2(new_n955), .A3(KEYINPUT44), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n952), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n948), .A2(new_n946), .A3(new_n952), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(KEYINPUT110), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n945), .A2(new_n966), .A3(new_n946), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n961), .B1(new_n968), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g544(.A(G1986), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n811), .A2(new_n970), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n971), .B(KEYINPUT112), .Z(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1996), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n737), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G2067), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n717), .B(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n736), .A2(G1996), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n975), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n820), .A2(new_n824), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n820), .A2(new_n824), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n973), .B(new_n982), .C1(new_n970), .C2(new_n811), .ZN(new_n983));
  INV_X1    g558(.A(G1384), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(new_n489), .B2(new_n495), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n467), .A2(new_n472), .A3(G40), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n983), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n991));
  OAI211_X1 g566(.A(KEYINPUT113), .B(new_n984), .C1(new_n489), .C2(new_n495), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n461), .A2(new_n463), .A3(G126), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n486), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(G2105), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n996), .A2(new_n485), .A3(new_n493), .A4(new_n494), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT113), .B1(new_n997), .B2(new_n984), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n991), .B1(new_n993), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n988), .B1(new_n985), .B2(KEYINPUT50), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G1961), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n493), .A2(new_n494), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n995), .A2(G2105), .B1(G102), .B2(new_n484), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1384), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n988), .B1(new_n1005), .B2(KEYINPUT45), .ZN(new_n1006));
  INV_X1    g581(.A(G2078), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1006), .A2(new_n1007), .A3(new_n987), .ZN(new_n1008));
  XNOR2_X1  g583(.A(KEYINPUT124), .B(KEYINPUT53), .ZN(new_n1009));
  AOI22_X1  g584(.A1(new_n1001), .A2(new_n1002), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n985), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1012), .A2(new_n986), .A3(new_n992), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1013), .A2(new_n1007), .A3(new_n1006), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT123), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1013), .A2(KEYINPUT123), .A3(new_n1007), .A4(new_n1006), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT53), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1010), .B(G301), .C1(new_n1016), .C2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1006), .A2(KEYINPUT53), .A3(new_n1007), .A4(new_n987), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT50), .B1(new_n1012), .B2(new_n992), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1000), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1020), .B(new_n1021), .C1(new_n1024), .C2(G1961), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(G171), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n1019), .A2(KEYINPUT54), .A3(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1010), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n580), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1010), .A2(G301), .A3(new_n1021), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT54), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1027), .B1(new_n1031), .B2(KEYINPUT125), .ZN(new_n1032));
  NAND2_X1  g607(.A1(G303), .A2(G8), .ZN(new_n1033));
  XNOR2_X1  g608(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1033), .B(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1012), .A2(KEYINPUT50), .A3(new_n992), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1005), .A2(new_n991), .ZN(new_n1037));
  INV_X1    g612(.A(new_n988), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1036), .A2(new_n707), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1006), .A2(new_n987), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n797), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G8), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1035), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1981), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n604), .A2(new_n1045), .A3(new_n605), .ZN(new_n1046));
  XNOR2_X1  g621(.A(KEYINPUT115), .B(G86), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n600), .B1(new_n542), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(G1981), .B1(new_n1048), .B2(new_n596), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT49), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1012), .A2(new_n992), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1043), .B1(new_n1053), .B2(new_n1038), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1046), .A2(KEYINPUT49), .A3(new_n1049), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1052), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1038), .B1(new_n993), .B2(new_n998), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n593), .A2(new_n594), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1058), .A2(G1976), .A3(new_n586), .A4(new_n591), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1057), .A2(new_n1059), .A3(G8), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT52), .ZN(new_n1061));
  INV_X1    g636(.A(G1976), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT52), .B1(G288), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1054), .A2(new_n1059), .A3(new_n1063), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1056), .A2(new_n1061), .A3(new_n1064), .ZN(new_n1065));
  XOR2_X1   g640(.A(new_n1033), .B(new_n1034), .Z(new_n1066));
  OAI21_X1  g641(.A(new_n1041), .B1(new_n1001), .B2(G2090), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1066), .A2(new_n1067), .A3(G8), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1044), .A2(new_n1065), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT126), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT126), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1044), .A2(new_n1065), .A3(new_n1071), .A4(new_n1068), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT125), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1025), .A2(new_n580), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(new_n580), .B2(new_n1028), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1074), .B1(new_n1076), .B2(KEYINPUT54), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1013), .A2(new_n1006), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n699), .ZN(new_n1079));
  INV_X1    g654(.A(G2084), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n999), .A2(new_n1080), .A3(new_n1000), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1043), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(G286), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1079), .A2(new_n1081), .A3(G168), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT122), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1084), .A2(new_n1085), .A3(G8), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT51), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1083), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1032), .A2(new_n1073), .A3(new_n1077), .A4(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n748), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n976), .B(new_n1038), .C1(new_n993), .C2(new_n998), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT117), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1053), .A2(KEYINPUT117), .A3(new_n976), .A4(new_n1038), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1093), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT118), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1093), .A2(new_n1096), .A3(new_n1100), .A4(new_n1097), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1103));
  INV_X1    g678(.A(G1956), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1006), .A2(new_n987), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT56), .B(G2072), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1103), .A2(new_n1104), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  XOR2_X1   g682(.A(G299), .B(KEYINPUT57), .Z(new_n1108));
  AND2_X1   g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1102), .A2(new_n1109), .A3(new_n616), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1102), .A2(KEYINPUT60), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT121), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT60), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1099), .A2(new_n1116), .A3(new_n1101), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1117), .A2(new_n624), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1102), .A2(KEYINPUT121), .A3(KEYINPUT60), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1115), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1117), .A2(new_n624), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT121), .B1(new_n1102), .B2(KEYINPUT60), .ZN(new_n1122));
  AOI211_X1 g697(.A(new_n1114), .B(new_n1116), .C1(new_n1099), .C2(new_n1101), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT61), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1125), .B1(new_n1107), .B2(KEYINPUT120), .ZN(new_n1126));
  OAI211_X1 g701(.A(KEYINPUT119), .B(new_n1126), .C1(new_n1109), .C2(new_n1111), .ZN(new_n1127));
  OR2_X1    g702(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(KEYINPUT120), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1131), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1127), .B(new_n1130), .C1(new_n1132), .C2(KEYINPUT61), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1040), .A2(G1996), .ZN(new_n1134));
  XNOR2_X1  g709(.A(KEYINPUT58), .B(G1341), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1135), .B1(new_n1053), .B2(new_n1038), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n555), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1137), .B(KEYINPUT59), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1120), .A2(new_n1124), .A3(new_n1133), .A4(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1092), .B1(new_n1112), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1067), .A2(G8), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n1035), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1142), .A2(G168), .A3(new_n1068), .A4(new_n1082), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1056), .A2(new_n1061), .A3(new_n1064), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(KEYINPUT116), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT116), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1056), .A2(new_n1061), .A3(new_n1064), .A4(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT63), .B1(new_n1143), .B2(new_n1148), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1068), .A2(G168), .A3(new_n1082), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT63), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1150), .A2(new_n1151), .A3(new_n1044), .A4(new_n1065), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1056), .A2(new_n1062), .A3(new_n900), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(new_n1046), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n1054), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1149), .A2(new_n1152), .A3(new_n1155), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n1148), .A2(new_n1068), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1029), .ZN(new_n1158));
  OR2_X1    g733(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1159), .A2(new_n1088), .B1(G286), .B2(new_n1082), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT62), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1158), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1073), .B1(new_n1091), .B2(KEYINPUT62), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1156), .B(new_n1157), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n990), .B1(new_n1140), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n972), .A2(new_n989), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1166), .B(KEYINPUT48), .ZN(new_n1167));
  INV_X1    g742(.A(new_n989), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1167), .B1(new_n1168), .B2(new_n982), .ZN(new_n1169));
  INV_X1    g744(.A(new_n980), .ZN(new_n1170));
  OAI22_X1  g745(.A1(new_n979), .A2(new_n1170), .B1(G2067), .B2(new_n717), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(new_n989), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1168), .B1(new_n737), .B2(new_n977), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n989), .A2(KEYINPUT46), .A3(new_n974), .ZN(new_n1174));
  AOI21_X1  g749(.A(KEYINPUT46), .B1(new_n989), .B2(new_n974), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g751(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1176), .B(new_n1177), .ZN(new_n1178));
  AND3_X1   g753(.A1(new_n1169), .A2(new_n1172), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1165), .A2(new_n1179), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g755(.A1(new_n884), .A2(G319), .ZN(new_n1182));
  NAND4_X1  g756(.A1(new_n965), .A2(new_n661), .A3(new_n1182), .A4(new_n967), .ZN(new_n1183));
  NOR2_X1   g757(.A1(G229), .A2(G227), .ZN(new_n1184));
  INV_X1    g758(.A(new_n1184), .ZN(new_n1185));
  NOR2_X1   g759(.A1(new_n1183), .A2(new_n1185), .ZN(G308));
  AND4_X1   g760(.A1(new_n966), .A2(new_n948), .A3(new_n946), .A4(new_n952), .ZN(new_n1187));
  AOI21_X1  g761(.A(new_n966), .B1(new_n962), .B2(KEYINPUT43), .ZN(new_n1188));
  AOI21_X1  g762(.A(new_n1187), .B1(new_n964), .B2(new_n1188), .ZN(new_n1189));
  NAND4_X1  g763(.A1(new_n1189), .A2(new_n661), .A3(new_n1184), .A4(new_n1182), .ZN(G225));
endmodule


