//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 0 1 0 0 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G140), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  AND2_X1   g003(.A1(new_n189), .A2(G227), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n188), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  OR2_X1    g006(.A1(KEYINPUT82), .A2(KEYINPUT3), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G104), .ZN(new_n195));
  AND2_X1   g009(.A1(KEYINPUT82), .A2(KEYINPUT3), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n193), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G101), .ZN(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G107), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(G107), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT82), .A2(KEYINPUT3), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n197), .A2(new_n198), .A3(new_n200), .A4(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n195), .A2(new_n200), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G101), .ZN(new_n206));
  AND2_X1   g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n208), .B1(new_n210), .B2(KEYINPUT1), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n209), .A2(KEYINPUT66), .A3(G143), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT66), .B1(new_n209), .B2(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(new_n210), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n211), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n208), .A2(KEYINPUT1), .ZN(new_n216));
  INV_X1    g030(.A(G143), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G146), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n216), .A2(new_n210), .A3(new_n218), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n207), .B(KEYINPUT10), .C1(new_n215), .C2(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n200), .B1(new_n193), .B2(new_n195), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT82), .A2(KEYINPUT3), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n202), .B1(new_n201), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(G101), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(KEYINPUT4), .A3(new_n204), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n226), .B1(new_n217), .B2(G146), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n217), .A2(G146), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n212), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT64), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n230), .B1(KEYINPUT0), .B2(G128), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT0), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(new_n208), .A3(KEYINPUT64), .ZN(new_n233));
  NAND2_X1  g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT65), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(KEYINPUT0), .A3(G128), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n231), .A2(new_n233), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(KEYINPUT0), .A2(G128), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n210), .A2(new_n218), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT67), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n210), .A2(new_n218), .A3(new_n239), .A4(new_n242), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n229), .A2(new_n238), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n245), .B(G101), .C1(new_n221), .C2(new_n223), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n225), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT11), .ZN(new_n248));
  INV_X1    g062(.A(G134), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n248), .B1(new_n249), .B2(G137), .ZN(new_n250));
  INV_X1    g064(.A(G137), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(KEYINPUT11), .A3(G134), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n249), .A2(G137), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G131), .ZN(new_n255));
  INV_X1    g069(.A(G131), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n250), .A2(new_n252), .A3(new_n256), .A4(new_n253), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n210), .A2(new_n218), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(new_n211), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n204), .B(new_n206), .C1(new_n261), .C2(new_n219), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT10), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n220), .A2(new_n247), .A3(new_n259), .A4(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n204), .A2(new_n206), .ZN(new_n266));
  INV_X1    g080(.A(new_n211), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n219), .B1(new_n229), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n262), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT12), .B1(new_n270), .B2(new_n258), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT12), .ZN(new_n272));
  AOI211_X1 g086(.A(new_n272), .B(new_n259), .C1(new_n269), .C2(new_n262), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n265), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT83), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT83), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n265), .B(new_n276), .C1(new_n271), .C2(new_n273), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n192), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n220), .A2(new_n247), .A3(new_n264), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n279), .A2(new_n258), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n265), .A2(new_n192), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n187), .B1(new_n278), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G469), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT84), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT84), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n283), .A2(new_n286), .A3(G469), .ZN(new_n287));
  INV_X1    g101(.A(new_n265), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n191), .B1(new_n280), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n270), .A2(new_n258), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n272), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n270), .A2(KEYINPUT12), .A3(new_n258), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(new_n192), .A3(new_n265), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G469), .ZN(new_n296));
  XOR2_X1   g110(.A(KEYINPUT74), .B(G902), .Z(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n285), .A2(new_n287), .A3(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT9), .B(G234), .ZN(new_n300));
  OAI21_X1  g114(.A(G221), .B1(new_n300), .B2(G902), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n301), .B(KEYINPUT81), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(G214), .B1(G237), .B2(G902), .ZN(new_n304));
  INV_X1    g118(.A(G119), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G116), .ZN(new_n306));
  INV_X1    g120(.A(G116), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G119), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(KEYINPUT2), .A2(G113), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT68), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT68), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(KEYINPUT2), .A3(G113), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(KEYINPUT2), .A2(G113), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n309), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT2), .ZN(new_n317));
  INV_X1    g131(.A(G113), .ZN(new_n318));
  AOI22_X1  g132(.A1(new_n311), .A2(new_n313), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n309), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n225), .A2(new_n322), .A3(new_n246), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT85), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n307), .A2(G119), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT5), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n318), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n306), .A2(new_n308), .A3(KEYINPUT5), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n321), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n324), .B1(new_n266), .B2(new_n330), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n319), .A2(new_n320), .B1(new_n327), .B2(new_n328), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n332), .A2(KEYINPUT85), .A3(new_n204), .A4(new_n206), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n323), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(G110), .B(G122), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n323), .A2(new_n331), .A3(new_n335), .A4(new_n333), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(KEYINPUT6), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT6), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n334), .A2(new_n340), .A3(new_n336), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n238), .A2(new_n229), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n241), .A2(new_n243), .ZN(new_n343));
  INV_X1    g157(.A(G125), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT78), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT78), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G125), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n342), .A2(new_n343), .A3(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n349), .B1(new_n268), .B2(new_n348), .ZN(new_n350));
  INV_X1    g164(.A(G224), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n351), .A2(G953), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n350), .B(new_n353), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n339), .A2(new_n341), .A3(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(G210), .B1(G237), .B2(G902), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n353), .A2(KEYINPUT7), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n349), .B(new_n358), .C1(new_n268), .C2(new_n348), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT86), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n353), .A2(KEYINPUT87), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT7), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT87), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n362), .B1(new_n352), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n350), .A2(new_n361), .A3(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n335), .B(KEYINPUT8), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n207), .A2(new_n332), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n266), .A2(new_n330), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OR2_X1    g183(.A1(new_n268), .A2(new_n348), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT86), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n370), .A2(new_n371), .A3(new_n349), .A4(new_n358), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n360), .A2(new_n365), .A3(new_n369), .A4(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n338), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n187), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n355), .A2(new_n357), .A3(new_n375), .ZN(new_n376));
  AND4_X1   g190(.A1(new_n372), .A2(new_n360), .A3(new_n365), .A4(new_n369), .ZN(new_n377));
  AOI21_X1  g191(.A(G902), .B1(new_n377), .B2(new_n338), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n339), .A2(new_n341), .A3(new_n354), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n356), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n304), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT90), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n345), .A2(new_n347), .A3(G140), .ZN(new_n383));
  INV_X1    g197(.A(G140), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G125), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT77), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT77), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n384), .A3(G125), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n383), .A2(KEYINPUT16), .A3(new_n386), .A4(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT16), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n348), .A2(new_n390), .A3(new_n384), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n389), .A2(G146), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(G146), .B1(new_n389), .B2(new_n391), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n382), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n389), .A2(new_n391), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n209), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(KEYINPUT90), .A3(new_n392), .ZN(new_n398));
  NOR2_X1   g212(.A1(G237), .A2(G953), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n399), .A2(G143), .A3(G214), .ZN(new_n400));
  AOI21_X1  g214(.A(G143), .B1(new_n399), .B2(G214), .ZN(new_n401));
  OAI21_X1  g215(.A(G131), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT17), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n399), .A2(G214), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n217), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n399), .A2(G143), .A3(G214), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(new_n256), .A3(new_n407), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n402), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n404), .B1(new_n409), .B2(new_n403), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n395), .A2(new_n398), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n344), .A2(G140), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n385), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(G146), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n383), .A2(new_n386), .A3(new_n388), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n414), .B1(new_n415), .B2(G146), .ZN(new_n416));
  NAND2_X1  g230(.A1(KEYINPUT18), .A2(G131), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n418), .B1(new_n400), .B2(new_n401), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n406), .A2(new_n407), .A3(new_n417), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OR2_X1    g235(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  XOR2_X1   g236(.A(G113), .B(G122), .Z(new_n423));
  XOR2_X1   g237(.A(KEYINPUT88), .B(G104), .Z(new_n424));
  XOR2_X1   g238(.A(new_n423), .B(new_n424), .Z(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n411), .A2(new_n422), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n426), .B1(new_n411), .B2(new_n422), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n187), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G475), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT89), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n416), .A2(new_n421), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n402), .A2(new_n408), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n392), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n413), .A2(KEYINPUT19), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n436), .B1(new_n415), .B2(KEYINPUT19), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n209), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n433), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n432), .B1(new_n439), .B2(new_n426), .ZN(new_n440));
  INV_X1    g254(.A(new_n438), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n392), .A2(new_n434), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n422), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(KEYINPUT89), .A3(new_n425), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n427), .A2(new_n440), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n446));
  NOR2_X1   g260(.A1(G475), .A2(G902), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n446), .B1(new_n445), .B2(new_n447), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n431), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G952), .ZN(new_n451));
  AOI211_X1 g265(.A(G953), .B(new_n451), .C1(G234), .C2(G237), .ZN(new_n452));
  AOI211_X1 g266(.A(new_n189), .B(new_n297), .C1(G234), .C2(G237), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(G898), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n297), .ZN(new_n457));
  INV_X1    g271(.A(G122), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT91), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT91), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G122), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n307), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n307), .A2(G122), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n194), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n464), .ZN(new_n466));
  NOR3_X1   g280(.A1(new_n462), .A2(G107), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT92), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT13), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT13), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(KEYINPUT92), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n469), .B(new_n471), .C1(G128), .C2(new_n217), .ZN(new_n472));
  XNOR2_X1  g286(.A(G128), .B(G143), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n472), .A2(G134), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n473), .B1(new_n472), .B2(G134), .ZN(new_n475));
  OAI22_X1  g289(.A1(new_n465), .A2(new_n467), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OR3_X1    g290(.A1(new_n458), .A2(KEYINPUT14), .A3(G116), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n464), .A2(KEYINPUT14), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(G107), .B1(new_n479), .B2(new_n462), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n463), .A2(new_n194), .A3(new_n464), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n473), .B(new_n249), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G217), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n300), .A2(new_n485), .A3(G953), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n476), .A2(new_n483), .A3(new_n486), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n457), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT93), .ZN(new_n491));
  INV_X1    g305(.A(G478), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n492), .A2(KEYINPUT15), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n490), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n476), .A2(new_n483), .A3(new_n486), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n486), .B1(new_n476), .B2(new_n483), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n491), .B(new_n297), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n493), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n495), .A2(KEYINPUT94), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(KEYINPUT94), .B1(new_n495), .B2(new_n499), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n456), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR3_X1   g316(.A1(new_n381), .A2(new_n450), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n299), .A2(new_n303), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT80), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n249), .A2(G137), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n251), .A2(G134), .ZN(new_n507));
  OAI21_X1  g321(.A(G131), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n257), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(KEYINPUT69), .B1(new_n268), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n257), .A2(new_n508), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT69), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n511), .B(new_n512), .C1(new_n215), .C2(new_n219), .ZN(new_n513));
  INV_X1    g327(.A(new_n322), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n258), .A2(new_n342), .A3(new_n343), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n510), .A2(new_n513), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n399), .A2(G210), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT27), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT26), .B(G101), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n519), .B(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT70), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n511), .B1(new_n215), .B2(new_n219), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n515), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT30), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n510), .A2(new_n513), .A3(KEYINPUT30), .A4(new_n515), .ZN(new_n529));
  AND4_X1   g343(.A1(new_n524), .A2(new_n528), .A3(new_n529), .A4(new_n322), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n514), .B1(new_n526), .B2(new_n527), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n524), .B1(new_n531), .B2(new_n529), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n523), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT31), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT28), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n535), .B1(new_n526), .B2(new_n322), .ZN(new_n536));
  XOR2_X1   g350(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n537));
  NAND2_X1  g351(.A1(new_n526), .A2(new_n322), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n537), .B1(new_n538), .B2(new_n516), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n536), .B1(new_n539), .B2(KEYINPUT72), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT72), .ZN(new_n541));
  AOI211_X1 g355(.A(new_n541), .B(new_n537), .C1(new_n538), .C2(new_n516), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n522), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT31), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n544), .B(new_n523), .C1(new_n530), .C2(new_n532), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n534), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(G472), .A2(G902), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT32), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT32), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n546), .A2(new_n550), .A3(new_n547), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT29), .ZN(new_n552));
  INV_X1    g366(.A(new_n536), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n538), .A2(new_n516), .ZN(new_n554));
  INV_X1    g368(.A(new_n537), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n553), .B1(new_n556), .B2(new_n541), .ZN(new_n557));
  INV_X1    g371(.A(new_n542), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n522), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n531), .A2(new_n529), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT70), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n531), .A2(new_n524), .A3(new_n529), .ZN(new_n562));
  AOI211_X1 g376(.A(new_n517), .B(new_n521), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n552), .B1(new_n559), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n322), .B1(new_n258), .B2(new_n244), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT73), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n566), .A2(new_n567), .A3(new_n510), .A4(new_n513), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n510), .A2(new_n513), .A3(new_n515), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n565), .A2(new_n568), .B1(new_n322), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n536), .B1(new_n570), .B2(new_n535), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n522), .A2(new_n552), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n297), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n564), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n549), .A2(new_n551), .B1(new_n576), .B2(G472), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n485), .B1(new_n297), .B2(G234), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT22), .B(G137), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n580), .B(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT75), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n584), .B1(new_n305), .B2(G128), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n208), .A2(KEYINPUT75), .A3(G119), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n305), .A2(G128), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT24), .B(G110), .ZN(new_n589));
  OR2_X1    g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT23), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n591), .B1(new_n305), .B2(G128), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n208), .A2(KEYINPUT23), .A3(G119), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n587), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT76), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n594), .A2(new_n595), .A3(G110), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n595), .B1(new_n594), .B2(G110), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n590), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n598), .B1(new_n397), .B2(new_n392), .ZN(new_n599));
  OR2_X1    g413(.A1(new_n594), .A2(G110), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n588), .A2(new_n589), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n414), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n602), .A2(new_n392), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n583), .B1(new_n599), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n392), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n393), .A2(new_n394), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n605), .B(new_n582), .C1(new_n606), .C2(new_n598), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT25), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n457), .B1(KEYINPUT79), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n604), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n608), .A2(KEYINPUT79), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n579), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n611), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n604), .A2(new_n607), .A3(new_n613), .A4(new_n609), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n578), .A2(G902), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n604), .A2(new_n616), .A3(new_n607), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n505), .B1(new_n577), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n517), .B1(new_n561), .B2(new_n562), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n522), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n521), .B1(new_n540), .B2(new_n542), .ZN(new_n622));
  AOI21_X1  g436(.A(KEYINPUT29), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(G472), .B1(new_n623), .B2(new_n574), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n546), .A2(new_n550), .A3(new_n547), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n550), .B1(new_n546), .B2(new_n547), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n618), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(KEYINPUT80), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n504), .B1(new_n619), .B2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(new_n198), .ZN(G3));
  AOI211_X1 g445(.A(G469), .B(new_n457), .C1(new_n289), .C2(new_n294), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n632), .B1(new_n284), .B2(KEYINPUT84), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n302), .B1(new_n633), .B2(new_n287), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n357), .B1(new_n355), .B2(new_n375), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n378), .A2(new_n356), .A3(new_n379), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n637), .A2(new_n304), .A3(new_n456), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n490), .A2(new_n492), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n488), .A2(new_n489), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT33), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT33), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n488), .A2(new_n642), .A3(new_n489), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n457), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n639), .B1(new_n644), .B2(new_n492), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(KEYINPUT95), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT95), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n647), .B(new_n639), .C1(new_n644), .C2(new_n492), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n450), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n638), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n548), .ZN(new_n651));
  INV_X1    g465(.A(G472), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n546), .B2(new_n297), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n651), .A2(new_n653), .A3(new_n618), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n634), .A2(new_n650), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT34), .B(G104), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT97), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT96), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n655), .B(new_n658), .ZN(G6));
  INV_X1    g473(.A(new_n449), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n500), .A2(new_n501), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n662), .A2(new_n663), .A3(new_n431), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n638), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n634), .A2(new_n654), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT35), .B(G107), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  NOR2_X1   g482(.A1(new_n583), .A2(KEYINPUT36), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n670), .B1(new_n599), .B2(new_n603), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n605), .B(new_n669), .C1(new_n606), .C2(new_n598), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n671), .A2(new_n616), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT98), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n671), .A2(KEYINPUT98), .A3(new_n616), .A4(new_n672), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(new_n614), .B2(new_n612), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT99), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n675), .A2(new_n676), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n615), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT99), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n684), .A2(new_n651), .A3(new_n653), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n634), .A2(new_n685), .A3(new_n503), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT37), .B(G110), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G12));
  AND3_X1   g502(.A1(new_n680), .A2(new_n615), .A3(KEYINPUT99), .ZN(new_n689));
  AOI21_X1  g503(.A(KEYINPUT99), .B1(new_n680), .B2(new_n615), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n381), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(G900), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n452), .B1(new_n453), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n664), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n634), .A2(new_n627), .A3(new_n691), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G128), .ZN(G30));
  XOR2_X1   g510(.A(new_n693), .B(KEYINPUT39), .Z(new_n697));
  NAND2_X1  g511(.A1(new_n634), .A2(new_n697), .ZN(new_n698));
  OR2_X1    g512(.A1(new_n698), .A2(KEYINPUT40), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(KEYINPUT40), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n637), .B(KEYINPUT38), .Z(new_n701));
  OR2_X1    g515(.A1(new_n620), .A2(new_n522), .ZN(new_n702));
  AOI21_X1  g516(.A(G902), .B1(new_n570), .B2(new_n522), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n652), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n704), .B1(new_n549), .B2(new_n551), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n450), .A2(new_n678), .A3(new_n663), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n304), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n701), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n699), .A2(new_n700), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G143), .ZN(G45));
  INV_X1    g524(.A(new_n693), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n450), .A2(new_n646), .A3(new_n648), .A4(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n634), .A2(new_n627), .A3(new_n691), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G146), .ZN(G48));
  NAND2_X1  g529(.A1(new_n295), .A2(new_n297), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(G469), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n303), .A3(new_n298), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n627), .A2(new_n650), .A3(new_n628), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT41), .B(G113), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT100), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n720), .B(new_n722), .ZN(G15));
  NAND4_X1  g537(.A1(new_n627), .A2(new_n665), .A3(new_n628), .A4(new_n719), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G116), .ZN(G18));
  NOR2_X1   g539(.A1(new_n502), .A2(new_n450), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n627), .A2(new_n691), .A3(new_n726), .A4(new_n719), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  INV_X1    g542(.A(new_n547), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n534), .A2(new_n545), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT101), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n571), .A2(new_n731), .ZN(new_n732));
  OAI211_X1 g546(.A(KEYINPUT101), .B(new_n536), .C1(new_n570), .C2(new_n535), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(new_n522), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n729), .B1(new_n730), .B2(new_n734), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n735), .A2(new_n653), .A3(new_n618), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n450), .A2(new_n663), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n381), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n718), .A2(new_n455), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n736), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G122), .ZN(G24));
  NOR3_X1   g555(.A1(new_n735), .A2(new_n653), .A3(new_n678), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n646), .A2(new_n648), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT102), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n743), .A2(new_n744), .A3(new_n450), .A4(new_n711), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n718), .A2(new_n381), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n712), .A2(KEYINPUT102), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n742), .A2(new_n745), .A3(new_n746), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G125), .ZN(G27));
  NOR2_X1   g563(.A1(new_n577), .A2(new_n618), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n712), .B(new_n744), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n632), .B1(new_n283), .B2(G469), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n635), .A2(new_n304), .A3(new_n636), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n752), .A2(new_n302), .A3(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n750), .A2(new_n751), .A3(KEYINPUT42), .A4(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT42), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n754), .A2(new_n627), .A3(new_n628), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n745), .A2(new_n747), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G131), .ZN(G33));
  NAND3_X1  g575(.A1(new_n750), .A2(new_n694), .A3(new_n754), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G134), .ZN(G36));
  INV_X1    g577(.A(KEYINPUT104), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n278), .A2(new_n282), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n765), .A2(KEYINPUT45), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(KEYINPUT45), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(G469), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(G469), .A2(G902), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(KEYINPUT46), .A3(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(KEYINPUT103), .A3(new_n298), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n768), .A2(new_n769), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n771), .B1(KEYINPUT46), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT103), .B1(new_n770), .B2(new_n298), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n303), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n697), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n764), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n773), .A2(new_n774), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n778), .A2(KEYINPUT104), .A3(new_n303), .A4(new_n697), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n681), .B1(new_n651), .B2(new_n653), .ZN(new_n780));
  XOR2_X1   g594(.A(new_n780), .B(KEYINPUT107), .Z(new_n781));
  INV_X1    g595(.A(new_n450), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n743), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT106), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n783), .A2(KEYINPUT106), .A3(new_n784), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT43), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n786), .B1(new_n787), .B2(new_n783), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n781), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT44), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n753), .B1(new_n789), .B2(new_n790), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n777), .A2(new_n779), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G137), .ZN(G39));
  INV_X1    g608(.A(KEYINPUT47), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n775), .B(new_n795), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n712), .A2(new_n628), .A3(new_n753), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n577), .A3(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  INV_X1    g613(.A(new_n655), .ZN(new_n800));
  OAI21_X1  g614(.A(KEYINPUT108), .B1(new_n630), .B2(new_n800), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n299), .A2(new_n303), .A3(new_n503), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n627), .A2(KEYINPUT80), .A3(new_n628), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT80), .B1(new_n627), .B2(new_n628), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT108), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(new_n806), .A3(new_n655), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n495), .A2(new_n499), .A3(KEYINPUT109), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n495), .A2(new_n499), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT109), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n782), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n638), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n634), .A2(new_n654), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n686), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT110), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n686), .A2(new_n814), .A3(KEYINPUT110), .ZN(new_n818));
  AOI22_X1  g632(.A1(new_n801), .A2(new_n807), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n695), .A2(new_n714), .A3(new_n748), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT111), .ZN(new_n822));
  INV_X1    g636(.A(new_n304), .ZN(new_n823));
  AOI211_X1 g637(.A(new_n823), .B(new_n693), .C1(new_n635), .C2(new_n636), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n276), .B1(new_n293), .B2(new_n265), .ZN(new_n825));
  INV_X1    g639(.A(new_n277), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n191), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n282), .ZN(new_n828));
  AOI21_X1  g642(.A(G902), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n298), .B1(new_n829), .B2(new_n296), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n706), .A2(new_n824), .A3(new_n830), .A4(new_n303), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n822), .B1(new_n831), .B2(new_n705), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n450), .A2(new_n678), .A3(new_n663), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n833), .A2(new_n381), .A3(new_n693), .ZN(new_n834));
  INV_X1    g648(.A(new_n704), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n835), .B1(new_n625), .B2(new_n626), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n752), .A2(new_n302), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n834), .A2(new_n836), .A3(KEYINPUT111), .A4(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n832), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n820), .B1(new_n821), .B2(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n299), .A2(new_n303), .A3(new_n691), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n841), .B(new_n627), .C1(new_n694), .C2(new_n713), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n832), .A2(new_n838), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(KEYINPUT52), .A3(new_n748), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n720), .A2(new_n724), .A3(new_n740), .A4(new_n727), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n693), .B1(new_n811), .B2(new_n808), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n431), .A3(new_n662), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n684), .A2(new_n848), .A3(new_n753), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n634), .A2(new_n849), .A3(new_n627), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n742), .A2(new_n745), .A3(new_n754), .A4(new_n747), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AND4_X1   g666(.A1(new_n760), .A2(new_n846), .A3(new_n762), .A4(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n819), .A2(new_n845), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT112), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n840), .A2(new_n857), .A3(new_n844), .ZN(new_n858));
  OAI211_X1 g672(.A(KEYINPUT112), .B(new_n820), .C1(new_n821), .C2(new_n839), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n819), .A2(KEYINPUT53), .A3(new_n853), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n856), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  XOR2_X1   g676(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n863));
  OR3_X1    g677(.A1(new_n862), .A2(KEYINPUT115), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT113), .ZN(new_n865));
  OR3_X1    g679(.A1(new_n854), .A2(new_n865), .A3(new_n855), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n819), .A2(new_n853), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n855), .B1(new_n860), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n865), .B1(new_n854), .B2(new_n855), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n866), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT54), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT115), .B1(new_n862), .B2(new_n863), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n864), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n452), .B(new_n736), .C1(new_n788), .C2(new_n785), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n753), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n717), .A2(new_n298), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n876), .A2(new_n303), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n875), .B1(new_n796), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n719), .A2(new_n823), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n879), .A2(KEYINPUT116), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(KEYINPUT116), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n880), .A2(new_n701), .A3(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n874), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT50), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT117), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n718), .A2(new_n753), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n452), .B(new_n886), .C1(new_n788), .C2(new_n785), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  AND4_X1   g702(.A1(new_n628), .A2(new_n705), .A3(new_n452), .A4(new_n886), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n743), .A2(new_n450), .ZN(new_n890));
  AOI22_X1  g704(.A1(new_n888), .A2(new_n742), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n884), .A2(new_n885), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n885), .B1(new_n884), .B2(new_n891), .ZN(new_n893));
  OAI211_X1 g707(.A(KEYINPUT51), .B(new_n878), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n649), .ZN(new_n895));
  AOI211_X1 g709(.A(new_n451), .B(G953), .C1(new_n889), .C2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n746), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n887), .A2(new_n577), .A3(new_n618), .ZN(new_n898));
  OAI221_X1 g712(.A(new_n896), .B1(new_n897), .B2(new_n874), .C1(new_n898), .C2(KEYINPUT48), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(KEYINPUT48), .B2(new_n898), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n878), .A2(new_n884), .A3(new_n891), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n894), .B(new_n900), .C1(new_n901), .C2(KEYINPUT51), .ZN(new_n902));
  OAI22_X1  g716(.A1(new_n873), .A2(new_n902), .B1(G952), .B2(G953), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n618), .A2(new_n302), .A3(new_n823), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n904), .B1(new_n876), .B2(KEYINPUT49), .ZN(new_n905));
  AOI211_X1 g719(.A(new_n783), .B(new_n905), .C1(KEYINPUT49), .C2(new_n876), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n705), .A3(new_n701), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n903), .A2(new_n907), .ZN(G75));
  NOR2_X1   g722(.A1(new_n189), .A2(G952), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n862), .A2(new_n457), .A3(new_n357), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n339), .A2(new_n341), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(new_n354), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT55), .ZN(new_n913));
  XNOR2_X1  g727(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n909), .B1(new_n910), .B2(new_n915), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n819), .A2(KEYINPUT53), .A3(new_n853), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n858), .A2(new_n859), .ZN(new_n918));
  AOI22_X1  g732(.A1(new_n917), .A2(new_n918), .B1(new_n855), .B2(new_n854), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n919), .A2(new_n297), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT56), .B1(new_n920), .B2(new_n357), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n916), .B1(new_n921), .B2(new_n913), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT119), .ZN(G51));
  XNOR2_X1  g737(.A(new_n862), .B(new_n863), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n769), .B(KEYINPUT57), .Z(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n295), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n768), .B(KEYINPUT120), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n920), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n909), .B1(new_n927), .B2(new_n929), .ZN(G54));
  NAND3_X1  g744(.A1(new_n920), .A2(KEYINPUT58), .A3(G475), .ZN(new_n931));
  INV_X1    g745(.A(new_n445), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n933), .A2(new_n934), .A3(new_n909), .ZN(G60));
  AND2_X1   g749(.A1(new_n641), .A2(new_n643), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(G478), .A2(G902), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT59), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n937), .B1(new_n873), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n924), .A2(new_n937), .A3(new_n939), .ZN(new_n941));
  INV_X1    g755(.A(new_n909), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n940), .A2(new_n943), .ZN(G63));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n945), .A2(KEYINPUT123), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT122), .ZN(new_n947));
  XNOR2_X1  g761(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n485), .A2(new_n187), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n947), .B1(new_n919), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n604), .A2(new_n607), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n854), .A2(new_n855), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n861), .A2(new_n860), .ZN(new_n955));
  OAI211_X1 g769(.A(KEYINPUT122), .B(new_n950), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n952), .A2(new_n953), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n909), .B1(KEYINPUT123), .B2(new_n945), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n671), .A2(new_n672), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n952), .B2(new_n956), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n946), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n952), .A2(new_n956), .ZN(new_n963));
  INV_X1    g777(.A(new_n960), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n946), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n965), .A2(new_n966), .A3(new_n957), .A4(new_n958), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n962), .A2(new_n967), .ZN(G66));
  OAI21_X1  g782(.A(G953), .B1(new_n454), .B2(new_n351), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n819), .A2(new_n846), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n969), .B1(new_n970), .B2(G953), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n911), .B1(G898), .B2(new_n189), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT124), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n971), .B(new_n973), .ZN(G69));
  AOI21_X1  g788(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n753), .B1(new_n812), .B2(new_n649), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n634), .A2(new_n976), .A3(new_n697), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n619), .B2(new_n629), .ZN(new_n978));
  INV_X1    g792(.A(new_n821), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n979), .A2(KEYINPUT126), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(KEYINPUT126), .ZN(new_n981));
  OR2_X1    g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n709), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT62), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n982), .A2(KEYINPUT62), .A3(new_n709), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n978), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n798), .A2(new_n793), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(G953), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n528), .A2(new_n529), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT125), .Z(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(new_n437), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n990), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n779), .A2(new_n777), .A3(new_n750), .A4(new_n738), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n996), .A2(new_n982), .A3(new_n760), .A4(new_n762), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n189), .B1(new_n988), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n692), .A2(G953), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT127), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n993), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n975), .B1(new_n995), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1001), .ZN(new_n1003));
  INV_X1    g817(.A(new_n975), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n1003), .B(new_n1004), .C1(new_n990), .C2(new_n994), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1002), .A2(new_n1005), .ZN(G72));
  NAND2_X1  g820(.A1(G472), .A2(G902), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT63), .Z(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n988), .A2(new_n997), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1009), .B1(new_n1010), .B2(new_n970), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n942), .B1(new_n1011), .B2(new_n621), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n987), .A2(new_n970), .A3(new_n989), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n702), .B1(new_n1013), .B2(new_n1008), .ZN(new_n1014));
  AND4_X1   g828(.A1(new_n621), .A2(new_n870), .A3(new_n702), .A4(new_n1008), .ZN(new_n1015));
  NOR3_X1   g829(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .ZN(G57));
endmodule


