//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 0 1 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969;
  XNOR2_X1  g000(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n187));
  XNOR2_X1  g001(.A(G113), .B(G122), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  INV_X1    g006(.A(G140), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G125), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT73), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n192), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n191), .A2(KEYINPUT73), .A3(G140), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT16), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n194), .A2(KEYINPUT16), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n199), .A2(G146), .A3(new_n201), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n192), .A2(new_n194), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT19), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n205), .B1(new_n198), .B2(new_n204), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n202), .B1(G146), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT89), .ZN(new_n208));
  OR2_X1    g022(.A1(new_n206), .A2(G146), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT89), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(new_n202), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT88), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G143), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT88), .ZN(new_n215));
  NOR2_X1   g029(.A1(G237), .A2(G953), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n213), .A2(new_n215), .A3(G214), .A4(new_n216), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n216), .A2(G214), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n217), .B1(new_n218), .B2(new_n213), .ZN(new_n219));
  INV_X1    g033(.A(G131), .ZN(new_n220));
  OR2_X1    g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n220), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n208), .A2(new_n211), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n219), .A2(new_n220), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT18), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT18), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n219), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G146), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n203), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n230), .B1(new_n198), .B2(new_n229), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n226), .A2(new_n228), .A3(new_n231), .A4(new_n222), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n190), .B1(new_n224), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT17), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n221), .A2(new_n234), .A3(new_n222), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT16), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n236), .B1(new_n196), .B2(new_n197), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n229), .B1(new_n237), .B2(new_n200), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n225), .A2(KEYINPUT17), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n235), .A2(new_n238), .A3(new_n202), .A4(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(new_n190), .A3(new_n232), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n233), .A2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(G475), .A2(G902), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n187), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(KEYINPUT90), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT90), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT20), .B1(new_n244), .B2(new_n248), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n247), .B(new_n249), .C1(new_n233), .C2(new_n242), .ZN(new_n250));
  INV_X1    g064(.A(G902), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n190), .B1(new_n240), .B2(new_n232), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n251), .B1(new_n242), .B2(new_n252), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n246), .A2(new_n250), .B1(G475), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G116), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(KEYINPUT14), .A3(G122), .ZN(new_n256));
  XOR2_X1   g070(.A(G116), .B(G122), .Z(new_n257));
  OAI211_X1 g071(.A(G107), .B(new_n256), .C1(new_n257), .C2(KEYINPUT14), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT93), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n258), .B(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n214), .A2(G128), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n214), .A2(G128), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G134), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  OR2_X1    g080(.A1(new_n257), .A2(G107), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n260), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT13), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n261), .B1(new_n263), .B2(new_n269), .ZN(new_n270));
  OR2_X1    g084(.A1(new_n270), .A2(KEYINPUT91), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n270), .B(KEYINPUT91), .C1(new_n269), .C2(new_n261), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(G134), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT92), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n257), .A2(G107), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n267), .A2(new_n276), .B1(new_n265), .B2(new_n264), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n271), .A2(new_n272), .A3(KEYINPUT92), .A4(G134), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n275), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  XOR2_X1   g093(.A(KEYINPUT9), .B(G234), .Z(new_n280));
  INV_X1    g094(.A(G953), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(G217), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n268), .A2(new_n279), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n283), .B1(new_n268), .B2(new_n279), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n251), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G478), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n287), .A2(KEYINPUT15), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n288), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n251), .B(new_n290), .C1(new_n284), .C2(new_n285), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n281), .A2(G952), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n292), .B1(G234), .B2(G237), .ZN(new_n293));
  XOR2_X1   g107(.A(KEYINPUT21), .B(G898), .Z(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  AOI211_X1 g109(.A(new_n251), .B(new_n281), .C1(G234), .C2(G237), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n293), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n289), .A2(new_n291), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(KEYINPUT94), .B1(new_n254), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n253), .A2(G475), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n223), .B1(new_n207), .B2(KEYINPUT89), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n210), .B1(new_n209), .B2(new_n202), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n232), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n190), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n245), .B1(new_n306), .B2(new_n241), .ZN(new_n307));
  INV_X1    g121(.A(new_n187), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n250), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AND4_X1   g123(.A1(KEYINPUT94), .A2(new_n299), .A3(new_n301), .A4(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n300), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT3), .ZN(new_n313));
  INV_X1    g127(.A(G107), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n314), .A3(G104), .ZN(new_n315));
  INV_X1    g129(.A(G101), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n189), .A2(G107), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n312), .A2(new_n315), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT78), .ZN(new_n319));
  OR2_X1    g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n319), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n314), .A2(G104), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n320), .A2(new_n321), .B1(G101), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G119), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G116), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n255), .A2(G119), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT2), .B(G113), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT65), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G113), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT2), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT2), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G113), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(G116), .B(G119), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT65), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n330), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n336), .A2(KEYINPUT5), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n340), .B(G113), .C1(KEYINPUT5), .C2(new_n326), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n324), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT4), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n312), .A2(new_n315), .A3(new_n317), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n343), .B1(new_n344), .B2(G101), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n318), .A2(new_n319), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n318), .A2(new_n319), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT79), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n344), .A2(new_n343), .A3(G101), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n318), .B(new_n319), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(KEYINPUT79), .A3(new_n345), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n350), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n335), .A2(new_n336), .ZN(new_n355));
  AOI211_X1 g169(.A(KEYINPUT66), .B(new_n355), .C1(new_n338), .C2(new_n330), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT66), .ZN(new_n357));
  INV_X1    g171(.A(new_n355), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n357), .B1(new_n339), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n342), .B1(new_n354), .B2(new_n360), .ZN(new_n361));
  XOR2_X1   g175(.A(G110), .B(G122), .Z(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n362), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n364), .B(new_n342), .C1(new_n354), .C2(new_n360), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n363), .A2(KEYINPUT6), .A3(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(G143), .B(G146), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT0), .ZN(new_n368));
  INV_X1    g182(.A(G128), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n214), .A2(G146), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n229), .A2(G143), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n368), .A2(new_n369), .ZN(new_n373));
  NOR2_X1   g187(.A1(KEYINPUT0), .A2(G128), .ZN(new_n374));
  OAI22_X1  g188(.A1(new_n371), .A2(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G125), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT1), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G128), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n229), .A2(new_n263), .B1(new_n372), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n379), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n367), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n191), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n377), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G224), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(G953), .ZN(new_n387));
  XOR2_X1   g201(.A(new_n385), .B(new_n387), .Z(new_n388));
  INV_X1    g202(.A(KEYINPUT6), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n361), .A2(new_n389), .A3(new_n362), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n366), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  XOR2_X1   g205(.A(new_n362), .B(KEYINPUT8), .Z(new_n392));
  AND3_X1   g206(.A1(new_n324), .A2(new_n339), .A3(new_n341), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n324), .B1(new_n339), .B2(new_n341), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n385), .B(KEYINPUT7), .C1(new_n386), .C2(G953), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT7), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n377), .B(new_n384), .C1(new_n397), .C2(new_n387), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT86), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n398), .B(new_n399), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n365), .A2(new_n395), .A3(new_n396), .A4(new_n400), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n401), .A2(new_n251), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n391), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(G210), .B1(G237), .B2(G902), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n391), .A2(new_n402), .A3(new_n404), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(G214), .B1(G237), .B2(G902), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(KEYINPUT85), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n311), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G221), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n413), .B1(new_n280), .B2(new_n251), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n323), .A2(G101), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n382), .A2(KEYINPUT80), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT80), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n367), .A2(new_n418), .A3(new_n381), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(new_n380), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n352), .A2(new_n416), .A3(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(new_n383), .B2(new_n324), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT81), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT11), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n424), .B1(new_n265), .B2(G137), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n265), .A2(G137), .ZN(new_n426));
  INV_X1    g240(.A(G137), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(KEYINPUT11), .A3(G134), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n425), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(G131), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n425), .A2(new_n428), .A3(new_n220), .A4(new_n426), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n422), .A2(new_n423), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT12), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n350), .A2(new_n353), .A3(new_n376), .A4(new_n351), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT10), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n436), .B1(new_n380), .B2(new_n382), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n421), .A2(new_n436), .B1(new_n324), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n432), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n435), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT12), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n422), .A2(new_n423), .A3(new_n441), .A4(new_n432), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n434), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  OR2_X1    g257(.A1(new_n443), .A2(KEYINPUT82), .ZN(new_n444));
  XNOR2_X1  g258(.A(G110), .B(G140), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n281), .A2(G227), .ZN(new_n446));
  XOR2_X1   g260(.A(new_n445), .B(new_n446), .Z(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(new_n443), .B2(KEYINPUT82), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n435), .A2(new_n438), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT83), .B1(new_n449), .B2(new_n432), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT83), .ZN(new_n451));
  AOI211_X1 g265(.A(new_n451), .B(new_n439), .C1(new_n435), .C2(new_n438), .ZN(new_n452));
  OR2_X1    g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n440), .A2(new_n447), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n444), .A2(new_n448), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(G469), .B1(new_n455), .B2(G902), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT84), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n440), .B1(new_n450), .B2(new_n452), .ZN(new_n458));
  INV_X1    g272(.A(new_n447), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n434), .A2(new_n442), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n454), .ZN(new_n462));
  AOI21_X1  g276(.A(G902), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G469), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n457), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n458), .A2(new_n459), .B1(new_n461), .B2(new_n454), .ZN(new_n466));
  NOR4_X1   g280(.A1(new_n466), .A2(KEYINPUT84), .A3(G469), .A4(G902), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n456), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n412), .A2(new_n415), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT95), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT70), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(G101), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n216), .A2(G210), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n473), .B(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n426), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n265), .A2(G137), .ZN(new_n477));
  OAI21_X1  g291(.A(G131), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n383), .A2(new_n431), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n432), .A2(new_n376), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT67), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n432), .A2(KEYINPUT67), .A3(new_n376), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n480), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n339), .A2(new_n358), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT66), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n339), .A2(new_n357), .A3(new_n358), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(KEYINPUT68), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT68), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n490), .B1(new_n356), .B2(new_n359), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n485), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT69), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n485), .A2(new_n489), .A3(new_n491), .A4(KEYINPUT69), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n481), .A2(KEYINPUT64), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT64), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n498), .B1(new_n432), .B2(new_n376), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n479), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n360), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT28), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT28), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n489), .A2(new_n491), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n481), .A2(new_n479), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n475), .B1(new_n504), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT30), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n510), .B(new_n479), .C1(new_n497), .C2(new_n499), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n510), .B2(new_n485), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n501), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n496), .A2(new_n475), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT31), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT31), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n496), .A2(new_n516), .A3(new_n475), .A4(new_n513), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n471), .B1(new_n509), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n494), .A2(new_n495), .B1(new_n501), .B2(new_n500), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n508), .B1(new_n520), .B2(new_n505), .ZN(new_n521));
  INV_X1    g335(.A(new_n475), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n523), .A2(KEYINPUT70), .A3(new_n515), .A4(new_n517), .ZN(new_n524));
  NOR2_X1   g338(.A1(G472), .A2(G902), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n519), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT32), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT32), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n519), .A2(new_n524), .A3(new_n528), .A4(new_n525), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n508), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT71), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n496), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n494), .A2(KEYINPUT71), .A3(new_n495), .ZN(new_n534));
  INV_X1    g348(.A(new_n506), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n533), .B(new_n534), .C1(new_n535), .C2(new_n485), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n531), .B1(new_n536), .B2(KEYINPUT28), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(KEYINPUT29), .A3(new_n475), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n504), .A2(new_n508), .A3(new_n475), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n475), .B1(new_n496), .B2(new_n513), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n540), .A2(KEYINPUT29), .ZN(new_n541));
  AOI21_X1  g355(.A(G902), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(G472), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n530), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n460), .A2(new_n462), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n251), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT84), .B1(new_n547), .B2(G469), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n463), .A2(new_n457), .A3(new_n464), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n414), .B1(new_n550), .B2(new_n456), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT95), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n552), .A3(new_n412), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n369), .A2(G119), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT23), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n554), .B1(KEYINPUT72), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n325), .A2(G128), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT72), .B(KEYINPUT23), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n556), .B(new_n557), .C1(new_n558), .C2(new_n554), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n554), .A2(new_n557), .ZN(new_n560));
  XOR2_X1   g374(.A(KEYINPUT24), .B(G110), .Z(new_n561));
  OAI22_X1  g375(.A1(new_n559), .A2(G110), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n202), .A2(new_n562), .A3(new_n230), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n202), .A2(new_n238), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT74), .ZN(new_n565));
  AOI22_X1  g379(.A1(new_n559), .A2(G110), .B1(new_n560), .B2(new_n561), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n565), .B1(new_n564), .B2(new_n566), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n563), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT75), .B(KEYINPUT22), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(G137), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n281), .A2(G221), .A3(G234), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n571), .B(new_n572), .Z(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n563), .B(new_n573), .C1(new_n567), .C2(new_n568), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n251), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT25), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n575), .A2(KEYINPUT25), .A3(new_n251), .A4(new_n576), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(G217), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n582), .B1(G234), .B2(new_n251), .ZN(new_n583));
  AOI21_X1  g397(.A(KEYINPUT76), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT76), .ZN(new_n585));
  INV_X1    g399(.A(new_n583), .ZN(new_n586));
  AOI211_X1 g400(.A(new_n585), .B(new_n586), .C1(new_n579), .C2(new_n580), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n577), .A2(new_n583), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT77), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n584), .A2(new_n587), .A3(new_n589), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT77), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n470), .A2(new_n545), .A3(new_n553), .A4(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G101), .ZN(G3));
  NAND3_X1  g412(.A1(new_n519), .A2(new_n251), .A3(new_n524), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(G472), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n594), .B1(new_n588), .B2(new_n590), .ZN(new_n601));
  NOR4_X1   g415(.A1(new_n584), .A2(new_n587), .A3(KEYINPUT77), .A4(new_n589), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n600), .B(new_n526), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n468), .A2(new_n415), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT96), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n600), .A2(new_n526), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT96), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n606), .A2(new_n607), .A3(new_n596), .A4(new_n551), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n408), .A2(new_n409), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n298), .ZN(new_n611));
  INV_X1    g425(.A(new_n286), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n287), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n287), .A2(new_n251), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  OR2_X1    g429(.A1(new_n284), .A2(new_n285), .ZN(new_n616));
  AOI21_X1  g430(.A(KEYINPUT97), .B1(new_n268), .B2(new_n279), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT33), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n616), .B(new_n619), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n613), .B(new_n615), .C1(new_n620), .C2(new_n287), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n254), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n611), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n609), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT34), .B(G104), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT98), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n625), .B(new_n627), .ZN(G6));
  INV_X1    g442(.A(new_n246), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n243), .A2(new_n245), .A3(new_n187), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n301), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n290), .B1(new_n616), .B2(new_n251), .ZN(new_n632));
  INV_X1    g446(.A(new_n291), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OR2_X1    g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n611), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n609), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT35), .B(G107), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G9));
  NAND2_X1  g453(.A1(new_n581), .A2(new_n583), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n585), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n574), .A2(KEYINPUT36), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n569), .B(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n643), .A2(new_n251), .A3(new_n586), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n581), .A2(KEYINPUT76), .A3(new_n583), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n641), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT99), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT99), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n588), .A2(new_n648), .A3(new_n644), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n470), .A2(new_n553), .A3(new_n606), .A4(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n652), .B(KEYINPUT37), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G110), .ZN(G12));
  AOI21_X1  g468(.A(new_n650), .B1(new_n530), .B2(new_n544), .ZN(new_n655));
  INV_X1    g469(.A(new_n296), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT100), .B(G900), .Z(new_n657));
  OR3_X1    g471(.A1(new_n656), .A2(KEYINPUT101), .A3(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n293), .ZN(new_n659));
  OAI21_X1  g473(.A(KEYINPUT101), .B1(new_n656), .B2(new_n657), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n468), .A2(new_n415), .A3(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n635), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n655), .A2(new_n610), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G128), .ZN(G30));
  XOR2_X1   g479(.A(new_n661), .B(KEYINPUT39), .Z(new_n666));
  OR2_X1    g480(.A1(new_n604), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT104), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT40), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n514), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n536), .B2(new_n522), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n673), .A2(KEYINPUT102), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n251), .B1(new_n673), .B2(KEYINPUT102), .ZN(new_n675));
  OAI21_X1  g489(.A(G472), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n530), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n409), .B1(new_n632), .B2(new_n633), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n254), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n650), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT103), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n678), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT38), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n408), .B(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n683), .B(new_n686), .C1(new_n682), .C2(new_n681), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n671), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT105), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n214), .ZN(G45));
  NOR2_X1   g504(.A1(new_n662), .A2(new_n623), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n655), .A2(new_n610), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G146), .ZN(G48));
  NAND2_X1  g507(.A1(new_n547), .A2(G469), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n550), .A2(new_n415), .A3(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n545), .A2(new_n624), .A3(new_n596), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT41), .B(G113), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G15));
  NAND4_X1  g513(.A1(new_n545), .A2(new_n636), .A3(new_n596), .A4(new_n696), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G116), .ZN(G18));
  INV_X1    g515(.A(new_n311), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n655), .A2(new_n702), .A3(new_n610), .A4(new_n696), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G119), .ZN(G21));
  INV_X1    g518(.A(new_n525), .ZN(new_n705));
  OR2_X1    g519(.A1(new_n537), .A2(new_n475), .ZN(new_n706));
  INV_X1    g520(.A(new_n518), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n600), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n599), .A2(KEYINPUT106), .A3(G472), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n708), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n680), .A2(new_n408), .A3(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n713), .B1(new_n680), .B2(new_n408), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n695), .A2(new_n297), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n712), .A2(new_n593), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G122), .ZN(G24));
  AND4_X1   g535(.A1(new_n415), .A2(new_n550), .A3(new_n610), .A4(new_n694), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n622), .A2(new_n661), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n712), .A2(new_n651), .A3(new_n722), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G125), .ZN(G27));
  INV_X1    g540(.A(new_n409), .ZN(new_n727));
  OAI21_X1  g541(.A(KEYINPUT108), .B1(new_n408), .B2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT108), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n406), .A2(new_n729), .A3(new_n407), .A4(new_n409), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n691), .A2(new_n545), .A3(new_n593), .A4(new_n732), .ZN(new_n733));
  AOI22_X1  g547(.A1(new_n527), .A2(new_n529), .B1(G472), .B2(new_n543), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n601), .A2(new_n602), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n734), .A2(new_n735), .A3(new_n731), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n662), .A2(KEYINPUT42), .A3(new_n623), .ZN(new_n737));
  AOI22_X1  g551(.A1(new_n733), .A2(KEYINPUT42), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G131), .ZN(G33));
  NAND4_X1  g553(.A1(new_n663), .A2(new_n545), .A3(new_n596), .A4(new_n732), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G134), .ZN(G36));
  XOR2_X1   g555(.A(new_n455), .B(KEYINPUT45), .Z(new_n742));
  OAI21_X1  g556(.A(G469), .B1(new_n742), .B2(G902), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(KEYINPUT46), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT46), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n745), .B(G469), .C1(new_n742), .C2(G902), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n744), .A2(new_n550), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n415), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(new_n666), .ZN(new_n749));
  INV_X1    g563(.A(new_n606), .ZN(new_n750));
  INV_X1    g564(.A(new_n254), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n621), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT43), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n750), .A2(new_n651), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT44), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n749), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n731), .B(KEYINPUT109), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(new_n754), .B2(new_n755), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(new_n427), .ZN(G39));
  XNOR2_X1  g575(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n748), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n764));
  AOI22_X1  g578(.A1(new_n747), .A2(new_n415), .B1(KEYINPUT110), .B2(new_n764), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n763), .A2(new_n765), .A3(new_n545), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n766), .A2(new_n735), .A3(new_n724), .A4(new_n732), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G140), .ZN(G42));
  NOR2_X1   g582(.A1(new_n717), .A2(new_n662), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n769), .A2(new_n588), .A3(new_n677), .A4(new_n644), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n725), .A2(new_n664), .A3(new_n770), .A4(new_n692), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT52), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n703), .A2(new_n720), .A3(new_n697), .A4(new_n700), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n408), .A2(new_n410), .A3(new_n298), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n254), .B1(new_n632), .B2(new_n633), .ZN(new_n778));
  OR3_X1    g592(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n777), .B1(new_n776), .B2(new_n778), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n779), .B(new_n780), .C1(new_n623), .C2(new_n776), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n605), .A2(new_n608), .A3(new_n781), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n782), .A2(new_n597), .A3(new_n652), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n775), .A2(new_n783), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n604), .A2(new_n731), .A3(new_n631), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n634), .A2(new_n661), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n655), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n655), .A2(new_n785), .A3(KEYINPUT113), .A4(new_n786), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n604), .A2(new_n731), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n712), .A2(new_n651), .A3(new_n724), .A4(new_n792), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n793), .A2(new_n740), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n791), .A2(new_n794), .A3(new_n738), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n773), .B1(new_n784), .B2(new_n795), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n791), .A2(new_n738), .A3(new_n794), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n782), .A2(new_n597), .A3(new_n652), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n798), .A2(new_n774), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n797), .A2(KEYINPUT114), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n772), .B1(new_n796), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n802), .B1(new_n772), .B2(new_n803), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n801), .A2(new_n804), .ZN(new_n806));
  OAI21_X1  g620(.A(KEYINPUT54), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n712), .A2(new_n593), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n753), .A2(new_n293), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n722), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n771), .B(new_n812), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n784), .A2(new_n795), .A3(new_n773), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT114), .B1(new_n797), .B2(new_n799), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n802), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n784), .A2(new_n795), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n818), .A2(KEYINPUT116), .A3(KEYINPUT53), .A4(new_n813), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n793), .A2(new_n740), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(new_n789), .B2(new_n790), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n799), .A2(KEYINPUT53), .A3(new_n822), .A4(new_n738), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n820), .B1(new_n823), .B2(new_n772), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n819), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n817), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n807), .A2(new_n811), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT51), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n696), .A2(new_n732), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT119), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n596), .A3(new_n293), .A4(new_n678), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n621), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(new_n751), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n809), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n831), .A2(new_n651), .A3(new_n712), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT120), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n836), .A2(new_n841), .A3(new_n838), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n829), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n550), .A2(new_n694), .ZN(new_n844));
  OAI22_X1  g658(.A1(new_n763), .A2(new_n765), .B1(new_n415), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n758), .A3(new_n810), .ZN(new_n846));
  NAND2_X1  g660(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n695), .A2(new_n409), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(KEYINPUT117), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n808), .A2(new_n849), .A3(new_n809), .ZN(new_n850));
  NOR2_X1   g664(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n686), .B1(new_n848), .B2(KEYINPUT117), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n851), .B1(new_n850), .B2(new_n852), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n847), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n843), .A2(new_n846), .A3(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n855), .A2(new_n836), .A3(new_n846), .A4(new_n838), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n292), .B1(new_n857), .B2(new_n829), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n833), .A2(new_n622), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n734), .A2(new_n591), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n831), .A2(new_n860), .A3(new_n837), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT48), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n856), .A2(new_n858), .A3(new_n859), .A4(new_n862), .ZN(new_n863));
  OAI22_X1  g677(.A1(new_n828), .A2(new_n863), .B1(G952), .B2(G953), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n844), .A2(KEYINPUT49), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT111), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n678), .A2(new_n410), .A3(new_n752), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n866), .A2(new_n414), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n844), .A2(KEYINPUT49), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n868), .A2(new_n685), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n864), .B1(new_n591), .B2(new_n870), .ZN(G75));
  NAND2_X1  g685(.A1(new_n796), .A2(new_n800), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT53), .B1(new_n872), .B2(new_n813), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n819), .A2(new_n824), .ZN(new_n874));
  OAI211_X1 g688(.A(G210), .B(G902), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT56), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n875), .A2(KEYINPUT121), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n366), .A2(new_n390), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n878), .B(new_n388), .Z(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT55), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n877), .A2(new_n880), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n281), .A2(G952), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(G51));
  OAI21_X1  g698(.A(KEYINPUT57), .B1(new_n464), .B2(new_n251), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n826), .B1(new_n817), .B2(new_n825), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n873), .A2(new_n874), .A3(KEYINPUT54), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n464), .A2(new_n251), .A3(KEYINPUT57), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n546), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n251), .B1(new_n817), .B2(new_n825), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n891), .A2(G469), .A3(new_n742), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n883), .B1(new_n890), .B2(new_n892), .ZN(G54));
  NAND3_X1  g707(.A1(new_n891), .A2(KEYINPUT58), .A3(G475), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n894), .A2(new_n243), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n243), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n895), .A2(new_n896), .A3(new_n883), .ZN(G60));
  INV_X1    g711(.A(new_n883), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n614), .B(KEYINPUT59), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n807), .B2(new_n827), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n898), .B1(new_n900), .B2(new_n620), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n886), .A2(new_n887), .ZN(new_n902));
  INV_X1    g716(.A(new_n620), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n902), .A2(new_n903), .A3(new_n899), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n901), .A2(new_n904), .ZN(G63));
  XNOR2_X1  g719(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(G217), .A2(G902), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT60), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n910), .B1(new_n873), .B2(new_n874), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n575), .A2(new_n576), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n883), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n643), .B(new_n910), .C1(new_n873), .C2(new_n874), .ZN(new_n914));
  AOI211_X1 g728(.A(KEYINPUT122), .B(new_n907), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n909), .B1(new_n817), .B2(new_n825), .ZN(new_n916));
  INV_X1    g730(.A(new_n912), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n898), .B(new_n914), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n906), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n915), .A2(new_n920), .ZN(G66));
  OAI21_X1  g735(.A(G953), .B1(new_n295), .B2(new_n386), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n922), .B1(new_n799), .B2(G953), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n878), .B1(G898), .B2(new_n281), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(G69));
  INV_X1    g739(.A(new_n760), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n767), .A2(new_n926), .A3(new_n738), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n725), .A2(new_n664), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n692), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n749), .A2(new_n718), .A3(new_n860), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n931), .A2(new_n932), .A3(new_n740), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n928), .A2(KEYINPUT126), .A3(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT126), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(new_n927), .B2(new_n933), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n935), .A2(new_n937), .A3(new_n281), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n512), .B(new_n206), .Z(new_n939));
  NAND2_X1  g753(.A1(G900), .A2(G953), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n939), .B(KEYINPUT124), .Z(new_n942));
  NAND2_X1  g756(.A1(new_n623), .A2(new_n778), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n669), .A2(new_n736), .A3(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n926), .A2(new_n767), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n947), .B1(new_n688), .B2(new_n930), .ZN(new_n948));
  OAI211_X1 g762(.A(KEYINPUT62), .B(new_n931), .C1(new_n671), .C2(new_n687), .ZN(new_n949));
  AOI211_X1 g763(.A(new_n945), .B(new_n946), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n942), .B1(new_n950), .B2(G953), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n941), .A2(KEYINPUT125), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n281), .B1(G227), .B2(G900), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n953), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n941), .A2(new_n951), .A3(KEYINPUT125), .A4(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n954), .A2(new_n956), .ZN(G72));
  NAND2_X1  g771(.A1(new_n935), .A2(new_n937), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n784), .B1(new_n958), .B2(new_n522), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n672), .A2(new_n540), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n496), .A2(new_n513), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n959), .B(new_n960), .C1(new_n962), .C2(new_n950), .ZN(new_n963));
  XNOR2_X1  g777(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n964));
  NAND2_X1  g778(.A1(G472), .A2(G902), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n883), .B1(new_n960), .B2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n966), .ZN(new_n968));
  OAI221_X1 g782(.A(new_n968), .B1(new_n672), .B2(new_n540), .C1(new_n805), .C2(new_n806), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n963), .A2(new_n967), .A3(new_n969), .ZN(G57));
endmodule


