//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1327, new_n1328;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n206), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n202), .A2(G50), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n208), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n211), .B1(new_n214), .B2(new_n215), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XOR2_X1   g0024(.A(G250), .B(G257), .Z(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT64), .ZN(new_n226));
  XNOR2_X1  g0026(.A(G264), .B(G270), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n228), .B(new_n233), .Z(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XNOR2_X1  g0035(.A(G107), .B(G116), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  INV_X1    g0037(.A(G50), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n238), .A2(G68), .ZN(new_n239));
  INV_X1    g0039(.A(G68), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G50), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n237), .B(new_n244), .ZN(G351));
  OAI21_X1  g0045(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n246));
  INV_X1    g0046(.A(G274), .ZN(new_n247));
  OR2_X1    g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G1), .A3(G13), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G226), .A3(new_n246), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(KEYINPUT65), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G1698), .ZN(new_n259));
  INV_X1    g0059(.A(G223), .ZN(new_n260));
  INV_X1    g0060(.A(G77), .ZN(new_n261));
  OAI22_X1  g0061(.A1(new_n259), .A2(new_n260), .B1(new_n261), .B2(new_n258), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  OAI211_X1 g0065(.A(G222), .B(new_n263), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  OR2_X1    g0066(.A1(new_n266), .A2(KEYINPUT66), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(KEYINPUT66), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n262), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n253), .B(G190), .C1(new_n269), .C2(new_n250), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT74), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n267), .A2(new_n268), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n264), .A2(new_n265), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(new_n263), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n275), .A2(G223), .B1(new_n274), .B2(G77), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n250), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n278), .A2(KEYINPUT74), .A3(G190), .A4(new_n253), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n272), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT9), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n212), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n202), .A2(G50), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(new_n206), .ZN(new_n286));
  XOR2_X1   g0086(.A(KEYINPUT8), .B(G58), .Z(new_n287));
  NOR2_X1   g0087(.A1(new_n255), .A2(G20), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n287), .A2(new_n288), .B1(G150), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT67), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n286), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT8), .B(G58), .ZN(new_n293));
  INV_X1    g0093(.A(new_n288), .ZN(new_n294));
  INV_X1    g0094(.A(G150), .ZN(new_n295));
  INV_X1    g0095(.A(new_n289), .ZN(new_n296));
  OAI22_X1  g0096(.A1(new_n293), .A2(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT67), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n284), .B1(new_n292), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n205), .A2(G20), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G50), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT69), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n301), .B(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT68), .ZN(new_n304));
  INV_X1    g0104(.A(G13), .ZN(new_n305));
  NOR3_X1   g0105(.A1(new_n305), .A2(new_n206), .A3(G1), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n304), .B1(new_n306), .B2(new_n283), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NOR3_X1   g0108(.A1(new_n306), .A2(new_n283), .A3(new_n304), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n303), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n306), .A2(new_n238), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n281), .B1(new_n299), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n298), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n297), .A2(KEYINPUT67), .B1(new_n206), .B2(new_n285), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n283), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n309), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n307), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n318), .A2(new_n303), .B1(new_n238), .B2(new_n306), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n316), .A2(new_n319), .A3(KEYINPUT9), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT73), .B(G200), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT65), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n252), .B(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n322), .B1(new_n277), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n313), .A2(new_n320), .A3(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT10), .B1(new_n280), .B2(new_n326), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n313), .A2(new_n320), .A3(new_n325), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n272), .A2(new_n279), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT10), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n306), .A2(new_n283), .ZN(new_n333));
  INV_X1    g0133(.A(new_n300), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(new_n261), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n333), .A2(new_n335), .B1(new_n261), .B2(new_n306), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n293), .A2(new_n296), .B1(new_n206), .B2(new_n261), .ZN(new_n337));
  XNOR2_X1  g0137(.A(KEYINPUT15), .B(G87), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n337), .A2(KEYINPUT71), .B1(new_n339), .B2(new_n288), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT71), .ZN(new_n341));
  OAI221_X1 g0141(.A(new_n341), .B1(new_n206), .B2(new_n261), .C1(new_n293), .C2(new_n296), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n284), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n343), .A2(KEYINPUT72), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n343), .A2(KEYINPUT72), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n336), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n258), .A2(G232), .A3(new_n263), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n274), .A2(G107), .ZN(new_n348));
  INV_X1    g0148(.A(G238), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n347), .B(new_n348), .C1(new_n259), .C2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n250), .A2(G244), .A3(new_n246), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n248), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT70), .ZN(new_n356));
  INV_X1    g0156(.A(G169), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT70), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n352), .A2(new_n358), .A3(new_n354), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n356), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G179), .ZN(new_n361));
  AND3_X1   g0161(.A1(new_n352), .A2(new_n358), .A3(new_n354), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n358), .B1(new_n352), .B2(new_n354), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n346), .A2(new_n360), .A3(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n343), .B(KEYINPUT72), .ZN(new_n366));
  OAI21_X1  g0166(.A(G190), .B1(new_n362), .B2(new_n363), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n356), .A2(new_n322), .A3(new_n359), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n366), .A2(new_n367), .A3(new_n368), .A4(new_n336), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n278), .A2(new_n361), .A3(new_n253), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n316), .A2(new_n319), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n357), .B1(new_n277), .B2(new_n324), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n365), .A2(new_n369), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n306), .A2(new_n240), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n375), .B(KEYINPUT12), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n289), .A2(G50), .B1(G20), .B2(new_n240), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n294), .B2(new_n261), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n378), .A2(KEYINPUT11), .A3(new_n283), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n333), .A2(G68), .A3(new_n300), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n376), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT11), .B1(new_n378), .B2(new_n283), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n357), .A2(KEYINPUT76), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n258), .A2(G232), .A3(G1698), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n258), .A2(G226), .A3(new_n263), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G33), .A2(G97), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n351), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n250), .A2(G238), .A3(new_n246), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT75), .B1(new_n248), .B2(new_n392), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n248), .A2(KEYINPUT75), .A3(new_n392), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n391), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT13), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT13), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n391), .B(new_n397), .C1(new_n393), .C2(new_n394), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n386), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT14), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n396), .A2(new_n398), .ZN(new_n401));
  OAI22_X1  g0201(.A1(new_n399), .A2(new_n400), .B1(new_n401), .B2(new_n361), .ZN(new_n402));
  AOI211_X1 g0202(.A(KEYINPUT14), .B(new_n386), .C1(new_n396), .C2(new_n398), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n384), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n401), .A2(G200), .ZN(new_n405));
  INV_X1    g0205(.A(G190), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n405), .B(new_n383), .C1(new_n401), .C2(new_n406), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n332), .A2(new_n374), .A3(new_n404), .A4(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n293), .A2(new_n334), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n318), .A2(new_n409), .B1(new_n306), .B2(new_n293), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G58), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n412), .A2(new_n240), .ZN(new_n413));
  OAI21_X1  g0213(.A(G20), .B1(new_n413), .B2(new_n201), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n289), .A2(G159), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n256), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n257), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT77), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n264), .B2(new_n265), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n256), .A2(KEYINPUT77), .A3(new_n257), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n422), .A3(new_n206), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT7), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n419), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI211_X1 g0225(.A(KEYINPUT16), .B(new_n417), .C1(new_n425), .C2(new_n240), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n426), .A2(new_n283), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT16), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT78), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n418), .B(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n424), .B1(new_n258), .B2(G20), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n240), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n428), .B1(new_n432), .B2(new_n416), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n411), .B1(new_n427), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(G226), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(G1698), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n258), .B(new_n436), .C1(G223), .C2(G1698), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G33), .A2(G87), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n250), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n250), .A2(new_n246), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n248), .B1(new_n440), .B2(new_n230), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n439), .A2(new_n361), .A3(new_n441), .ZN(new_n442));
  OR2_X1    g0242(.A1(new_n439), .A2(new_n441), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n442), .B1(G169), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT18), .B1(new_n434), .B2(new_n444), .ZN(new_n445));
  AND2_X1   g0245(.A1(KEYINPUT79), .A2(G190), .ZN(new_n446));
  NOR2_X1   g0246(.A1(KEYINPUT79), .A2(G190), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n439), .A2(new_n448), .A3(new_n441), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n449), .B1(G200), .B2(new_n443), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n434), .A2(KEYINPUT17), .A3(new_n450), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n418), .A2(new_n429), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n418), .A2(new_n429), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n431), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n416), .B1(new_n454), .B2(G68), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n283), .B(new_n426), .C1(new_n455), .C2(KEYINPUT16), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n410), .ZN(new_n457));
  INV_X1    g0257(.A(new_n444), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT18), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n456), .A2(new_n450), .A3(new_n410), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT17), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n445), .A2(new_n451), .A3(new_n460), .A4(new_n463), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n464), .A2(KEYINPUT80), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n464), .A2(KEYINPUT80), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n408), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n205), .A2(G33), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n333), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(G107), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n306), .A2(KEYINPUT25), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT25), .B1(new_n306), .B2(new_n470), .ZN(new_n472));
  OAI22_X1  g0272(.A1(new_n469), .A2(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n470), .A2(G20), .ZN(new_n474));
  XNOR2_X1  g0274(.A(new_n474), .B(KEYINPUT23), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT87), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G116), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n476), .B1(new_n477), .B2(G20), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n206), .A2(KEYINPUT87), .A3(G33), .A4(G116), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n206), .B(G87), .C1(new_n264), .C2(new_n265), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n482), .A2(KEYINPUT22), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n482), .A2(KEYINPUT22), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT24), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT24), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n481), .B(new_n487), .C1(new_n483), .C2(new_n484), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n473), .B1(new_n489), .B2(new_n283), .ZN(new_n490));
  OAI211_X1 g0290(.A(G257), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n491));
  OAI211_X1 g0291(.A(G250), .B(new_n263), .C1(new_n264), .C2(new_n265), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G33), .A2(G294), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT88), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT88), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n491), .A2(new_n492), .A3(new_n496), .A4(new_n493), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n495), .A2(new_n497), .A3(new_n351), .ZN(new_n498));
  XNOR2_X1  g0298(.A(KEYINPUT5), .B(G41), .ZN(new_n499));
  INV_X1    g0299(.A(G45), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n500), .A2(G1), .ZN(new_n501));
  INV_X1    g0301(.A(new_n212), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n499), .A2(new_n501), .B1(new_n502), .B2(new_n249), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G264), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT89), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT89), .ZN(new_n506));
  AND2_X1   g0306(.A1(KEYINPUT5), .A2(G41), .ZN(new_n507));
  NOR2_X1   g0307(.A1(KEYINPUT5), .A2(G41), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n501), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AND4_X1   g0309(.A1(new_n506), .A2(new_n509), .A3(G264), .A4(new_n250), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(KEYINPUT90), .B1(new_n498), .B2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n499), .A2(G274), .A3(new_n250), .A4(new_n501), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n506), .B1(new_n503), .B2(G264), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n515), .A2(new_n510), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n495), .A2(new_n497), .A3(new_n351), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT90), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n513), .A2(G179), .A3(new_n514), .A4(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n516), .A2(new_n517), .A3(new_n514), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G169), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n490), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n513), .A2(new_n514), .A3(new_n519), .ZN(new_n524));
  INV_X1    g0324(.A(G200), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OR2_X1    g0326(.A1(new_n521), .A2(G190), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n523), .B1(new_n528), .B2(new_n490), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n509), .A2(G270), .A3(new_n250), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n530), .A2(new_n514), .ZN(new_n531));
  OAI211_X1 g0331(.A(G264), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n532));
  OAI211_X1 g0332(.A(G257), .B(new_n263), .C1(new_n264), .C2(new_n265), .ZN(new_n533));
  INV_X1    g0333(.A(G303), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n532), .B(new_n533), .C1(new_n534), .C2(new_n258), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n351), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n333), .A2(G116), .A3(new_n468), .ZN(new_n538));
  INV_X1    g0338(.A(G116), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n306), .A2(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n282), .A2(new_n212), .B1(G20), .B2(new_n539), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G283), .ZN(new_n542));
  INV_X1    g0342(.A(G97), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n542), .B(new_n206), .C1(G33), .C2(new_n543), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n541), .A2(KEYINPUT20), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(KEYINPUT20), .B1(new_n541), .B2(new_n544), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n538), .B(new_n540), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT86), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n548), .A2(KEYINPUT21), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n537), .A2(new_n547), .A3(G169), .A4(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n547), .ZN(new_n552));
  INV_X1    g0352(.A(new_n448), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n531), .A2(new_n536), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n537), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n552), .B(new_n554), .C1(new_n555), .C2(new_n525), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n537), .A2(new_n547), .A3(G169), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n549), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n555), .A2(G179), .A3(new_n547), .ZN(new_n559));
  AND4_X1   g0359(.A1(new_n551), .A2(new_n556), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n306), .A2(new_n543), .ZN(new_n561));
  XNOR2_X1  g0361(.A(new_n561), .B(KEYINPUT82), .ZN(new_n562));
  INV_X1    g0362(.A(new_n469), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n562), .B1(G97), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n289), .A2(G77), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT81), .ZN(new_n566));
  XNOR2_X1  g0366(.A(new_n565), .B(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT6), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n568), .A2(new_n543), .A3(G107), .ZN(new_n569));
  XNOR2_X1  g0369(.A(G97), .B(G107), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n569), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n567), .B1(new_n206), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(G107), .B2(new_n454), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n564), .B1(new_n573), .B2(new_n284), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n509), .A2(G257), .A3(new_n250), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n514), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n263), .A2(G244), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n577), .B1(new_n256), .B2(new_n257), .ZN(new_n578));
  OAI21_X1  g0378(.A(KEYINPUT83), .B1(new_n578), .B2(KEYINPUT4), .ZN(new_n579));
  OAI211_X1 g0379(.A(G250), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n580), .A2(new_n542), .ZN(new_n581));
  INV_X1    g0381(.A(G244), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n582), .A2(G1698), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n258), .A2(KEYINPUT4), .A3(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n583), .B1(new_n264), .B2(new_n265), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT83), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT4), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n579), .A2(new_n581), .A3(new_n584), .A4(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n576), .B1(new_n589), .B2(new_n351), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n590), .A2(new_n525), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n574), .A2(new_n591), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n586), .B1(new_n585), .B2(new_n587), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n584), .A2(new_n542), .A3(new_n580), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n250), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(KEYINPUT84), .B1(new_n597), .B2(new_n576), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT84), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n590), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n598), .A2(new_n600), .A3(G190), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n592), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n589), .A2(new_n351), .ZN(new_n603));
  INV_X1    g0403(.A(new_n576), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n599), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI211_X1 g0405(.A(KEYINPUT84), .B(new_n576), .C1(new_n589), .C2(new_n351), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n357), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n470), .B1(new_n430), .B2(new_n431), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n283), .B1(new_n608), .B2(new_n572), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n609), .A2(new_n564), .B1(new_n361), .B2(new_n590), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n205), .A2(G45), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(G250), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n351), .A2(new_n613), .B1(new_n247), .B2(new_n612), .ZN(new_n614));
  OAI211_X1 g0414(.A(G244), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n615));
  OAI211_X1 g0415(.A(G238), .B(new_n263), .C1(new_n264), .C2(new_n265), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n616), .A3(new_n477), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n614), .B1(new_n617), .B2(new_n351), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n618), .A2(G169), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n619), .B1(new_n361), .B2(new_n618), .ZN(new_n620));
  INV_X1    g0420(.A(new_n306), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n339), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n258), .A2(new_n206), .A3(G68), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(KEYINPUT85), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT19), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n288), .A2(new_n625), .A3(G97), .ZN(new_n626));
  NOR2_X1   g0426(.A1(G97), .A2(G107), .ZN(new_n627));
  INV_X1    g0427(.A(G87), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n627), .A2(new_n628), .B1(new_n389), .B2(new_n206), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n626), .B1(new_n629), .B2(new_n625), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT85), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n258), .A2(new_n631), .A3(new_n206), .A4(G68), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n624), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n622), .B1(new_n633), .B2(new_n283), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n469), .B2(new_n338), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n618), .A2(new_n321), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(G190), .B2(new_n618), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n469), .A2(new_n628), .ZN(new_n638));
  AOI211_X1 g0438(.A(new_n622), .B(new_n638), .C1(new_n633), .C2(new_n283), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n620), .A2(new_n635), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  AND4_X1   g0440(.A1(new_n560), .A2(new_n602), .A3(new_n611), .A4(new_n640), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n467), .A2(new_n529), .A3(new_n641), .ZN(G372));
  NAND2_X1  g0442(.A1(new_n520), .A2(new_n522), .ZN(new_n643));
  INV_X1    g0443(.A(new_n490), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n558), .A2(new_n559), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(new_n551), .A3(new_n646), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n602), .A2(new_n611), .A3(new_n640), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n644), .B1(new_n526), .B2(new_n527), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n620), .A2(new_n635), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT26), .ZN(new_n653));
  INV_X1    g0453(.A(new_n640), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n653), .B1(new_n654), .B2(new_n611), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n640), .A2(new_n607), .A3(KEYINPUT26), .A4(new_n610), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n652), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n467), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n373), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n445), .A2(new_n460), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n404), .A2(new_n365), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n407), .A2(new_n463), .A3(new_n451), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT91), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n330), .B1(new_n328), .B2(new_n329), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n327), .A2(KEYINPUT91), .A3(new_n331), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n660), .B1(new_n664), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n659), .A2(new_n671), .ZN(G369));
  NAND3_X1  g0472(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(new_n675), .A3(G213), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n644), .A2(new_n678), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n529), .A2(new_n679), .B1(new_n523), .B2(new_n678), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n646), .A2(new_n551), .ZN(new_n681));
  INV_X1    g0481(.A(new_n678), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n552), .A2(new_n682), .ZN(new_n683));
  MUX2_X1   g0483(.A(new_n560), .B(new_n681), .S(new_n683), .Z(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G330), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n681), .A2(new_n682), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n688), .A2(new_n649), .A3(new_n523), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n689), .B1(new_n523), .B2(new_n682), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n687), .A2(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n209), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n627), .A2(new_n628), .A3(new_n539), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n694), .A2(G1), .A3(new_n696), .ZN(new_n697));
  OAI22_X1  g0497(.A1(new_n697), .A2(KEYINPUT92), .B1(new_n215), .B2(new_n694), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n698), .B1(KEYINPUT92), .B2(new_n697), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT28), .Z(new_n700));
  NAND2_X1  g0500(.A1(new_n658), .A2(new_n682), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(KEYINPUT29), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n678), .B1(new_n651), .B2(new_n657), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT29), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  INV_X1    g0507(.A(new_n618), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n537), .A2(new_n708), .A3(new_n361), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n598), .A2(new_n600), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n513), .A2(new_n519), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n707), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n605), .A2(new_n606), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n518), .B1(new_n516), .B2(new_n517), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n713), .A2(new_n716), .A3(KEYINPUT30), .A4(new_n709), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT93), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n537), .A2(new_n708), .A3(new_n718), .A4(new_n361), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n603), .A2(new_n604), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n537), .A2(new_n708), .A3(new_n361), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT93), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n524), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n712), .A2(new_n717), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n678), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT31), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n641), .A2(new_n529), .A3(new_n682), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G330), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n706), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n700), .B1(new_n733), .B2(G1), .ZN(G364));
  NOR2_X1   g0534(.A1(new_n305), .A2(G20), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n205), .B1(new_n735), .B2(G45), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n693), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n212), .B1(G20), .B2(new_n357), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR4_X1   g0541(.A1(new_n321), .A2(new_n206), .A3(G179), .A4(G190), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n742), .A2(KEYINPUT96), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(KEYINPUT96), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G107), .ZN(new_n747));
  NAND3_X1  g0547(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n448), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n748), .A2(G190), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n750), .A2(new_n238), .B1(new_n240), .B2(new_n752), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n206), .A2(new_n361), .A3(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n553), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n274), .B(new_n753), .C1(G58), .C2(new_n756), .ZN(new_n757));
  NOR4_X1   g0557(.A1(new_n321), .A2(new_n206), .A3(G179), .A4(new_n406), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G179), .A2(G200), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(G20), .A3(new_n406), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n761), .A2(KEYINPUT32), .A3(G159), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT32), .ZN(new_n763));
  INV_X1    g0563(.A(G159), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n763), .B1(new_n760), .B2(new_n764), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n758), .A2(G87), .B1(new_n762), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n754), .A2(new_n406), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n767), .A2(KEYINPUT95), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(KEYINPUT95), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n206), .B1(new_n759), .B2(G190), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n771), .B(KEYINPUT97), .Z(new_n772));
  AOI22_X1  g0572(.A1(new_n770), .A2(G77), .B1(new_n772), .B2(G97), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n747), .A2(new_n757), .A3(new_n766), .A4(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n258), .B1(new_n761), .B2(G329), .ZN(new_n775));
  INV_X1    g0575(.A(G294), .ZN(new_n776));
  INV_X1    g0576(.A(new_n758), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n775), .B1(new_n776), .B2(new_n771), .C1(new_n777), .C2(new_n534), .ZN(new_n778));
  INV_X1    g0578(.A(G326), .ZN(new_n779));
  INV_X1    g0579(.A(G322), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n750), .A2(new_n779), .B1(new_n755), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G311), .ZN(new_n782));
  XOR2_X1   g0582(.A(KEYINPUT33), .B(G317), .Z(new_n783));
  OAI22_X1  g0583(.A1(new_n767), .A2(new_n782), .B1(new_n752), .B2(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n778), .A2(new_n781), .A3(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G283), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n785), .B1(new_n786), .B2(new_n745), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n741), .B1(new_n774), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G13), .A2(G33), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(G20), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n740), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n692), .A2(new_n274), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n793), .A2(G355), .B1(new_n539), .B2(new_n692), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n421), .A2(new_n422), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n692), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(G45), .B2(new_n215), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n244), .A2(new_n500), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n794), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n739), .B(new_n788), .C1(new_n792), .C2(new_n799), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT98), .Z(new_n801));
  INV_X1    g0601(.A(new_n791), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n684), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n684), .A2(G330), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n804), .A2(KEYINPUT94), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(KEYINPUT94), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n805), .A2(new_n685), .A3(new_n806), .A4(new_n739), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n803), .A2(new_n807), .ZN(G396));
  OAI21_X1  g0608(.A(new_n274), .B1(new_n760), .B2(new_n782), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n750), .A2(new_n534), .B1(new_n755), .B2(new_n776), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n809), .B(new_n810), .C1(G283), .C2(new_n751), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n746), .A2(G87), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n758), .A2(G107), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n770), .A2(G116), .B1(new_n772), .B2(G97), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n811), .A2(new_n812), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n756), .A2(G143), .B1(G137), .B2(new_n749), .ZN(new_n816));
  INV_X1    g0616(.A(new_n770), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n816), .B1(new_n295), .B2(new_n752), .C1(new_n817), .C2(new_n764), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT34), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n746), .A2(G68), .ZN(new_n821));
  INV_X1    g0621(.A(G132), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n795), .B1(new_n412), .B2(new_n771), .C1(new_n822), .C2(new_n760), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(G50), .B2(new_n758), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n820), .A2(new_n821), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n818), .A2(new_n819), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n815), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n740), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n740), .A2(new_n789), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n739), .B1(new_n261), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n365), .A2(new_n678), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n346), .A2(new_n678), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n369), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(new_n365), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n828), .B(new_n830), .C1(new_n837), .C2(new_n790), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n701), .A2(new_n836), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n703), .A2(new_n837), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n839), .A2(KEYINPUT99), .A3(new_n840), .ZN(new_n841));
  OR3_X1    g0641(.A1(new_n703), .A2(KEYINPUT99), .A3(new_n837), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n841), .A2(new_n732), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n739), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n732), .B1(new_n841), .B2(new_n842), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n838), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT100), .ZN(G384));
  INV_X1    g0647(.A(new_n571), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n539), .B(new_n214), .C1(new_n848), .C2(KEYINPUT35), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(KEYINPUT35), .B2(new_n848), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT36), .Z(new_n851));
  OR3_X1    g0651(.A1(new_n215), .A2(new_n261), .A3(new_n413), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n205), .B(G13), .C1(new_n852), .C2(new_n239), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n456), .A2(new_n410), .A3(new_n450), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n444), .B1(new_n456), .B2(new_n410), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT37), .ZN(new_n858));
  INV_X1    g0658(.A(new_n676), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT101), .B1(new_n457), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT101), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n861), .B(new_n676), .C1(new_n456), .C2(new_n410), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n857), .B(new_n858), .C1(new_n860), .C2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n417), .B1(new_n425), .B2(new_n240), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n864), .A2(new_n428), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n426), .A2(new_n283), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n410), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n859), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n461), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n867), .A2(new_n458), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT37), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n863), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n868), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n464), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n872), .A2(KEYINPUT38), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT102), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT102), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n872), .A2(new_n877), .A3(KEYINPUT38), .A4(new_n874), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n872), .A2(new_n874), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n876), .A2(new_n878), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n384), .A2(new_n678), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n404), .A2(new_n407), .A3(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n384), .B(new_n678), .C1(new_n402), .C2(new_n403), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n836), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(KEYINPUT105), .A2(KEYINPUT31), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n725), .A2(new_n678), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n887), .B1(new_n725), .B2(new_n678), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n729), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT40), .B1(new_n882), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n886), .A2(new_n890), .A3(KEYINPUT40), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n863), .A2(KEYINPUT103), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n861), .B1(new_n434), .B2(new_n676), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n457), .A2(KEYINPUT101), .A3(new_n859), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT103), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n897), .A2(new_n898), .A3(new_n858), .A4(new_n857), .ZN(new_n899));
  INV_X1    g0699(.A(new_n857), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n860), .A2(new_n862), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT37), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n894), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n464), .A2(new_n901), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT104), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n464), .A2(KEYINPUT104), .A3(new_n901), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n880), .B1(new_n903), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n893), .B1(new_n909), .B2(new_n875), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n892), .A2(new_n910), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n911), .A2(new_n467), .A3(new_n890), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n911), .B1(new_n467), .B2(new_n890), .ZN(new_n913));
  INV_X1    g0713(.A(G330), .ZN(new_n914));
  OR3_X1    g0714(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n909), .A2(new_n916), .A3(new_n875), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n863), .A2(new_n871), .B1(new_n464), .B2(new_n873), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n878), .B1(KEYINPUT38), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n877), .B1(new_n918), .B2(KEYINPUT38), .ZN(new_n920));
  OAI21_X1  g0720(.A(KEYINPUT39), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n404), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n682), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n661), .A2(new_n859), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n840), .A2(new_n832), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n884), .A2(new_n885), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n882), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n926), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n467), .B1(new_n702), .B2(new_n705), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n671), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n931), .B(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n915), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n205), .B2(new_n735), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n915), .A2(new_n934), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n854), .B1(new_n936), .B2(new_n937), .ZN(G367));
  NAND2_X1  g0738(.A1(new_n574), .A2(new_n678), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n602), .A2(new_n611), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n611), .B2(new_n682), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT106), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n523), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n678), .B1(new_n944), .B2(new_n611), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT43), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n640), .B1(new_n639), .B2(new_n682), .ZN(new_n948));
  INV_X1    g0748(.A(new_n639), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n652), .A2(new_n949), .A3(new_n678), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n689), .A2(new_n941), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT42), .Z(new_n954));
  NAND4_X1  g0754(.A1(new_n946), .A2(new_n947), .A3(new_n952), .A4(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n687), .A2(new_n942), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n952), .A2(new_n947), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n958));
  INV_X1    g0758(.A(new_n954), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n957), .B(new_n958), .C1(new_n945), .C2(new_n959), .ZN(new_n960));
  AND3_X1   g0760(.A1(new_n955), .A2(new_n956), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n956), .B1(new_n955), .B2(new_n960), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n693), .B(KEYINPUT41), .Z(new_n964));
  NOR2_X1   g0764(.A1(new_n690), .A2(new_n941), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT44), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n690), .A2(new_n941), .ZN(new_n967));
  XOR2_X1   g0767(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n968));
  XNOR2_X1  g0768(.A(new_n967), .B(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n686), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n706), .A2(new_n732), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT108), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n689), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(KEYINPUT108), .B1(new_n680), .B2(new_n688), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n975), .B2(new_n689), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n976), .A2(G330), .A3(new_n684), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n685), .B(new_n974), .C1(new_n975), .C2(new_n689), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n972), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n966), .A2(new_n687), .A3(new_n969), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n971), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n964), .B1(new_n981), .B2(new_n733), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n963), .B1(new_n982), .B2(new_n737), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n228), .A2(new_n796), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n984), .B(new_n792), .C1(new_n209), .C2(new_n338), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT109), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n985), .A2(new_n986), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n987), .A2(new_n988), .A3(new_n739), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n770), .A2(G50), .B1(G159), .B2(new_n751), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT111), .ZN(new_n991));
  INV_X1    g0791(.A(G137), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n258), .B1(new_n992), .B2(new_n760), .C1(new_n755), .C2(new_n295), .ZN(new_n993));
  INV_X1    g0793(.A(new_n742), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n412), .A2(new_n777), .B1(new_n994), .B2(new_n261), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n993), .B(new_n995), .C1(G143), .C2(new_n749), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n772), .A2(G68), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n991), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n777), .A2(new_n539), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n999), .A2(KEYINPUT46), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(G283), .B2(new_n770), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n750), .A2(new_n782), .B1(new_n755), .B2(new_n534), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT110), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n752), .A2(new_n776), .B1(new_n470), .B2(new_n771), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n795), .ZN(new_n1006));
  INV_X1    g0806(.A(G317), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1006), .B1(new_n1007), .B2(new_n760), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1005), .B(new_n1008), .C1(G97), .C2(new_n742), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n999), .A2(KEYINPUT46), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1001), .A2(new_n1004), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n998), .A2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT47), .Z(new_n1013));
  OAI221_X1 g0813(.A(new_n989), .B1(new_n802), .B2(new_n951), .C1(new_n1013), .C2(new_n741), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n983), .A2(new_n1014), .ZN(G387));
  NAND2_X1  g0815(.A1(new_n977), .A2(new_n978), .ZN(new_n1016));
  OAI21_X1  g0816(.A(KEYINPUT114), .B1(new_n733), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT114), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n972), .A2(new_n978), .A3(new_n1018), .A4(new_n977), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n733), .A2(new_n1016), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1017), .A2(new_n1019), .A3(new_n693), .A4(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n793), .A2(new_n695), .B1(new_n470), .B2(new_n692), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n233), .A2(new_n500), .ZN(new_n1023));
  AOI21_X1  g0823(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n287), .A2(new_n238), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n696), .B(new_n1024), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n796), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1022), .B1(new_n1023), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n739), .B1(new_n1030), .B2(new_n792), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1006), .B1(G150), .B2(new_n761), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n749), .A2(KEYINPUT113), .A3(G159), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n758), .A2(G77), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT113), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n750), .B2(new_n764), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .A4(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n772), .A2(new_n339), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n767), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n1039), .A2(G68), .B1(new_n287), .B2(new_n751), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1038), .B(new_n1040), .C1(new_n238), .C2(new_n755), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1037), .B(new_n1041), .C1(G97), .C2(new_n746), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n994), .A2(new_n539), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1006), .B1(new_n779), .B2(new_n760), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n749), .A2(G322), .B1(G311), .B2(new_n751), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n1007), .B2(new_n755), .C1(new_n817), .C2(new_n534), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1047), .A2(KEYINPUT48), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1047), .A2(KEYINPUT48), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n777), .A2(new_n776), .B1(new_n786), .B2(new_n771), .ZN(new_n1050));
  NOR3_X1   g0850(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n1043), .B(new_n1044), .C1(new_n1051), .C2(KEYINPUT49), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1051), .A2(KEYINPUT49), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1042), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1031), .B1(new_n1054), .B2(new_n741), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n680), .B2(new_n791), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n1016), .B2(new_n737), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1021), .A2(new_n1057), .ZN(G393));
  NAND3_X1  g0858(.A1(new_n971), .A2(new_n737), .A3(new_n980), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n796), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n792), .B1(new_n543), .B2(new_n209), .C1(new_n1060), .C2(new_n237), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n738), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n750), .A2(new_n1007), .B1(new_n755), .B2(new_n782), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT52), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n767), .A2(new_n776), .B1(new_n539), .B2(new_n771), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n274), .B1(new_n780), .B2(new_n760), .C1(new_n752), .C2(new_n534), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(G283), .C2(new_n758), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n747), .A2(new_n1064), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1006), .B1(G143), .B2(new_n761), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n812), .B(new_n1069), .C1(new_n240), .C2(new_n777), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT115), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n770), .A2(new_n287), .B1(G50), .B2(new_n751), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1073), .A2(KEYINPUT116), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(KEYINPUT116), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n772), .A2(G77), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n750), .A2(new_n295), .B1(new_n755), .B2(new_n764), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT51), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .A4(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1068), .B1(new_n1071), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1062), .B1(new_n1080), .B2(new_n740), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n943), .B2(new_n802), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n981), .A2(new_n693), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n979), .B1(new_n971), .B2(new_n980), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1059), .B(new_n1082), .C1(new_n1083), .C2(new_n1084), .ZN(G390));
  AOI21_X1  g0885(.A(new_n831), .B1(new_n703), .B2(new_n837), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n891), .A2(G330), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n929), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n732), .B2(new_n836), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1086), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n731), .A2(new_n886), .A3(G330), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT118), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n731), .A2(new_n886), .A3(KEYINPUT118), .A4(G330), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n890), .A2(G330), .A3(new_n837), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n929), .A2(KEYINPUT117), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT117), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n884), .A2(new_n1099), .A3(new_n885), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1097), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT120), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1097), .A2(new_n1101), .A3(KEYINPUT120), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1096), .A2(new_n1104), .A3(new_n1086), .A4(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT121), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n1097), .A2(KEYINPUT120), .A3(new_n1101), .ZN(new_n1109));
  AOI21_X1  g0909(.A(KEYINPUT120), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n928), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1112));
  AOI21_X1  g0912(.A(KEYINPUT121), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1091), .B1(new_n1108), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n924), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n917), .A2(new_n1115), .A3(new_n921), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n907), .ZN(new_n1117));
  AOI21_X1  g0917(.A(KEYINPUT104), .B1(new_n464), .B2(new_n901), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n894), .A2(new_n902), .A3(new_n899), .ZN(new_n1120));
  AOI21_X1  g0920(.A(KEYINPUT38), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n875), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n924), .B1(new_n1086), .B2(new_n1101), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  AND3_X1   g0923(.A1(new_n1116), .A2(new_n1123), .A3(new_n1096), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1087), .B1(new_n1116), .B2(new_n1123), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n467), .A2(G330), .A3(new_n890), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n932), .A2(new_n1127), .A3(new_n671), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(KEYINPUT119), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT119), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n932), .A2(new_n1127), .A3(new_n1130), .A4(new_n671), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1114), .A2(new_n1126), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1116), .A2(new_n1123), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1087), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1116), .A2(new_n1123), .A3(new_n1096), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1111), .A2(KEYINPUT121), .A3(new_n1112), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1090), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1139), .B1(new_n1142), .B2(new_n1132), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1134), .A2(new_n1143), .A3(new_n693), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT123), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n739), .B1(new_n293), .B2(new_n829), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n1146), .B(KEYINPUT122), .Z(new_n1147));
  OAI21_X1  g0947(.A(new_n274), .B1(new_n760), .B2(new_n776), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n750), .A2(new_n786), .B1(new_n755), .B2(new_n539), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1148), .B(new_n1149), .C1(G107), .C2(new_n751), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n758), .A2(G87), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n770), .A2(G97), .B1(new_n772), .B2(G77), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1150), .A2(new_n821), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n755), .A2(new_n822), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n274), .B1(new_n761), .B2(G125), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n992), .B2(new_n752), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1154), .B(new_n1156), .C1(G128), .C2(new_n749), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT54), .B(G143), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n770), .A2(new_n1159), .B1(new_n772), .B2(G159), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1157), .B(new_n1160), .C1(new_n238), .C2(new_n994), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n758), .A2(G150), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT53), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1153), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1147), .B1(new_n1164), .B2(new_n740), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n922), .B2(new_n790), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1145), .B(new_n1166), .C1(new_n1139), .C2(new_n736), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1166), .B1(new_n1139), .B2(new_n736), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(KEYINPUT123), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1144), .A2(new_n1167), .A3(new_n1169), .ZN(G378));
  OAI21_X1  g0970(.A(new_n1133), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n668), .A2(new_n669), .A3(new_n373), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n371), .A2(new_n859), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n668), .A2(new_n669), .A3(new_n373), .A4(new_n1173), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1177), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n911), .B2(G330), .ZN(new_n1182));
  NOR4_X1   g0982(.A1(new_n892), .A2(new_n910), .A3(new_n1180), .A4(new_n914), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n931), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(KEYINPUT40), .B(new_n891), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n882), .A2(new_n891), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1185), .B(G330), .C1(new_n1186), .C2(KEYINPUT40), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n1180), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n930), .A2(new_n927), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n925), .B2(new_n922), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n911), .A2(G330), .A3(new_n1181), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1188), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1184), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1171), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT57), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n694), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT125), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1184), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1197), .B1(new_n1184), .B2(new_n1192), .ZN(new_n1199));
  OAI211_X1 g0999(.A(KEYINPUT57), .B(new_n1171), .C1(new_n1198), .C2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1196), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1193), .A2(new_n737), .ZN(new_n1202));
  INV_X1    g1002(.A(G41), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1006), .A2(new_n1203), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1034), .B1(new_n786), .B2(new_n760), .C1(new_n338), .C2(new_n767), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1204), .B(new_n1205), .C1(G58), .C2(new_n742), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n749), .A2(G116), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n756), .A2(G107), .B1(G97), .B2(new_n751), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1206), .A2(new_n997), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT58), .ZN(new_n1210));
  AOI21_X1  g1010(.A(G50), .B1(new_n255), .B2(new_n1203), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1209), .A2(new_n1210), .B1(new_n1204), .B2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n1210), .B2(new_n1209), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n767), .A2(new_n992), .B1(new_n752), .B2(new_n822), .ZN(new_n1214));
  AND2_X1   g1014(.A1(new_n756), .A2(G128), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1214), .B(new_n1215), .C1(G125), .C2(new_n749), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n772), .A2(G150), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(new_n777), .C2(new_n1158), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n742), .A2(G159), .ZN(new_n1220));
  AOI211_X1 g1020(.A(G33), .B(G41), .C1(new_n761), .C2(G124), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n740), .B1(new_n1213), .B2(new_n1224), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT124), .Z(new_n1226));
  AOI21_X1  g1026(.A(new_n739), .B1(new_n238), .B2(new_n829), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1226), .B(new_n1227), .C1(new_n1181), .C2(new_n790), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1202), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1201), .A2(new_n1230), .ZN(G375));
  AOI21_X1  g1031(.A(new_n739), .B1(new_n240), .B2(new_n829), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1038), .B1(new_n817), .B2(new_n470), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n274), .B1(new_n760), .B2(new_n534), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n750), .A2(new_n776), .B1(new_n755), .B2(new_n786), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1234), .B(new_n1235), .C1(G116), .C2(new_n751), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n543), .B2(new_n777), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n1233), .B(new_n1237), .C1(G77), .C2(new_n746), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1039), .A2(G150), .B1(new_n749), .B2(G132), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1239), .B1(new_n992), .B2(new_n755), .C1(new_n752), .C2(new_n1158), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1006), .B1(G128), .B2(new_n761), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1241), .B1(new_n994), .B2(new_n412), .C1(new_n764), .C2(new_n777), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1240), .B(new_n1242), .C1(G50), .C2(new_n772), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1238), .A2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1232), .B1(new_n1244), .B2(new_n741), .ZN(new_n1245));
  XOR2_X1   g1045(.A(new_n1245), .B(KEYINPUT126), .Z(new_n1246));
  NAND2_X1  g1046(.A1(new_n1101), .A2(new_n789), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n1142), .B2(new_n736), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n964), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n1142), .B2(new_n1132), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1142), .A2(new_n1132), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1250), .B1(new_n1252), .B2(new_n1254), .ZN(G381));
  AOI21_X1  g1055(.A(new_n1229), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1144), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(G390), .ZN(new_n1259));
  INV_X1    g1059(.A(G384), .ZN(new_n1260));
  INV_X1    g1060(.A(G396), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1021), .A2(new_n1261), .A3(new_n1057), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1259), .A2(new_n1260), .A3(new_n1263), .ZN(new_n1264));
  OR4_X1    g1064(.A1(G387), .A2(new_n1258), .A3(G381), .A4(new_n1264), .ZN(G407));
  OAI211_X1 g1065(.A(G407), .B(G213), .C1(G343), .C2(new_n1258), .ZN(G409));
  NAND3_X1  g1066(.A1(new_n1171), .A2(new_n1251), .A3(new_n1193), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1267), .A2(new_n1228), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n737), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1257), .A2(new_n1268), .A3(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n677), .A2(G213), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1270), .B(new_n1271), .C1(new_n1256), .C2(new_n1257), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1273), .A2(KEYINPUT60), .A3(new_n1132), .A4(new_n1091), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n693), .ZN(new_n1275));
  OAI21_X1  g1075(.A(KEYINPUT60), .B1(new_n1142), .B2(new_n1132), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1275), .B1(new_n1253), .B2(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(G384), .B1(new_n1277), .B2(new_n1249), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1275), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1276), .A2(new_n1253), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1249), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1260), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1278), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(KEYINPUT62), .B1(new_n1272), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT61), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1281), .A2(new_n1260), .ZN(new_n1287));
  AOI211_X1 g1087(.A(G384), .B(new_n1249), .C1(new_n1279), .C2(new_n1280), .ZN(new_n1288));
  INV_X1    g1088(.A(G2897), .ZN(new_n1289));
  OAI22_X1  g1089(.A1(new_n1287), .A2(new_n1288), .B1(new_n1289), .B2(new_n1271), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1271), .A2(new_n1289), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1278), .A2(new_n1282), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1257), .B1(new_n1201), .B2(new_n1230), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1290), .B(new_n1292), .C1(new_n1293), .C2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(G375), .A2(G378), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1267), .A2(new_n1228), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(G378), .A2(new_n1297), .ZN(new_n1298));
  AOI22_X1  g1098(.A1(new_n1298), .A2(new_n1269), .B1(G213), .B2(new_n677), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT62), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1296), .A2(new_n1299), .A3(new_n1300), .A4(new_n1283), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1285), .A2(new_n1286), .A3(new_n1295), .A4(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1261), .B1(new_n1021), .B2(new_n1057), .ZN(new_n1303));
  OAI21_X1  g1103(.A(KEYINPUT127), .B1(new_n1263), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1303), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT127), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1305), .A2(new_n1306), .A3(new_n1262), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1304), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n983), .A2(new_n1014), .A3(G390), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(G390), .B1(new_n983), .B2(new_n1014), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1308), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(G387), .A2(new_n1259), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1313), .A2(new_n1304), .A3(new_n1307), .A4(new_n1309), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1312), .A2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1302), .A2(new_n1316), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1278), .A2(new_n1282), .A3(new_n1291), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1291), .B1(new_n1278), .B2(new_n1282), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(KEYINPUT61), .B1(new_n1320), .B2(new_n1272), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1296), .A2(new_n1299), .A3(KEYINPUT63), .A4(new_n1283), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT63), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1323), .B1(new_n1272), .B2(new_n1284), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1321), .A2(new_n1322), .A3(new_n1315), .A4(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1317), .A2(new_n1325), .ZN(G405));
  XNOR2_X1  g1126(.A(new_n1315), .B(new_n1283), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1296), .A2(new_n1258), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(new_n1327), .B(new_n1328), .ZN(G402));
endmodule


