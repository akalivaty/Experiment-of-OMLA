

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U553 ( .A1(n737), .A2(n736), .ZN(n754) );
  NOR2_X4 U554 ( .A1(G2105), .A2(n533), .ZN(n882) );
  NOR2_X2 U555 ( .A1(n793), .A2(n693), .ZN(n721) );
  BUF_X1 U556 ( .A(n619), .Z(n620) );
  AND2_X2 U557 ( .A1(G2104), .A2(G2105), .ZN(n887) );
  NAND2_X1 U558 ( .A1(n714), .A2(n713), .ZN(n716) );
  AND2_X1 U559 ( .A1(n519), .A2(n810), .ZN(n518) );
  XOR2_X1 U560 ( .A(n809), .B(KEYINPUT100), .Z(n519) );
  OR2_X1 U561 ( .A1(n771), .A2(n770), .ZN(n520) );
  AND2_X1 U562 ( .A1(n774), .A2(n773), .ZN(n521) );
  INV_X1 U563 ( .A(KEYINPUT104), .ZN(n715) );
  AND2_X1 U564 ( .A1(n772), .A2(n520), .ZN(n773) );
  NOR2_X2 U565 ( .A1(G2104), .A2(n524), .ZN(n619) );
  NOR2_X1 U566 ( .A1(G651), .A2(n648), .ZN(n651) );
  NOR2_X1 U567 ( .A1(n536), .A2(n535), .ZN(G160) );
  INV_X1 U568 ( .A(KEYINPUT66), .ZN(n523) );
  NAND2_X1 U569 ( .A1(G113), .A2(n887), .ZN(n522) );
  XNOR2_X1 U570 ( .A(n523), .B(n522), .ZN(n527) );
  INV_X1 U571 ( .A(G2105), .ZN(n524) );
  NAND2_X1 U572 ( .A1(G125), .A2(n619), .ZN(n525) );
  XNOR2_X1 U573 ( .A(KEYINPUT65), .B(n525), .ZN(n526) );
  NOR2_X1 U574 ( .A1(n527), .A2(n526), .ZN(n532) );
  XNOR2_X1 U575 ( .A(KEYINPUT68), .B(KEYINPUT17), .ZN(n529) );
  NOR2_X1 U576 ( .A1(G2104), .A2(G2105), .ZN(n528) );
  XNOR2_X1 U577 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U578 ( .A(KEYINPUT67), .B(n530), .ZN(n625) );
  NAND2_X1 U579 ( .A1(G137), .A2(n625), .ZN(n531) );
  NAND2_X1 U580 ( .A1(n532), .A2(n531), .ZN(n536) );
  INV_X1 U581 ( .A(G2104), .ZN(n533) );
  NAND2_X1 U582 ( .A1(G101), .A2(n882), .ZN(n534) );
  XNOR2_X1 U583 ( .A(KEYINPUT23), .B(n534), .ZN(n535) );
  NOR2_X1 U584 ( .A1(G543), .A2(G651), .ZN(n653) );
  NAND2_X1 U585 ( .A1(G85), .A2(n653), .ZN(n538) );
  XOR2_X1 U586 ( .A(G543), .B(KEYINPUT0), .Z(n648) );
  INV_X1 U587 ( .A(G651), .ZN(n539) );
  NOR2_X1 U588 ( .A1(n648), .A2(n539), .ZN(n657) );
  NAND2_X1 U589 ( .A1(G72), .A2(n657), .ZN(n537) );
  NAND2_X1 U590 ( .A1(n538), .A2(n537), .ZN(n545) );
  NAND2_X1 U591 ( .A1(G47), .A2(n651), .ZN(n543) );
  NOR2_X1 U592 ( .A1(G543), .A2(n539), .ZN(n541) );
  XNOR2_X1 U593 ( .A(KEYINPUT1), .B(KEYINPUT69), .ZN(n540) );
  XNOR2_X1 U594 ( .A(n541), .B(n540), .ZN(n654) );
  NAND2_X1 U595 ( .A1(G60), .A2(n654), .ZN(n542) );
  NAND2_X1 U596 ( .A1(n543), .A2(n542), .ZN(n544) );
  OR2_X1 U597 ( .A1(n545), .A2(n544), .ZN(G290) );
  NAND2_X1 U598 ( .A1(n625), .A2(G138), .ZN(n552) );
  NAND2_X1 U599 ( .A1(G102), .A2(n882), .ZN(n547) );
  NAND2_X1 U600 ( .A1(G126), .A2(n619), .ZN(n546) );
  AND2_X1 U601 ( .A1(n547), .A2(n546), .ZN(n550) );
  NAND2_X1 U602 ( .A1(G114), .A2(n887), .ZN(n548) );
  XOR2_X1 U603 ( .A(KEYINPUT91), .B(n548), .Z(n549) );
  AND2_X1 U604 ( .A1(n550), .A2(n549), .ZN(n551) );
  AND2_X1 U605 ( .A1(n552), .A2(n551), .ZN(G164) );
  NAND2_X1 U606 ( .A1(n654), .A2(G64), .ZN(n553) );
  XNOR2_X1 U607 ( .A(n553), .B(KEYINPUT70), .ZN(n555) );
  NAND2_X1 U608 ( .A1(G52), .A2(n651), .ZN(n554) );
  NAND2_X1 U609 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U610 ( .A(KEYINPUT71), .B(n556), .Z(n564) );
  NAND2_X1 U611 ( .A1(n657), .A2(G77), .ZN(n557) );
  XNOR2_X1 U612 ( .A(KEYINPUT73), .B(n557), .ZN(n560) );
  NAND2_X1 U613 ( .A1(n653), .A2(G90), .ZN(n558) );
  XOR2_X1 U614 ( .A(n558), .B(KEYINPUT72), .Z(n559) );
  NOR2_X1 U615 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U616 ( .A(KEYINPUT74), .B(n561), .Z(n562) );
  XOR2_X1 U617 ( .A(KEYINPUT9), .B(n562), .Z(n563) );
  NOR2_X1 U618 ( .A1(n564), .A2(n563), .ZN(G171) );
  INV_X1 U619 ( .A(G171), .ZN(G301) );
  AND2_X1 U620 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U621 ( .A(G57), .ZN(G237) );
  INV_X1 U622 ( .A(G69), .ZN(G235) );
  INV_X1 U623 ( .A(G108), .ZN(G238) );
  INV_X1 U624 ( .A(G120), .ZN(G236) );
  NAND2_X1 U625 ( .A1(G51), .A2(n651), .ZN(n566) );
  NAND2_X1 U626 ( .A1(G63), .A2(n654), .ZN(n565) );
  NAND2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U628 ( .A(KEYINPUT6), .B(n567), .ZN(n575) );
  NAND2_X1 U629 ( .A1(G89), .A2(n653), .ZN(n568) );
  XNOR2_X1 U630 ( .A(n568), .B(KEYINPUT82), .ZN(n569) );
  XNOR2_X1 U631 ( .A(KEYINPUT4), .B(n569), .ZN(n572) );
  NAND2_X1 U632 ( .A1(n657), .A2(G76), .ZN(n570) );
  XOR2_X1 U633 ( .A(KEYINPUT83), .B(n570), .Z(n571) );
  NAND2_X1 U634 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U635 ( .A(n573), .B(KEYINPUT5), .Z(n574) );
  NOR2_X1 U636 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U637 ( .A(KEYINPUT84), .B(n576), .Z(n577) );
  XNOR2_X1 U638 ( .A(KEYINPUT7), .B(n577), .ZN(G168) );
  XOR2_X1 U639 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  XOR2_X1 U640 ( .A(KEYINPUT10), .B(KEYINPUT79), .Z(n579) );
  NAND2_X1 U641 ( .A1(G7), .A2(G661), .ZN(n578) );
  XOR2_X1 U642 ( .A(n579), .B(n578), .Z(n920) );
  NAND2_X1 U643 ( .A1(n920), .A2(G567), .ZN(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT11), .B(n580), .Z(G234) );
  NAND2_X1 U645 ( .A1(n653), .A2(G81), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(KEYINPUT12), .ZN(n583) );
  NAND2_X1 U647 ( .A1(G68), .A2(n657), .ZN(n582) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(KEYINPUT13), .ZN(n586) );
  NAND2_X1 U650 ( .A1(G43), .A2(n651), .ZN(n585) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U652 ( .A1(n654), .A2(G56), .ZN(n587) );
  XOR2_X1 U653 ( .A(KEYINPUT14), .B(n587), .Z(n588) );
  NOR2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n979) );
  NAND2_X1 U655 ( .A1(n979), .A2(G860), .ZN(G153) );
  NAND2_X1 U656 ( .A1(G301), .A2(G868), .ZN(n590) );
  XNOR2_X1 U657 ( .A(n590), .B(KEYINPUT80), .ZN(n600) );
  INV_X1 U658 ( .A(G868), .ZN(n674) );
  NAND2_X1 U659 ( .A1(G92), .A2(n653), .ZN(n592) );
  NAND2_X1 U660 ( .A1(G79), .A2(n657), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U662 ( .A1(G54), .A2(n651), .ZN(n594) );
  NAND2_X1 U663 ( .A1(G66), .A2(n654), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U665 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U666 ( .A(KEYINPUT15), .B(n597), .Z(n598) );
  XOR2_X1 U667 ( .A(KEYINPUT81), .B(n598), .Z(n899) );
  INV_X1 U668 ( .A(n899), .ZN(n980) );
  NAND2_X1 U669 ( .A1(n674), .A2(n980), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n600), .A2(n599), .ZN(G284) );
  NAND2_X1 U671 ( .A1(n653), .A2(G91), .ZN(n601) );
  XOR2_X1 U672 ( .A(KEYINPUT75), .B(n601), .Z(n603) );
  NAND2_X1 U673 ( .A1(n657), .A2(G78), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U675 ( .A(KEYINPUT76), .B(n604), .Z(n610) );
  NAND2_X1 U676 ( .A1(n654), .A2(G65), .ZN(n605) );
  XOR2_X1 U677 ( .A(KEYINPUT77), .B(n605), .Z(n607) );
  NAND2_X1 U678 ( .A1(n651), .A2(G53), .ZN(n606) );
  NAND2_X1 U679 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U680 ( .A(KEYINPUT78), .B(n608), .Z(n609) );
  NAND2_X1 U681 ( .A1(n610), .A2(n609), .ZN(G299) );
  NAND2_X1 U682 ( .A1(G868), .A2(G286), .ZN(n612) );
  NAND2_X1 U683 ( .A1(G299), .A2(n674), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n612), .A2(n611), .ZN(G297) );
  INV_X1 U685 ( .A(G860), .ZN(n613) );
  NAND2_X1 U686 ( .A1(n613), .A2(G559), .ZN(n614) );
  NAND2_X1 U687 ( .A1(n614), .A2(n899), .ZN(n615) );
  XNOR2_X1 U688 ( .A(n615), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U689 ( .A1(n899), .A2(G868), .ZN(n616) );
  NOR2_X1 U690 ( .A1(G559), .A2(n616), .ZN(n618) );
  AND2_X1 U691 ( .A1(n674), .A2(n979), .ZN(n617) );
  NOR2_X1 U692 ( .A1(n618), .A2(n617), .ZN(G282) );
  NAND2_X1 U693 ( .A1(G123), .A2(n620), .ZN(n621) );
  XOR2_X1 U694 ( .A(KEYINPUT85), .B(n621), .Z(n622) );
  XNOR2_X1 U695 ( .A(n622), .B(KEYINPUT18), .ZN(n624) );
  NAND2_X1 U696 ( .A1(G111), .A2(n887), .ZN(n623) );
  NAND2_X1 U697 ( .A1(n624), .A2(n623), .ZN(n629) );
  NAND2_X1 U698 ( .A1(n882), .A2(G99), .ZN(n627) );
  BUF_X1 U699 ( .A(n625), .Z(n883) );
  NAND2_X1 U700 ( .A1(G135), .A2(n883), .ZN(n626) );
  NAND2_X1 U701 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U702 ( .A1(n629), .A2(n628), .ZN(n1004) );
  XNOR2_X1 U703 ( .A(G2096), .B(n1004), .ZN(n630) );
  INV_X1 U704 ( .A(G2100), .ZN(n850) );
  NAND2_X1 U705 ( .A1(n630), .A2(n850), .ZN(G156) );
  NAND2_X1 U706 ( .A1(G93), .A2(n653), .ZN(n632) );
  NAND2_X1 U707 ( .A1(G80), .A2(n657), .ZN(n631) );
  NAND2_X1 U708 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U709 ( .A1(G55), .A2(n651), .ZN(n634) );
  NAND2_X1 U710 ( .A1(G67), .A2(n654), .ZN(n633) );
  NAND2_X1 U711 ( .A1(n634), .A2(n633), .ZN(n635) );
  OR2_X1 U712 ( .A1(n636), .A2(n635), .ZN(n673) );
  NAND2_X1 U713 ( .A1(n899), .A2(G559), .ZN(n669) );
  XOR2_X1 U714 ( .A(n979), .B(n669), .Z(n637) );
  NOR2_X1 U715 ( .A1(G860), .A2(n637), .ZN(n638) );
  XOR2_X1 U716 ( .A(n673), .B(n638), .Z(G145) );
  NAND2_X1 U717 ( .A1(G88), .A2(n653), .ZN(n640) );
  NAND2_X1 U718 ( .A1(G75), .A2(n657), .ZN(n639) );
  NAND2_X1 U719 ( .A1(n640), .A2(n639), .ZN(n644) );
  NAND2_X1 U720 ( .A1(G50), .A2(n651), .ZN(n642) );
  NAND2_X1 U721 ( .A1(G62), .A2(n654), .ZN(n641) );
  NAND2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U723 ( .A1(n644), .A2(n643), .ZN(G166) );
  INV_X1 U724 ( .A(G166), .ZN(G303) );
  NAND2_X1 U725 ( .A1(G49), .A2(n651), .ZN(n646) );
  NAND2_X1 U726 ( .A1(G74), .A2(G651), .ZN(n645) );
  NAND2_X1 U727 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U728 ( .A1(n654), .A2(n647), .ZN(n650) );
  NAND2_X1 U729 ( .A1(n648), .A2(G87), .ZN(n649) );
  NAND2_X1 U730 ( .A1(n650), .A2(n649), .ZN(G288) );
  NAND2_X1 U731 ( .A1(G48), .A2(n651), .ZN(n652) );
  XNOR2_X1 U732 ( .A(n652), .B(KEYINPUT86), .ZN(n662) );
  NAND2_X1 U733 ( .A1(G86), .A2(n653), .ZN(n656) );
  NAND2_X1 U734 ( .A1(G61), .A2(n654), .ZN(n655) );
  NAND2_X1 U735 ( .A1(n656), .A2(n655), .ZN(n660) );
  NAND2_X1 U736 ( .A1(n657), .A2(G73), .ZN(n658) );
  XOR2_X1 U737 ( .A(KEYINPUT2), .B(n658), .Z(n659) );
  NOR2_X1 U738 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U739 ( .A1(n662), .A2(n661), .ZN(G305) );
  XOR2_X1 U740 ( .A(G303), .B(G290), .Z(n668) );
  XOR2_X1 U741 ( .A(G299), .B(KEYINPUT19), .Z(n664) );
  XNOR2_X1 U742 ( .A(G288), .B(n979), .ZN(n663) );
  XNOR2_X1 U743 ( .A(n664), .B(n663), .ZN(n665) );
  XOR2_X1 U744 ( .A(n673), .B(n665), .Z(n666) );
  XNOR2_X1 U745 ( .A(n666), .B(G305), .ZN(n667) );
  XNOR2_X1 U746 ( .A(n668), .B(n667), .ZN(n898) );
  XNOR2_X1 U747 ( .A(n898), .B(KEYINPUT87), .ZN(n670) );
  XNOR2_X1 U748 ( .A(n670), .B(n669), .ZN(n671) );
  NAND2_X1 U749 ( .A1(n671), .A2(G868), .ZN(n672) );
  XNOR2_X1 U750 ( .A(n672), .B(KEYINPUT88), .ZN(n676) );
  NAND2_X1 U751 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U752 ( .A1(n676), .A2(n675), .ZN(G295) );
  NAND2_X1 U753 ( .A1(G2078), .A2(G2084), .ZN(n677) );
  XOR2_X1 U754 ( .A(KEYINPUT20), .B(n677), .Z(n678) );
  NAND2_X1 U755 ( .A1(G2090), .A2(n678), .ZN(n679) );
  XNOR2_X1 U756 ( .A(KEYINPUT21), .B(n679), .ZN(n680) );
  NAND2_X1 U757 ( .A1(n680), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U758 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U759 ( .A(KEYINPUT89), .B(KEYINPUT22), .Z(n682) );
  NAND2_X1 U760 ( .A1(G132), .A2(G82), .ZN(n681) );
  XNOR2_X1 U761 ( .A(n682), .B(n681), .ZN(n683) );
  NOR2_X1 U762 ( .A1(n683), .A2(G218), .ZN(n684) );
  NAND2_X1 U763 ( .A1(G96), .A2(n684), .ZN(n831) );
  NAND2_X1 U764 ( .A1(G2106), .A2(n831), .ZN(n689) );
  NOR2_X1 U765 ( .A1(G236), .A2(G238), .ZN(n686) );
  NOR2_X1 U766 ( .A1(G235), .A2(G237), .ZN(n685) );
  NAND2_X1 U767 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U768 ( .A(KEYINPUT90), .B(n687), .ZN(n832) );
  NAND2_X1 U769 ( .A1(n832), .A2(G567), .ZN(n688) );
  NAND2_X1 U770 ( .A1(n689), .A2(n688), .ZN(n833) );
  NAND2_X1 U771 ( .A1(G661), .A2(G483), .ZN(n690) );
  NOR2_X1 U772 ( .A1(n833), .A2(n690), .ZN(n830) );
  NAND2_X1 U773 ( .A1(n830), .A2(G36), .ZN(G176) );
  NOR2_X1 U774 ( .A1(G1976), .A2(G288), .ZN(n759) );
  NOR2_X1 U775 ( .A1(G1971), .A2(G303), .ZN(n691) );
  NOR2_X1 U776 ( .A1(n759), .A2(n691), .ZN(n976) );
  NAND2_X1 U777 ( .A1(G160), .A2(G40), .ZN(n793) );
  NOR2_X1 U778 ( .A1(G164), .A2(G1384), .ZN(n794) );
  INV_X1 U779 ( .A(n794), .ZN(n693) );
  INV_X1 U780 ( .A(n721), .ZN(n738) );
  NAND2_X1 U781 ( .A1(G1956), .A2(n738), .ZN(n694) );
  XNOR2_X1 U782 ( .A(KEYINPUT102), .B(n694), .ZN(n697) );
  NAND2_X1 U783 ( .A1(n721), .A2(G2072), .ZN(n695) );
  XOR2_X1 U784 ( .A(KEYINPUT27), .B(n695), .Z(n696) );
  NAND2_X1 U785 ( .A1(n697), .A2(n696), .ZN(n712) );
  NAND2_X1 U786 ( .A1(G299), .A2(n712), .ZN(n698) );
  XOR2_X1 U787 ( .A(KEYINPUT28), .B(n698), .Z(n718) );
  NAND2_X1 U788 ( .A1(n721), .A2(G1996), .ZN(n699) );
  XNOR2_X1 U789 ( .A(n699), .B(KEYINPUT26), .ZN(n701) );
  NAND2_X1 U790 ( .A1(G1341), .A2(n738), .ZN(n700) );
  NAND2_X1 U791 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U792 ( .A(n702), .B(KEYINPUT103), .ZN(n703) );
  NAND2_X1 U793 ( .A1(n703), .A2(n979), .ZN(n704) );
  XNOR2_X1 U794 ( .A(KEYINPUT64), .B(n704), .ZN(n709) );
  OR2_X1 U795 ( .A1(n980), .A2(n709), .ZN(n708) );
  NOR2_X1 U796 ( .A1(n721), .A2(G1348), .ZN(n706) );
  NOR2_X1 U797 ( .A1(G2067), .A2(n738), .ZN(n705) );
  NOR2_X1 U798 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U799 ( .A1(n708), .A2(n707), .ZN(n711) );
  NAND2_X1 U800 ( .A1(n709), .A2(n980), .ZN(n710) );
  NAND2_X1 U801 ( .A1(n711), .A2(n710), .ZN(n714) );
  OR2_X1 U802 ( .A1(G299), .A2(n712), .ZN(n713) );
  XNOR2_X1 U803 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X1 U804 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U805 ( .A(n719), .B(KEYINPUT29), .ZN(n725) );
  NOR2_X1 U806 ( .A1(n721), .A2(G1961), .ZN(n720) );
  XNOR2_X1 U807 ( .A(n720), .B(KEYINPUT101), .ZN(n723) );
  XNOR2_X1 U808 ( .A(KEYINPUT25), .B(G2078), .ZN(n951) );
  NAND2_X1 U809 ( .A1(n721), .A2(n951), .ZN(n722) );
  NAND2_X1 U810 ( .A1(n723), .A2(n722), .ZN(n729) );
  NAND2_X1 U811 ( .A1(G171), .A2(n729), .ZN(n724) );
  NAND2_X1 U812 ( .A1(n725), .A2(n724), .ZN(n747) );
  NAND2_X1 U813 ( .A1(G8), .A2(n738), .ZN(n771) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n771), .ZN(n734) );
  NOR2_X1 U815 ( .A1(G2084), .A2(n738), .ZN(n733) );
  NOR2_X1 U816 ( .A1(n734), .A2(n733), .ZN(n726) );
  NAND2_X1 U817 ( .A1(G8), .A2(n726), .ZN(n727) );
  XNOR2_X1 U818 ( .A(KEYINPUT30), .B(n727), .ZN(n728) );
  NOR2_X1 U819 ( .A1(G168), .A2(n728), .ZN(n731) );
  NOR2_X1 U820 ( .A1(G171), .A2(n729), .ZN(n730) );
  NOR2_X1 U821 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U822 ( .A(KEYINPUT31), .B(n732), .Z(n745) );
  AND2_X1 U823 ( .A1(n747), .A2(n745), .ZN(n737) );
  AND2_X1 U824 ( .A1(G8), .A2(n733), .ZN(n735) );
  OR2_X1 U825 ( .A1(n735), .A2(n734), .ZN(n736) );
  INV_X1 U826 ( .A(G8), .ZN(n744) );
  NOR2_X1 U827 ( .A1(G2090), .A2(n738), .ZN(n739) );
  XNOR2_X1 U828 ( .A(KEYINPUT105), .B(n739), .ZN(n742) );
  NOR2_X1 U829 ( .A1(G1971), .A2(n771), .ZN(n740) );
  NOR2_X1 U830 ( .A1(G166), .A2(n740), .ZN(n741) );
  NAND2_X1 U831 ( .A1(n742), .A2(n741), .ZN(n743) );
  OR2_X1 U832 ( .A1(n744), .A2(n743), .ZN(n748) );
  AND2_X1 U833 ( .A1(n745), .A2(n748), .ZN(n746) );
  NAND2_X1 U834 ( .A1(n747), .A2(n746), .ZN(n751) );
  INV_X1 U835 ( .A(n748), .ZN(n749) );
  OR2_X1 U836 ( .A1(n749), .A2(G286), .ZN(n750) );
  NAND2_X1 U837 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U838 ( .A(n752), .B(KEYINPUT32), .ZN(n753) );
  NAND2_X1 U839 ( .A1(n754), .A2(n753), .ZN(n766) );
  AND2_X1 U840 ( .A1(n976), .A2(n766), .ZN(n757) );
  NAND2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n975) );
  INV_X1 U842 ( .A(n771), .ZN(n755) );
  NAND2_X1 U843 ( .A1(n975), .A2(n755), .ZN(n756) );
  NOR2_X1 U844 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X1 U845 ( .A1(n758), .A2(KEYINPUT33), .ZN(n762) );
  NAND2_X1 U846 ( .A1(n759), .A2(KEYINPUT33), .ZN(n760) );
  NOR2_X1 U847 ( .A1(n760), .A2(n771), .ZN(n761) );
  NOR2_X1 U848 ( .A1(n762), .A2(n761), .ZN(n763) );
  XOR2_X1 U849 ( .A(G1981), .B(G305), .Z(n971) );
  NAND2_X1 U850 ( .A1(n763), .A2(n971), .ZN(n774) );
  NOR2_X1 U851 ( .A1(G2090), .A2(G303), .ZN(n764) );
  NAND2_X1 U852 ( .A1(G8), .A2(n764), .ZN(n765) );
  NAND2_X1 U853 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U854 ( .A1(n771), .A2(n767), .ZN(n768) );
  XNOR2_X1 U855 ( .A(n768), .B(KEYINPUT106), .ZN(n772) );
  NOR2_X1 U856 ( .A1(G1981), .A2(G305), .ZN(n769) );
  XOR2_X1 U857 ( .A(n769), .B(KEYINPUT24), .Z(n770) );
  XNOR2_X1 U858 ( .A(n521), .B(KEYINPUT107), .ZN(n811) );
  XNOR2_X1 U859 ( .A(KEYINPUT98), .B(G1991), .ZN(n950) );
  NAND2_X1 U860 ( .A1(G107), .A2(n887), .ZN(n775) );
  XNOR2_X1 U861 ( .A(n775), .B(KEYINPUT96), .ZN(n782) );
  NAND2_X1 U862 ( .A1(G95), .A2(n882), .ZN(n777) );
  NAND2_X1 U863 ( .A1(G119), .A2(n620), .ZN(n776) );
  NAND2_X1 U864 ( .A1(n777), .A2(n776), .ZN(n780) );
  NAND2_X1 U865 ( .A1(G131), .A2(n883), .ZN(n778) );
  XNOR2_X1 U866 ( .A(KEYINPUT97), .B(n778), .ZN(n779) );
  NOR2_X1 U867 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U868 ( .A1(n782), .A2(n781), .ZN(n869) );
  AND2_X1 U869 ( .A1(n950), .A2(n869), .ZN(n792) );
  NAND2_X1 U870 ( .A1(G105), .A2(n882), .ZN(n783) );
  XOR2_X1 U871 ( .A(KEYINPUT38), .B(n783), .Z(n788) );
  NAND2_X1 U872 ( .A1(G117), .A2(n887), .ZN(n785) );
  NAND2_X1 U873 ( .A1(G129), .A2(n620), .ZN(n784) );
  NAND2_X1 U874 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U875 ( .A(KEYINPUT99), .B(n786), .Z(n787) );
  NOR2_X1 U876 ( .A1(n788), .A2(n787), .ZN(n790) );
  NAND2_X1 U877 ( .A1(G141), .A2(n883), .ZN(n789) );
  NAND2_X1 U878 ( .A1(n790), .A2(n789), .ZN(n862) );
  AND2_X1 U879 ( .A1(n862), .A2(G1996), .ZN(n791) );
  NOR2_X1 U880 ( .A1(n792), .A2(n791), .ZN(n1001) );
  INV_X1 U881 ( .A(n1001), .ZN(n795) );
  NOR2_X1 U882 ( .A1(n794), .A2(n793), .ZN(n823) );
  NAND2_X1 U883 ( .A1(n795), .A2(n823), .ZN(n812) );
  XOR2_X1 U884 ( .A(G2067), .B(KEYINPUT37), .Z(n796) );
  XOR2_X1 U885 ( .A(KEYINPUT92), .B(n796), .Z(n821) );
  NAND2_X1 U886 ( .A1(G116), .A2(n887), .ZN(n798) );
  NAND2_X1 U887 ( .A1(G128), .A2(n620), .ZN(n797) );
  NAND2_X1 U888 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U889 ( .A(KEYINPUT35), .B(n799), .ZN(n806) );
  XNOR2_X1 U890 ( .A(KEYINPUT94), .B(KEYINPUT34), .ZN(n804) );
  NAND2_X1 U891 ( .A1(G140), .A2(n883), .ZN(n802) );
  NAND2_X1 U892 ( .A1(n882), .A2(G104), .ZN(n800) );
  XOR2_X1 U893 ( .A(KEYINPUT93), .B(n800), .Z(n801) );
  NAND2_X1 U894 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U895 ( .A(n804), .B(n803), .Z(n805) );
  NAND2_X1 U896 ( .A1(n806), .A2(n805), .ZN(n807) );
  XOR2_X1 U897 ( .A(KEYINPUT36), .B(n807), .Z(n894) );
  OR2_X1 U898 ( .A1(n821), .A2(n894), .ZN(n808) );
  XNOR2_X1 U899 ( .A(n808), .B(KEYINPUT95), .ZN(n1017) );
  NAND2_X1 U900 ( .A1(n823), .A2(n1017), .ZN(n819) );
  NAND2_X1 U901 ( .A1(n812), .A2(n819), .ZN(n809) );
  XNOR2_X1 U902 ( .A(G1986), .B(G290), .ZN(n978) );
  NAND2_X1 U903 ( .A1(n978), .A2(n823), .ZN(n810) );
  NAND2_X1 U904 ( .A1(n811), .A2(n518), .ZN(n826) );
  NOR2_X1 U905 ( .A1(G1996), .A2(n862), .ZN(n996) );
  INV_X1 U906 ( .A(n812), .ZN(n816) );
  NOR2_X1 U907 ( .A1(n950), .A2(n869), .ZN(n813) );
  XNOR2_X1 U908 ( .A(KEYINPUT108), .B(n813), .ZN(n1000) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n814) );
  NOR2_X1 U910 ( .A1(n1000), .A2(n814), .ZN(n815) );
  NOR2_X1 U911 ( .A1(n816), .A2(n815), .ZN(n817) );
  NOR2_X1 U912 ( .A1(n996), .A2(n817), .ZN(n818) );
  XNOR2_X1 U913 ( .A(n818), .B(KEYINPUT39), .ZN(n820) );
  NAND2_X1 U914 ( .A1(n820), .A2(n819), .ZN(n822) );
  NAND2_X1 U915 ( .A1(n821), .A2(n894), .ZN(n1005) );
  NAND2_X1 U916 ( .A1(n822), .A2(n1005), .ZN(n824) );
  NAND2_X1 U917 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U918 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U919 ( .A(n827), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n920), .ZN(G217) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n828) );
  NAND2_X1 U922 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U924 ( .A1(n830), .A2(n829), .ZN(G188) );
  INV_X1 U926 ( .A(G132), .ZN(G219) );
  INV_X1 U927 ( .A(G96), .ZN(G221) );
  INV_X1 U928 ( .A(G82), .ZN(G220) );
  NOR2_X1 U929 ( .A1(n832), .A2(n831), .ZN(G325) );
  INV_X1 U930 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U931 ( .A(KEYINPUT111), .B(n833), .ZN(G319) );
  XOR2_X1 U932 ( .A(KEYINPUT41), .B(G1986), .Z(n835) );
  XNOR2_X1 U933 ( .A(G1996), .B(G1991), .ZN(n834) );
  XNOR2_X1 U934 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U935 ( .A(n836), .B(G2474), .Z(n838) );
  XNOR2_X1 U936 ( .A(G1981), .B(G1966), .ZN(n837) );
  XNOR2_X1 U937 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U938 ( .A(G1956), .B(G1961), .Z(n840) );
  XNOR2_X1 U939 ( .A(G1976), .B(G1971), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U941 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U942 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(G229) );
  XOR2_X1 U944 ( .A(G2096), .B(KEYINPUT43), .Z(n846) );
  XNOR2_X1 U945 ( .A(G2090), .B(G2678), .ZN(n845) );
  XNOR2_X1 U946 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U947 ( .A(n847), .B(KEYINPUT112), .Z(n849) );
  XNOR2_X1 U948 ( .A(G2067), .B(G2072), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n854) );
  XNOR2_X1 U950 ( .A(KEYINPUT42), .B(n850), .ZN(n852) );
  XNOR2_X1 U951 ( .A(G2078), .B(G2084), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n854), .B(n853), .ZN(G227) );
  NAND2_X1 U954 ( .A1(G124), .A2(n620), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n855), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U956 ( .A1(n887), .A2(G112), .ZN(n856) );
  NAND2_X1 U957 ( .A1(n857), .A2(n856), .ZN(n861) );
  NAND2_X1 U958 ( .A1(n882), .A2(G100), .ZN(n859) );
  NAND2_X1 U959 ( .A1(G136), .A2(n883), .ZN(n858) );
  NAND2_X1 U960 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U961 ( .A1(n861), .A2(n860), .ZN(G162) );
  XNOR2_X1 U962 ( .A(G162), .B(n862), .ZN(n864) );
  XNOR2_X1 U963 ( .A(G164), .B(G160), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(n868) );
  XOR2_X1 U965 ( .A(KEYINPUT119), .B(KEYINPUT118), .Z(n866) );
  XNOR2_X1 U966 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n865) );
  XNOR2_X1 U967 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U968 ( .A(n868), .B(n867), .Z(n871) );
  XOR2_X1 U969 ( .A(n869), .B(n1004), .Z(n870) );
  XNOR2_X1 U970 ( .A(n871), .B(n870), .ZN(n881) );
  NAND2_X1 U971 ( .A1(n882), .A2(G106), .ZN(n873) );
  NAND2_X1 U972 ( .A1(G142), .A2(n883), .ZN(n872) );
  NAND2_X1 U973 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U974 ( .A(n874), .B(KEYINPUT45), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G118), .A2(n887), .ZN(n875) );
  NAND2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n879) );
  NAND2_X1 U977 ( .A1(G130), .A2(n620), .ZN(n877) );
  XNOR2_X1 U978 ( .A(KEYINPUT115), .B(n877), .ZN(n878) );
  NOR2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U980 ( .A(n881), .B(n880), .Z(n896) );
  NAND2_X1 U981 ( .A1(n882), .A2(G103), .ZN(n885) );
  NAND2_X1 U982 ( .A1(G139), .A2(n883), .ZN(n884) );
  NAND2_X1 U983 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U984 ( .A(KEYINPUT116), .B(n886), .ZN(n893) );
  NAND2_X1 U985 ( .A1(G115), .A2(n887), .ZN(n889) );
  NAND2_X1 U986 ( .A1(G127), .A2(n620), .ZN(n888) );
  NAND2_X1 U987 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U988 ( .A(KEYINPUT47), .B(n890), .ZN(n891) );
  XNOR2_X1 U989 ( .A(KEYINPUT117), .B(n891), .ZN(n892) );
  NOR2_X1 U990 ( .A1(n893), .A2(n892), .ZN(n1007) );
  XOR2_X1 U991 ( .A(n894), .B(n1007), .Z(n895) );
  XNOR2_X1 U992 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U993 ( .A1(G37), .A2(n897), .ZN(G395) );
  XNOR2_X1 U994 ( .A(G286), .B(n898), .ZN(n901) );
  XOR2_X1 U995 ( .A(G301), .B(n899), .Z(n900) );
  XNOR2_X1 U996 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U997 ( .A1(G37), .A2(n902), .ZN(G397) );
  XNOR2_X1 U998 ( .A(G2446), .B(G2443), .ZN(n912) );
  XOR2_X1 U999 ( .A(G2430), .B(KEYINPUT110), .Z(n904) );
  XNOR2_X1 U1000 ( .A(G2454), .B(G2435), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n908) );
  XOR2_X1 U1002 ( .A(G2438), .B(G2427), .Z(n906) );
  XNOR2_X1 U1003 ( .A(G1348), .B(G1341), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1005 ( .A(n908), .B(n907), .Z(n910) );
  XNOR2_X1 U1006 ( .A(KEYINPUT109), .B(G2451), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(n912), .B(n911), .ZN(n913) );
  NAND2_X1 U1009 ( .A1(n913), .A2(G14), .ZN(n919) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n919), .ZN(n916) );
  NOR2_X1 U1011 ( .A1(G229), .A2(G227), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n914), .ZN(n915) );
  NOR2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(n919), .ZN(G401) );
  INV_X1 U1018 ( .A(n920), .ZN(G223) );
  XNOR2_X1 U1019 ( .A(G1966), .B(G21), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(G5), .B(G1961), .ZN(n921) );
  NOR2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n933) );
  XNOR2_X1 U1022 ( .A(KEYINPUT59), .B(KEYINPUT125), .ZN(n923) );
  XNOR2_X1 U1023 ( .A(n923), .B(G4), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(G1348), .B(n924), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(G1956), .B(G20), .ZN(n925) );
  NOR2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n930) );
  XNOR2_X1 U1027 ( .A(G1981), .B(G6), .ZN(n928) );
  XNOR2_X1 U1028 ( .A(G19), .B(G1341), .ZN(n927) );
  NOR2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1031 ( .A(KEYINPUT60), .B(n931), .Z(n932) );
  NAND2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n941) );
  XNOR2_X1 U1033 ( .A(G1976), .B(G23), .ZN(n935) );
  XNOR2_X1 U1034 ( .A(G1971), .B(G22), .ZN(n934) );
  NOR2_X1 U1035 ( .A1(n935), .A2(n934), .ZN(n938) );
  XOR2_X1 U1036 ( .A(G1986), .B(KEYINPUT126), .Z(n936) );
  XNOR2_X1 U1037 ( .A(G24), .B(n936), .ZN(n937) );
  NAND2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1039 ( .A(KEYINPUT58), .B(n939), .ZN(n940) );
  NOR2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1041 ( .A(KEYINPUT61), .B(n942), .Z(n943) );
  NOR2_X1 U1042 ( .A1(G16), .A2(n943), .ZN(n944) );
  XOR2_X1 U1043 ( .A(KEYINPUT127), .B(n944), .Z(n1025) );
  XOR2_X1 U1044 ( .A(G34), .B(KEYINPUT122), .Z(n946) );
  XNOR2_X1 U1045 ( .A(G2084), .B(KEYINPUT54), .ZN(n945) );
  XNOR2_X1 U1046 ( .A(n946), .B(n945), .ZN(n962) );
  XNOR2_X1 U1047 ( .A(G2090), .B(G35), .ZN(n960) );
  XOR2_X1 U1048 ( .A(G32), .B(G1996), .Z(n947) );
  NAND2_X1 U1049 ( .A1(n947), .A2(G28), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(G2067), .B(G26), .ZN(n949) );
  XNOR2_X1 U1051 ( .A(G33), .B(G2072), .ZN(n948) );
  NOR2_X1 U1052 ( .A1(n949), .A2(n948), .ZN(n955) );
  XNOR2_X1 U1053 ( .A(n950), .B(G25), .ZN(n953) );
  XOR2_X1 U1054 ( .A(n951), .B(G27), .Z(n952) );
  NOR2_X1 U1055 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1056 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1057 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1058 ( .A(KEYINPUT53), .B(n958), .ZN(n959) );
  NOR2_X1 U1059 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1061 ( .A(KEYINPUT55), .B(n963), .Z(n965) );
  INV_X1 U1062 ( .A(G29), .ZN(n964) );
  NAND2_X1 U1063 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1064 ( .A1(G11), .A2(n966), .ZN(n994) );
  XNOR2_X1 U1065 ( .A(G16), .B(KEYINPUT56), .ZN(n967) );
  XNOR2_X1 U1066 ( .A(n967), .B(KEYINPUT123), .ZN(n992) );
  XOR2_X1 U1067 ( .A(G299), .B(G1956), .Z(n969) );
  XOR2_X1 U1068 ( .A(G301), .B(G1961), .Z(n968) );
  NAND2_X1 U1069 ( .A1(n969), .A2(n968), .ZN(n990) );
  XNOR2_X1 U1070 ( .A(G1966), .B(KEYINPUT124), .ZN(n970) );
  XNOR2_X1 U1071 ( .A(n970), .B(G168), .ZN(n972) );
  NAND2_X1 U1072 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1073 ( .A(n973), .B(KEYINPUT57), .ZN(n988) );
  NAND2_X1 U1074 ( .A1(G1971), .A2(G303), .ZN(n974) );
  NAND2_X1 U1075 ( .A1(n975), .A2(n974), .ZN(n986) );
  INV_X1 U1076 ( .A(n976), .ZN(n977) );
  NOR2_X1 U1077 ( .A1(n978), .A2(n977), .ZN(n984) );
  XOR2_X1 U1078 ( .A(n979), .B(G1341), .Z(n982) );
  XNOR2_X1 U1079 ( .A(G1348), .B(n980), .ZN(n981) );
  NOR2_X1 U1080 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1081 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1082 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1084 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n1023) );
  XOR2_X1 U1087 ( .A(G2090), .B(G162), .Z(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1089 ( .A(KEYINPUT51), .B(n997), .Z(n998) );
  XOR2_X1 U1090 ( .A(KEYINPUT120), .B(n998), .Z(n999) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1015) );
  XNOR2_X1 U1092 ( .A(G160), .B(G2084), .ZN(n1002) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1013) );
  XOR2_X1 U1096 ( .A(n1007), .B(KEYINPUT121), .Z(n1008) );
  XOR2_X1 U1097 ( .A(G2072), .B(n1008), .Z(n1010) );
  XOR2_X1 U1098 ( .A(G164), .B(G2078), .Z(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1100 ( .A(KEYINPUT50), .B(n1011), .Z(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(KEYINPUT52), .B(n1018), .ZN(n1020) );
  INV_X1 U1105 ( .A(KEYINPUT55), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1107 ( .A1(n1021), .A2(G29), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1026), .Z(G150) );
  INV_X1 U1111 ( .A(G150), .ZN(G311) );
endmodule

