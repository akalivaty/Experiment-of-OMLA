//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 1 0 0 1 0 0 1 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015;
  INV_X1    g000(.A(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G214), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT18), .A2(G131), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G125), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G140), .ZN(new_n194));
  INV_X1    g008(.A(G140), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G125), .ZN(new_n196));
  NOR3_X1   g010(.A1(new_n194), .A2(new_n196), .A3(G146), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(KEYINPUT74), .A3(G125), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT74), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n199), .B1(new_n193), .B2(G140), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n198), .B1(new_n200), .B2(new_n194), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n197), .B1(G146), .B2(new_n201), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n192), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n190), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT67), .B(G131), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(KEYINPUT17), .A3(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n190), .B(new_n207), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n208), .B1(new_n210), .B2(KEYINPUT17), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n194), .A2(KEYINPUT16), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n212), .B1(new_n201), .B2(KEYINPUT16), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n213), .B(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n204), .B1(new_n211), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(G113), .B(G122), .ZN(new_n217));
  INV_X1    g031(.A(G104), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n217), .B(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n216), .B(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G902), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G475), .ZN(new_n224));
  NOR2_X1   g038(.A1(G475), .A2(G902), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n216), .A2(new_n220), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n201), .A2(KEYINPUT19), .ZN(new_n228));
  OR3_X1    g042(.A1(new_n194), .A2(new_n196), .A3(KEYINPUT19), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n228), .A2(new_n214), .A3(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT76), .B1(new_n213), .B2(new_n214), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT76), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT16), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n195), .A2(G125), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n234), .B1(new_n196), .B2(new_n199), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n233), .B1(new_n235), .B2(new_n198), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n232), .B(G146), .C1(new_n236), .C2(new_n212), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n230), .B1(new_n231), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT88), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n210), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AOI211_X1 g054(.A(KEYINPUT88), .B(new_n230), .C1(new_n231), .C2(new_n237), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n204), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n220), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n227), .B1(new_n243), .B2(KEYINPUT89), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT89), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n245), .A3(new_n220), .ZN(new_n246));
  AOI211_X1 g060(.A(KEYINPUT20), .B(new_n226), .C1(new_n244), .C2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT20), .ZN(new_n248));
  INV_X1    g062(.A(new_n230), .ZN(new_n249));
  INV_X1    g063(.A(new_n212), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n195), .A2(KEYINPUT74), .A3(G125), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n193), .A2(G140), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT74), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n251), .B1(new_n253), .B2(new_n234), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n250), .B1(new_n254), .B2(new_n233), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n232), .B1(new_n255), .B2(G146), .ZN(new_n256));
  NOR3_X1   g070(.A1(new_n213), .A2(KEYINPUT76), .A3(new_n214), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n249), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n209), .B1(new_n258), .B2(KEYINPUT88), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n238), .A2(new_n239), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n203), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT89), .B1(new_n261), .B2(new_n219), .ZN(new_n262));
  INV_X1    g076(.A(new_n227), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(new_n263), .A3(new_n246), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n248), .B1(new_n264), .B2(new_n225), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n224), .B1(new_n247), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G952), .ZN(new_n267));
  AOI211_X1 g081(.A(G953), .B(new_n267), .C1(G234), .C2(G237), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  XOR2_X1   g083(.A(KEYINPUT73), .B(G902), .Z(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  AOI211_X1 g085(.A(new_n188), .B(new_n271), .C1(G234), .C2(G237), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  XOR2_X1   g087(.A(KEYINPUT21), .B(G898), .Z(new_n274));
  OAI21_X1  g088(.A(new_n269), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  XOR2_X1   g089(.A(new_n275), .B(KEYINPUT97), .Z(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  XOR2_X1   g091(.A(KEYINPUT9), .B(G234), .Z(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(G217), .A3(new_n188), .ZN(new_n279));
  XNOR2_X1  g093(.A(G128), .B(G143), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT93), .B(G134), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n280), .B(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G122), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT90), .B1(new_n283), .B2(G116), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT90), .ZN(new_n285));
  INV_X1    g099(.A(G116), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n286), .A3(G122), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n283), .A2(G116), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT91), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT91), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n288), .A2(new_n292), .A3(new_n289), .ZN(new_n293));
  AOI21_X1  g107(.A(G107), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G107), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n288), .A2(KEYINPUT14), .B1(G116), .B2(new_n283), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT14), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n284), .A2(new_n287), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n295), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT94), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n294), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n300), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n282), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT95), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT92), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n288), .A2(new_n292), .A3(new_n289), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n292), .B1(new_n288), .B2(new_n289), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n307), .A2(new_n308), .A3(new_n295), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n306), .B1(new_n309), .B2(new_n294), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n295), .B1(new_n307), .B2(new_n308), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n291), .A2(G107), .A3(new_n293), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n312), .A3(KEYINPUT92), .ZN(new_n313));
  INV_X1    g127(.A(G128), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT13), .B1(new_n314), .B2(G143), .ZN(new_n315));
  INV_X1    g129(.A(G134), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(new_n280), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n310), .A2(new_n313), .A3(new_n318), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n304), .A2(new_n305), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n305), .B1(new_n304), .B2(new_n319), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n279), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n313), .A2(new_n318), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT92), .B1(new_n311), .B2(new_n312), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n282), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n296), .A2(new_n298), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G107), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(KEYINPUT94), .A3(new_n311), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n326), .B1(new_n329), .B2(new_n302), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT95), .B1(new_n325), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n279), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n304), .A2(new_n319), .A3(new_n305), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n322), .A2(new_n271), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G478), .ZN(new_n336));
  NOR2_X1   g150(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n336), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n340), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n322), .A2(new_n271), .A3(new_n334), .A4(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NOR3_X1   g158(.A1(new_n266), .A2(new_n277), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G110), .ZN(new_n346));
  INV_X1    g160(.A(G119), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G128), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n314), .A2(G119), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n349), .A2(KEYINPUT23), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT23), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n351), .B1(G119), .B2(new_n314), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n346), .B(new_n348), .C1(new_n350), .C2(new_n352), .ZN(new_n353));
  OR2_X1    g167(.A1(new_n353), .A2(KEYINPUT75), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n349), .A2(new_n348), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT24), .B(G110), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n353), .A2(KEYINPUT75), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n197), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n358), .B1(new_n256), .B2(new_n257), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n355), .A2(new_n356), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n348), .B1(new_n352), .B2(new_n350), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n360), .B1(new_n361), .B2(G110), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n215), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT22), .B(G137), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n366));
  XOR2_X1   g180(.A(new_n365), .B(new_n366), .Z(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n359), .A2(new_n363), .A3(new_n367), .ZN(new_n370));
  INV_X1    g184(.A(G217), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n371), .B1(new_n271), .B2(G234), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(G902), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n369), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT77), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n374), .B(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n372), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n369), .A2(new_n271), .A3(new_n370), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT25), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n369), .A2(KEYINPUT25), .A3(new_n271), .A4(new_n370), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n377), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT30), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT0), .ZN(new_n386));
  INV_X1    g200(.A(G143), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G146), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n214), .A2(G143), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n386), .B1(new_n390), .B2(new_n314), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT64), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n214), .A3(G143), .ZN(new_n393));
  AOI21_X1  g207(.A(KEYINPUT64), .B1(new_n387), .B2(G146), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n387), .A2(G146), .ZN(new_n395));
  OAI211_X1 g209(.A(G128), .B(new_n393), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n390), .A2(G128), .ZN(new_n397));
  AOI22_X1  g211(.A1(new_n391), .A2(new_n396), .B1(new_n397), .B2(new_n386), .ZN(new_n398));
  INV_X1    g212(.A(G137), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G134), .ZN(new_n400));
  AND2_X1   g214(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n401));
  NOR2_X1   g215(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT66), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n400), .B(KEYINPUT66), .C1(new_n401), .C2(new_n402), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n399), .A2(KEYINPUT11), .A3(G134), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n316), .A2(G137), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n405), .A2(new_n406), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G131), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n405), .A2(new_n406), .A3(new_n410), .A4(new_n206), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n398), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT1), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(G143), .B2(new_n214), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n390), .B1(new_n416), .B2(new_n314), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n417), .B1(new_n396), .B2(KEYINPUT1), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT68), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n400), .A2(new_n408), .A3(new_n419), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n420), .B(G131), .C1(new_n419), .C2(new_n400), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n413), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n385), .B1(new_n414), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n391), .A2(new_n396), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n397), .A2(new_n386), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n413), .ZN(new_n427));
  INV_X1    g241(.A(G131), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n409), .B1(new_n403), .B2(new_n404), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n428), .B1(new_n429), .B2(new_n406), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n426), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n413), .A2(new_n418), .A3(new_n421), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(KEYINPUT30), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n347), .A2(G116), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n286), .A2(G119), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(KEYINPUT2), .B(G113), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(KEYINPUT69), .B1(new_n434), .B2(new_n435), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(G116), .B(G119), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT69), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n438), .B1(new_n443), .B2(new_n437), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n423), .A2(new_n433), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n187), .A2(new_n188), .A3(G210), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(G101), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n448), .B(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n431), .A2(new_n444), .A3(new_n432), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n446), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT31), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT70), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g269(.A(KEYINPUT70), .B(KEYINPUT31), .Z(new_n456));
  NAND4_X1  g270(.A1(new_n446), .A2(new_n450), .A3(new_n451), .A4(new_n456), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n414), .A2(new_n422), .A3(new_n445), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(KEYINPUT28), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT28), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n444), .B1(new_n431), .B2(new_n432), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n460), .B1(new_n461), .B2(KEYINPUT71), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n445), .B1(new_n414), .B2(new_n422), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT71), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n451), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n459), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n455), .B(new_n457), .C1(new_n450), .C2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(G472), .A2(G902), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(KEYINPUT32), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT32), .B1(new_n467), .B2(new_n468), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT28), .B1(new_n458), .B2(new_n461), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n459), .B1(new_n473), .B2(KEYINPUT72), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT72), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n475), .B(KEYINPUT28), .C1(new_n458), .C2(new_n461), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n474), .A2(KEYINPUT29), .A3(new_n450), .A4(new_n476), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n466), .A2(new_n450), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n450), .B1(new_n446), .B2(new_n451), .ZN(new_n479));
  OR2_X1    g293(.A1(new_n479), .A2(KEYINPUT29), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n477), .B(new_n271), .C1(new_n478), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(G472), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n384), .B1(new_n472), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(G214), .B1(G237), .B2(G902), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  OAI22_X1  g299(.A1(new_n218), .A2(G107), .B1(KEYINPUT79), .B2(KEYINPUT3), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT80), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n218), .A3(G107), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT81), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n218), .A2(G107), .ZN(new_n491));
  AND2_X1   g305(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n492));
  NOR2_X1   g306(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT80), .B1(new_n295), .B2(G104), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n489), .A2(new_n490), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n486), .A2(new_n495), .A3(new_n488), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n295), .A2(G104), .ZN(new_n498));
  OR2_X1    g312(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n499));
  NAND2_X1  g313(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(KEYINPUT81), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n496), .A2(new_n502), .A3(G101), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT4), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(KEYINPUT82), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n496), .A2(new_n502), .A3(G101), .A4(new_n505), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n494), .A2(new_n495), .A3(new_n488), .A4(new_n486), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT83), .B(G101), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT4), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n507), .A2(new_n508), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n445), .ZN(new_n514));
  XOR2_X1   g328(.A(G110), .B(G122), .Z(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n438), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n434), .A2(new_n435), .A3(KEYINPUT69), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT5), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n518), .A2(new_n439), .A3(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(G113), .B1(new_n434), .B2(KEYINPUT5), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT84), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n295), .B2(G104), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n218), .A2(KEYINPUT84), .A3(G107), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n498), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G101), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n527), .B1(new_n509), .B2(new_n510), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT85), .B1(new_n522), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n440), .A2(new_n442), .A3(KEYINPUT5), .ZN(new_n530));
  INV_X1    g344(.A(new_n521), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n438), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n497), .A2(new_n501), .ZN(new_n533));
  INV_X1    g347(.A(new_n510), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n533), .A2(new_n534), .B1(G101), .B2(new_n526), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT85), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n532), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n529), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n514), .A2(new_n516), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT86), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n513), .A2(new_n445), .B1(new_n529), .B2(new_n537), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(KEYINPUT86), .A3(new_n516), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n515), .B(KEYINPUT8), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n522), .A2(new_n535), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n436), .A2(new_n519), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n517), .B1(new_n521), .B2(new_n547), .ZN(new_n548));
  AOI211_X1 g362(.A(new_n545), .B(new_n546), .C1(new_n535), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n418), .A2(new_n193), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n193), .B2(new_n398), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n188), .A2(G224), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(KEYINPUT7), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n551), .B1(KEYINPUT7), .B2(new_n552), .ZN(new_n555));
  NOR3_X1   g369(.A1(new_n549), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(G902), .B1(new_n544), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n542), .ZN(new_n558));
  AOI21_X1  g372(.A(KEYINPUT6), .B1(new_n558), .B2(new_n515), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n515), .ZN(new_n560));
  AND4_X1   g374(.A1(KEYINPUT86), .A2(new_n514), .A3(new_n516), .A4(new_n538), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT86), .B1(new_n542), .B2(new_n516), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n559), .B1(new_n563), .B2(KEYINPUT6), .ZN(new_n564));
  XOR2_X1   g378(.A(new_n551), .B(new_n552), .Z(new_n565));
  XOR2_X1   g379(.A(new_n565), .B(KEYINPUT87), .Z(new_n566));
  OAI21_X1  g380(.A(new_n557), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(G210), .B1(G237), .B2(G902), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n559), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n541), .A2(new_n543), .B1(new_n515), .B2(new_n558), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT6), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n566), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(new_n568), .A3(new_n557), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n485), .B1(new_n570), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(G221), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(new_n278), .B2(new_n222), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n412), .A2(new_n413), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n396), .A2(KEYINPUT1), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n584), .B1(new_n314), .B2(new_n416), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n528), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n535), .A2(new_n418), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n582), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT12), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI211_X1 g404(.A(KEYINPUT12), .B(new_n582), .C1(new_n586), .C2(new_n587), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n513), .A2(new_n426), .ZN(new_n593));
  INV_X1    g407(.A(new_n582), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n583), .A2(new_n585), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n535), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT10), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n418), .A2(KEYINPUT10), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n596), .A2(new_n597), .B1(new_n598), .B2(new_n535), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n593), .A2(new_n594), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n592), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n188), .A2(G227), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(KEYINPUT78), .ZN(new_n603));
  XNOR2_X1  g417(.A(G110), .B(G140), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n503), .A2(new_n506), .B1(KEYINPUT4), .B2(new_n511), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n398), .B1(new_n607), .B2(new_n508), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n598), .A2(new_n535), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n609), .B1(new_n586), .B2(KEYINPUT10), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n582), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n605), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(new_n600), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n606), .A2(G469), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(G469), .A2(G902), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n608), .A2(new_n610), .A3(new_n582), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n594), .B1(new_n593), .B2(new_n599), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n605), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n592), .A2(new_n600), .A3(new_n612), .ZN(new_n620));
  AOI211_X1 g434(.A(G469), .B(new_n270), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n581), .B1(new_n616), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n345), .A2(new_n483), .A3(new_n578), .A4(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(new_n510), .ZN(G3));
  NOR2_X1   g439(.A1(new_n567), .A2(new_n569), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n568), .B1(new_n576), .B2(new_n557), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n484), .B(new_n623), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(KEYINPUT99), .A2(KEYINPUT33), .ZN(new_n629));
  OR2_X1    g443(.A1(KEYINPUT99), .A2(KEYINPUT33), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n320), .A2(new_n321), .A3(new_n279), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n332), .B1(new_n331), .B2(new_n333), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n629), .B(new_n630), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n322), .A2(KEYINPUT99), .A3(new_n334), .A4(KEYINPUT33), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n270), .A2(new_n336), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n335), .A2(new_n336), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n639), .A2(new_n276), .A3(new_n266), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n467), .A2(new_n468), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT98), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n455), .A2(new_n457), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n462), .A2(new_n465), .ZN(new_n644));
  INV_X1    g458(.A(new_n459), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n450), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n642), .B(new_n271), .C1(new_n643), .C2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(G472), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n642), .B1(new_n467), .B2(new_n271), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n641), .B(new_n383), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n628), .A2(new_n640), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT34), .B(G104), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  OAI211_X1 g467(.A(new_n344), .B(new_n224), .C1(new_n247), .C2(new_n265), .ZN(new_n654));
  OR3_X1    g468(.A1(new_n654), .A2(KEYINPUT100), .A3(new_n277), .ZN(new_n655));
  AOI211_X1 g469(.A(new_n485), .B(new_n622), .C1(new_n570), .C2(new_n577), .ZN(new_n656));
  INV_X1    g470(.A(new_n650), .ZN(new_n657));
  OAI21_X1  g471(.A(KEYINPUT100), .B1(new_n654), .B2(new_n277), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n655), .A2(new_n656), .A3(new_n657), .A4(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n659), .B(KEYINPUT101), .Z(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT35), .B(G107), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  NOR2_X1   g476(.A1(new_n368), .A2(KEYINPUT36), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n364), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n373), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n380), .A2(new_n381), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n665), .B1(new_n666), .B2(new_n377), .ZN(new_n667));
  OAI211_X1 g481(.A(new_n667), .B(new_n641), .C1(new_n648), .C2(new_n649), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n345), .A2(new_n578), .A3(new_n623), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT37), .B(G110), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT102), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n670), .B(new_n672), .ZN(G12));
  INV_X1    g487(.A(G900), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n268), .B1(new_n272), .B2(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n654), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n667), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(new_n472), .B2(new_n482), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n656), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G128), .ZN(G30));
  NAND2_X1  g494(.A1(new_n570), .A2(new_n577), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT38), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n224), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n262), .A2(new_n263), .A3(new_n246), .ZN(new_n685));
  OAI21_X1  g499(.A(KEYINPUT20), .B1(new_n685), .B2(new_n226), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n264), .A2(new_n248), .A3(new_n225), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n684), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n344), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n691));
  INV_X1    g505(.A(new_n450), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n692), .B1(new_n458), .B2(new_n461), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n452), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n222), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n691), .B1(new_n452), .B2(new_n693), .ZN(new_n696));
  OAI21_X1  g510(.A(G472), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n667), .B1(new_n472), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n690), .A2(new_n698), .A3(new_n484), .ZN(new_n699));
  OAI21_X1  g513(.A(KEYINPUT104), .B1(new_n683), .B2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n681), .B(KEYINPUT38), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT104), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n690), .A2(new_n698), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n701), .A2(new_n702), .A3(new_n703), .A4(new_n484), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n675), .B(KEYINPUT39), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n623), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g521(.A(new_n707), .B(KEYINPUT40), .Z(new_n708));
  NAND3_X1  g522(.A1(new_n700), .A2(new_n704), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT105), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n700), .A2(new_n704), .A3(new_n711), .A4(new_n708), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n387), .ZN(G45));
  INV_X1    g528(.A(new_n675), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n639), .A2(new_n266), .A3(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n639), .A2(KEYINPUT106), .A3(new_n266), .A4(new_n715), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n718), .A2(new_n656), .A3(new_n678), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT107), .B(G146), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G48));
  AND3_X1   g536(.A1(new_n592), .A2(new_n600), .A3(new_n612), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n612), .B1(new_n611), .B2(new_n600), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n271), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(G469), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n619), .A2(new_n620), .ZN(new_n727));
  INV_X1    g541(.A(G469), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n728), .A3(new_n271), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n726), .A2(new_n581), .A3(new_n729), .ZN(new_n730));
  AOI211_X1 g544(.A(new_n485), .B(new_n730), .C1(new_n570), .C2(new_n577), .ZN(new_n731));
  AOI22_X1  g545(.A1(new_n635), .A2(new_n636), .B1(new_n336), .B2(new_n335), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n688), .A2(new_n732), .A3(new_n277), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n731), .A2(new_n483), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT41), .B(G113), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G15));
  NAND4_X1  g550(.A1(new_n655), .A2(new_n731), .A3(new_n483), .A4(new_n658), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G116), .ZN(G18));
  NOR3_X1   g552(.A1(new_n266), .A2(new_n677), .A3(new_n344), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n277), .B1(new_n472), .B2(new_n482), .ZN(new_n740));
  INV_X1    g554(.A(new_n730), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n739), .A2(new_n740), .A3(new_n578), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  NAND2_X1  g557(.A1(new_n467), .A2(new_n271), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(G472), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n450), .B1(new_n474), .B2(new_n476), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n468), .B1(new_n746), .B2(new_n643), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n748), .A2(new_n384), .A3(new_n277), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n690), .A2(new_n749), .A3(new_n578), .A4(new_n741), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G122), .ZN(G24));
  NOR2_X1   g565(.A1(new_n748), .A2(new_n677), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n718), .A2(new_n719), .A3(new_n731), .A4(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT108), .B(G125), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G27));
  NAND2_X1  g569(.A1(new_n718), .A2(new_n719), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n626), .A2(new_n627), .A3(new_n485), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(new_n470), .B2(new_n471), .ZN(new_n759));
  INV_X1    g573(.A(new_n471), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(KEYINPUT109), .A3(new_n469), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n759), .A2(new_n761), .A3(new_n482), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n757), .A2(new_n383), .A3(new_n762), .A4(new_n623), .ZN(new_n763));
  OAI21_X1  g577(.A(KEYINPUT42), .B1(new_n756), .B2(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n623), .A2(new_n570), .A3(new_n484), .A4(new_n577), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n482), .A2(new_n760), .A3(new_n469), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n383), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT42), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n768), .A2(new_n718), .A3(new_n769), .A4(new_n719), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n764), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(new_n428), .ZN(G33));
  NAND2_X1  g586(.A1(new_n768), .A2(new_n676), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G134), .ZN(G36));
  INV_X1    g588(.A(KEYINPUT110), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n688), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n266), .A2(KEYINPUT110), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n777), .A3(new_n639), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT43), .ZN(new_n779));
  OR3_X1    g593(.A1(new_n266), .A2(new_n732), .A3(KEYINPUT43), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n779), .A2(new_n780), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT111), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n648), .A2(new_n649), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n677), .B1(new_n786), .B2(new_n641), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n783), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT44), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n783), .A2(KEYINPUT44), .A3(new_n785), .A4(new_n787), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n617), .A2(new_n605), .ZN(new_n792));
  AOI22_X1  g606(.A1(new_n792), .A2(new_n611), .B1(new_n601), .B2(new_n605), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n793), .A2(KEYINPUT45), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(KEYINPUT45), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(G469), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(KEYINPUT46), .A3(new_n615), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n729), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT46), .B1(new_n796), .B2(new_n615), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(new_n581), .A3(new_n706), .ZN(new_n801));
  INV_X1    g615(.A(new_n757), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n790), .A2(new_n791), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G137), .ZN(G39));
  NOR4_X1   g619(.A1(new_n756), .A2(new_n766), .A3(new_n802), .A4(new_n383), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n800), .A2(new_n581), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT47), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n807), .A2(KEYINPUT47), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n806), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G140), .ZN(G42));
  NAND2_X1  g625(.A1(new_n726), .A2(new_n729), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(KEYINPUT49), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT112), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n472), .A2(new_n383), .A3(new_n697), .ZN(new_n815));
  AOI211_X1 g629(.A(new_n485), .B(new_n580), .C1(new_n812), .C2(KEYINPUT49), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  OR3_X1    g631(.A1(new_n817), .A2(new_n701), .A3(new_n778), .ZN(new_n818));
  NOR4_X1   g632(.A1(new_n681), .A2(new_n485), .A3(new_n269), .A4(new_n730), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n781), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n762), .A2(new_n383), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(KEYINPUT118), .B2(KEYINPUT48), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n824));
  OR2_X1    g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n748), .A2(new_n384), .A3(new_n269), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n781), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n731), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n819), .A2(new_n815), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n639), .A2(new_n266), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  AOI211_X1 g646(.A(new_n267), .B(G953), .C1(new_n830), .C2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n825), .A2(new_n826), .A3(new_n829), .A4(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n701), .A2(new_n484), .A3(new_n730), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n835), .A2(new_n781), .A3(new_n827), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT50), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n639), .A2(new_n266), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n830), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n820), .A2(new_n752), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n812), .A2(new_n581), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n845), .B1(new_n809), .B2(new_n808), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n828), .A2(new_n757), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT51), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n838), .A2(new_n844), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n842), .B(new_n843), .C1(new_n846), .C2(new_n847), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT51), .B1(new_n851), .B2(new_n837), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n834), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n737), .A2(new_n734), .A3(new_n742), .A4(new_n750), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n771), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n656), .A2(new_n715), .A3(new_n690), .A4(new_n698), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n720), .A2(new_n753), .A3(new_n679), .A4(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n857), .A2(new_n858), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n855), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n656), .A2(new_n733), .A3(new_n657), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT113), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n862), .A2(new_n863), .A3(new_n624), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n863), .B1(new_n862), .B2(new_n624), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n654), .A2(new_n277), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n867), .A2(new_n578), .A3(new_n657), .A4(new_n623), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n670), .A2(new_n868), .A3(KEYINPUT114), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT114), .B1(new_n670), .B2(new_n868), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n765), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n718), .A2(new_n872), .A3(new_n719), .A4(new_n752), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n872), .A2(new_n766), .A3(new_n715), .A4(new_n739), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n873), .A2(new_n874), .A3(new_n773), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n866), .A2(new_n871), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT53), .B1(new_n861), .B2(new_n877), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n734), .A2(new_n742), .A3(new_n750), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n879), .A2(new_n764), .A3(new_n737), .A4(new_n770), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n720), .A2(new_n679), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n881), .A2(KEYINPUT52), .A3(new_n753), .A4(new_n856), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n857), .A2(new_n858), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n880), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n688), .A2(new_n276), .A3(new_n689), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n628), .A2(new_n885), .A3(new_n767), .ZN(new_n886));
  OAI21_X1  g700(.A(KEYINPUT113), .B1(new_n651), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n670), .A2(new_n868), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT114), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n862), .A2(new_n863), .A3(new_n624), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n670), .A2(new_n868), .A3(KEYINPUT114), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n887), .A2(new_n890), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n875), .ZN(new_n894));
  XOR2_X1   g708(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n884), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n878), .A2(KEYINPUT54), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n896), .B1(new_n861), .B2(new_n877), .ZN(new_n899));
  OAI21_X1  g713(.A(KEYINPUT116), .B1(new_n893), .B2(new_n875), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT116), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n866), .A2(new_n901), .A3(new_n871), .A4(new_n876), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n884), .A2(new_n900), .A3(KEYINPUT53), .A4(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT54), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n899), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n853), .A2(new_n898), .A3(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(G952), .A2(G953), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT119), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n818), .B1(new_n906), .B2(new_n908), .ZN(G75));
  NAND2_X1  g723(.A1(new_n900), .A2(new_n902), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n855), .B(KEYINPUT53), .C1(new_n859), .C2(new_n860), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n895), .B1(new_n884), .B2(new_n894), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n270), .B(new_n569), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT56), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n271), .B1(new_n899), .B2(new_n903), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT120), .B1(new_n917), .B2(new_n569), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n564), .B(new_n575), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT55), .Z(new_n920));
  OAI21_X1  g734(.A(new_n916), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n920), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n914), .A2(KEYINPUT120), .A3(new_n915), .A4(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n188), .A2(G952), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n921), .A2(new_n923), .A3(new_n925), .ZN(G51));
  OAI21_X1  g740(.A(KEYINPUT54), .B1(new_n912), .B2(new_n913), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n905), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n615), .B(KEYINPUT57), .Z(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n727), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n917), .A2(G469), .A3(new_n795), .A4(new_n794), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n924), .B1(new_n931), .B2(new_n932), .ZN(G54));
  NAND3_X1  g747(.A1(new_n917), .A2(KEYINPUT58), .A3(G475), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n925), .B1(new_n934), .B2(new_n685), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n685), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(KEYINPUT121), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT121), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n934), .A2(new_n938), .A3(new_n685), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n935), .B1(new_n937), .B2(new_n939), .ZN(G60));
  XNOR2_X1  g754(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n941));
  NAND2_X1  g755(.A1(G478), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n941), .B(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n898), .B2(new_n905), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n925), .B1(new_n944), .B2(new_n635), .ZN(new_n945));
  INV_X1    g759(.A(new_n635), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n946), .A2(new_n943), .ZN(new_n947));
  AOI21_X1  g761(.A(KEYINPUT123), .B1(new_n928), .B2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT123), .ZN(new_n949));
  INV_X1    g763(.A(new_n947), .ZN(new_n950));
  AOI211_X1 g764(.A(new_n949), .B(new_n950), .C1(new_n927), .C2(new_n905), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n945), .A2(new_n948), .A3(new_n951), .ZN(G63));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n953));
  NAND2_X1  g767(.A1(G217), .A2(G902), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT60), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n955), .B1(new_n899), .B2(new_n903), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n664), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n925), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n369), .A2(new_n370), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n953), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n960), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n962), .A2(KEYINPUT61), .A3(new_n925), .A4(new_n957), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(new_n963), .ZN(G66));
  NOR2_X1   g778(.A1(new_n893), .A2(new_n854), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT124), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n966), .A2(G953), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n188), .B1(new_n274), .B2(G224), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n564), .B1(G898), .B2(new_n188), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT125), .Z(new_n971));
  XNOR2_X1  g785(.A(new_n969), .B(new_n971), .ZN(G69));
  INV_X1    g786(.A(G227), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n423), .A2(new_n433), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n228), .A2(new_n229), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  OAI221_X1 g791(.A(G953), .B1(new_n973), .B2(new_n674), .C1(new_n977), .C2(KEYINPUT126), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n757), .A2(new_n483), .A3(new_n623), .A4(new_n706), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n980), .B1(new_n831), .B2(new_n654), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT62), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n881), .A2(new_n753), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n982), .B1(new_n713), .B2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n983), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n985), .A2(new_n710), .A3(KEYINPUT62), .A4(new_n712), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n981), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n804), .A2(new_n810), .ZN(new_n988));
  AOI21_X1  g802(.A(G953), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n989), .A2(new_n976), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n674), .A2(new_n188), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n762), .A2(new_n690), .A3(new_n578), .A4(new_n383), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n773), .B1(new_n801), .B2(new_n992), .ZN(new_n993));
  NOR3_X1   g807(.A1(new_n983), .A2(new_n993), .A3(new_n771), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n804), .A2(new_n994), .A3(new_n810), .ZN(new_n995));
  AOI211_X1 g809(.A(new_n977), .B(new_n991), .C1(new_n995), .C2(new_n188), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n979), .B1(new_n990), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n995), .A2(new_n188), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n977), .A2(new_n991), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n1000), .B(new_n978), .C1(new_n989), .C2(new_n976), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n997), .A2(new_n1001), .ZN(G72));
  NAND2_X1  g816(.A1(new_n446), .A2(new_n451), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT127), .Z(new_n1004));
  NAND2_X1  g818(.A1(new_n995), .A2(new_n966), .ZN(new_n1005));
  NAND2_X1  g819(.A1(G472), .A2(G902), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n1006), .B(KEYINPUT63), .Z(new_n1007));
  AOI211_X1 g821(.A(new_n450), .B(new_n1004), .C1(new_n1005), .C2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1004), .A2(new_n450), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n987), .A2(new_n988), .A3(new_n966), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1009), .B1(new_n1010), .B2(new_n1007), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n878), .A2(new_n897), .ZN(new_n1012));
  INV_X1    g826(.A(new_n452), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1007), .B1(new_n1013), .B2(new_n479), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n925), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  NOR3_X1   g829(.A1(new_n1008), .A2(new_n1011), .A3(new_n1015), .ZN(G57));
endmodule


