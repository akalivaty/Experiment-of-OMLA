

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U553 ( .A1(n766), .A2(n765), .ZN(n520) );
  AND2_X1 U554 ( .A1(n797), .A2(n809), .ZN(n521) );
  INV_X1 U555 ( .A(KEYINPUT99), .ZN(n689) );
  NOR2_X1 U556 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U557 ( .A1(n695), .A2(n694), .ZN(n697) );
  BUF_X1 U558 ( .A(n698), .Z(n735) );
  AND2_X1 U559 ( .A1(n685), .A2(n684), .ZN(n730) );
  AND2_X1 U560 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U561 ( .A1(n682), .A2(n786), .ZN(n698) );
  XNOR2_X1 U562 ( .A(n683), .B(KEYINPUT93), .ZN(n684) );
  NOR2_X1 U563 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  NOR2_X1 U564 ( .A1(n803), .A2(n521), .ZN(n798) );
  NOR2_X1 U565 ( .A1(G651), .A2(n632), .ZN(n640) );
  NOR2_X1 U566 ( .A1(n532), .A2(n531), .ZN(G160) );
  INV_X1 U567 ( .A(G2104), .ZN(n527) );
  NOR2_X1 U568 ( .A1(G2105), .A2(n527), .ZN(n882) );
  NAND2_X1 U569 ( .A1(G101), .A2(n882), .ZN(n522) );
  XOR2_X1 U570 ( .A(KEYINPUT23), .B(n522), .Z(n526) );
  NAND2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  XOR2_X2 U572 ( .A(KEYINPUT64), .B(n523), .Z(n875) );
  NAND2_X1 U573 ( .A1(G113), .A2(n875), .ZN(n524) );
  XOR2_X1 U574 ( .A(KEYINPUT65), .B(n524), .Z(n525) );
  NAND2_X1 U575 ( .A1(n526), .A2(n525), .ZN(n532) );
  AND2_X1 U576 ( .A1(n527), .A2(G2105), .ZN(n874) );
  NAND2_X1 U577 ( .A1(G125), .A2(n874), .ZN(n530) );
  XOR2_X2 U578 ( .A(KEYINPUT17), .B(n528), .Z(n879) );
  NAND2_X1 U579 ( .A1(G137), .A2(n879), .ZN(n529) );
  NAND2_X1 U580 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U581 ( .A1(G138), .A2(n879), .ZN(n534) );
  NAND2_X1 U582 ( .A1(G102), .A2(n882), .ZN(n533) );
  NAND2_X1 U583 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U584 ( .A(n535), .B(KEYINPUT90), .ZN(n539) );
  NAND2_X1 U585 ( .A1(n874), .A2(G126), .ZN(n537) );
  NAND2_X1 U586 ( .A1(G114), .A2(n875), .ZN(n536) );
  NAND2_X1 U587 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U588 ( .A1(n539), .A2(n538), .ZN(G164) );
  NOR2_X1 U589 ( .A1(G651), .A2(G543), .ZN(n645) );
  NAND2_X1 U590 ( .A1(G85), .A2(n645), .ZN(n542) );
  INV_X1 U591 ( .A(G651), .ZN(n543) );
  NOR2_X1 U592 ( .A1(G543), .A2(n543), .ZN(n540) );
  XOR2_X1 U593 ( .A(KEYINPUT1), .B(n540), .Z(n639) );
  NAND2_X1 U594 ( .A1(G60), .A2(n639), .ZN(n541) );
  NAND2_X1 U595 ( .A1(n542), .A2(n541), .ZN(n547) );
  XOR2_X1 U596 ( .A(KEYINPUT0), .B(G543), .Z(n632) );
  NOR2_X1 U597 ( .A1(n632), .A2(n543), .ZN(n643) );
  NAND2_X1 U598 ( .A1(G72), .A2(n643), .ZN(n545) );
  NAND2_X1 U599 ( .A1(G47), .A2(n640), .ZN(n544) );
  NAND2_X1 U600 ( .A1(n545), .A2(n544), .ZN(n546) );
  OR2_X1 U601 ( .A1(n547), .A2(n546), .ZN(G290) );
  AND2_X1 U602 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U603 ( .A(G108), .ZN(G238) );
  INV_X1 U604 ( .A(G69), .ZN(G235) );
  NAND2_X1 U605 ( .A1(n643), .A2(G76), .ZN(n548) );
  XNOR2_X1 U606 ( .A(KEYINPUT74), .B(n548), .ZN(n551) );
  NAND2_X1 U607 ( .A1(n645), .A2(G89), .ZN(n549) );
  XNOR2_X1 U608 ( .A(KEYINPUT4), .B(n549), .ZN(n550) );
  NAND2_X1 U609 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U610 ( .A(n552), .B(KEYINPUT5), .ZN(n558) );
  NAND2_X1 U611 ( .A1(n639), .A2(G63), .ZN(n553) );
  XOR2_X1 U612 ( .A(KEYINPUT75), .B(n553), .Z(n555) );
  NAND2_X1 U613 ( .A1(n640), .A2(G51), .ZN(n554) );
  NAND2_X1 U614 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U615 ( .A(KEYINPUT6), .B(n556), .Z(n557) );
  NAND2_X1 U616 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U617 ( .A(n559), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U618 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U619 ( .A1(G7), .A2(G661), .ZN(n560) );
  XNOR2_X1 U620 ( .A(n560), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U621 ( .A(G567), .ZN(n677) );
  NOR2_X1 U622 ( .A1(n677), .A2(G223), .ZN(n561) );
  XNOR2_X1 U623 ( .A(n561), .B(KEYINPUT11), .ZN(G234) );
  NAND2_X1 U624 ( .A1(n645), .A2(G81), .ZN(n562) );
  XNOR2_X1 U625 ( .A(n562), .B(KEYINPUT12), .ZN(n564) );
  NAND2_X1 U626 ( .A1(G68), .A2(n643), .ZN(n563) );
  NAND2_X1 U627 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U628 ( .A(n565), .B(KEYINPUT13), .ZN(n567) );
  NAND2_X1 U629 ( .A1(G43), .A2(n640), .ZN(n566) );
  NAND2_X1 U630 ( .A1(n567), .A2(n566), .ZN(n570) );
  NAND2_X1 U631 ( .A1(n639), .A2(G56), .ZN(n568) );
  XOR2_X1 U632 ( .A(KEYINPUT14), .B(n568), .Z(n569) );
  NOR2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n1005) );
  NAND2_X1 U634 ( .A1(n1005), .A2(G860), .ZN(G153) );
  NAND2_X1 U635 ( .A1(n643), .A2(G77), .ZN(n571) );
  XNOR2_X1 U636 ( .A(KEYINPUT68), .B(n571), .ZN(n574) );
  NAND2_X1 U637 ( .A1(n645), .A2(G90), .ZN(n572) );
  XOR2_X1 U638 ( .A(KEYINPUT67), .B(n572), .Z(n573) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(KEYINPUT9), .ZN(n577) );
  NAND2_X1 U641 ( .A1(G52), .A2(n640), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n639), .A2(G64), .ZN(n578) );
  XOR2_X1 U644 ( .A(KEYINPUT66), .B(n578), .Z(n579) );
  NOR2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(KEYINPUT69), .B(n581), .ZN(G301) );
  NAND2_X1 U647 ( .A1(G868), .A2(G301), .ZN(n591) );
  NAND2_X1 U648 ( .A1(n640), .A2(G54), .ZN(n588) );
  NAND2_X1 U649 ( .A1(G92), .A2(n645), .ZN(n583) );
  NAND2_X1 U650 ( .A1(G79), .A2(n643), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U652 ( .A1(G66), .A2(n639), .ZN(n584) );
  XNOR2_X1 U653 ( .A(KEYINPUT73), .B(n584), .ZN(n585) );
  NOR2_X1 U654 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U655 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U656 ( .A(KEYINPUT15), .B(n589), .Z(n1004) );
  INV_X1 U657 ( .A(G868), .ZN(n652) );
  NAND2_X1 U658 ( .A1(n1004), .A2(n652), .ZN(n590) );
  NAND2_X1 U659 ( .A1(n591), .A2(n590), .ZN(G284) );
  NAND2_X1 U660 ( .A1(G91), .A2(n645), .ZN(n593) );
  NAND2_X1 U661 ( .A1(G78), .A2(n643), .ZN(n592) );
  NAND2_X1 U662 ( .A1(n593), .A2(n592), .ZN(n596) );
  NAND2_X1 U663 ( .A1(n640), .A2(G53), .ZN(n594) );
  XOR2_X1 U664 ( .A(KEYINPUT70), .B(n594), .Z(n595) );
  NOR2_X1 U665 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U666 ( .A1(n639), .A2(G65), .ZN(n597) );
  NAND2_X1 U667 ( .A1(n598), .A2(n597), .ZN(n994) );
  XOR2_X1 U668 ( .A(KEYINPUT71), .B(n994), .Z(G299) );
  NAND2_X1 U669 ( .A1(G286), .A2(G868), .ZN(n600) );
  NAND2_X1 U670 ( .A1(G299), .A2(n652), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(G297) );
  INV_X1 U672 ( .A(G860), .ZN(n601) );
  NAND2_X1 U673 ( .A1(n601), .A2(G559), .ZN(n602) );
  INV_X1 U674 ( .A(n1004), .ZN(n890) );
  NAND2_X1 U675 ( .A1(n602), .A2(n890), .ZN(n603) );
  XNOR2_X1 U676 ( .A(n603), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U677 ( .A1(n890), .A2(G868), .ZN(n604) );
  NOR2_X1 U678 ( .A1(G559), .A2(n604), .ZN(n606) );
  AND2_X1 U679 ( .A1(n652), .A2(n1005), .ZN(n605) );
  NOR2_X1 U680 ( .A1(n606), .A2(n605), .ZN(G282) );
  NAND2_X1 U681 ( .A1(G123), .A2(n874), .ZN(n607) );
  XNOR2_X1 U682 ( .A(n607), .B(KEYINPUT18), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n882), .A2(G99), .ZN(n608) );
  NAND2_X1 U684 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U685 ( .A1(n879), .A2(G135), .ZN(n611) );
  NAND2_X1 U686 ( .A1(G111), .A2(n875), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U688 ( .A1(n613), .A2(n612), .ZN(n925) );
  XNOR2_X1 U689 ( .A(n925), .B(G2096), .ZN(n615) );
  INV_X1 U690 ( .A(G2100), .ZN(n614) );
  NAND2_X1 U691 ( .A1(n615), .A2(n614), .ZN(G156) );
  NAND2_X1 U692 ( .A1(G88), .A2(n645), .ZN(n617) );
  NAND2_X1 U693 ( .A1(G75), .A2(n643), .ZN(n616) );
  NAND2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U695 ( .A(KEYINPUT83), .B(n618), .ZN(n622) );
  NAND2_X1 U696 ( .A1(G62), .A2(n639), .ZN(n620) );
  NAND2_X1 U697 ( .A1(G50), .A2(n640), .ZN(n619) );
  AND2_X1 U698 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n622), .A2(n621), .ZN(G303) );
  INV_X1 U700 ( .A(G303), .ZN(G166) );
  NAND2_X1 U701 ( .A1(n643), .A2(G73), .ZN(n624) );
  XNOR2_X1 U702 ( .A(KEYINPUT2), .B(KEYINPUT82), .ZN(n623) );
  XNOR2_X1 U703 ( .A(n624), .B(n623), .ZN(n631) );
  NAND2_X1 U704 ( .A1(G86), .A2(n645), .ZN(n626) );
  NAND2_X1 U705 ( .A1(G48), .A2(n640), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U707 ( .A1(G61), .A2(n639), .ZN(n627) );
  XNOR2_X1 U708 ( .A(KEYINPUT81), .B(n627), .ZN(n628) );
  NOR2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n631), .A2(n630), .ZN(G305) );
  NAND2_X1 U711 ( .A1(G74), .A2(G651), .ZN(n637) );
  NAND2_X1 U712 ( .A1(G49), .A2(n640), .ZN(n634) );
  NAND2_X1 U713 ( .A1(G87), .A2(n632), .ZN(n633) );
  NAND2_X1 U714 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U715 ( .A1(n639), .A2(n635), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U717 ( .A(n638), .B(KEYINPUT80), .ZN(G288) );
  NAND2_X1 U718 ( .A1(G67), .A2(n639), .ZN(n642) );
  NAND2_X1 U719 ( .A1(G55), .A2(n640), .ZN(n641) );
  NAND2_X1 U720 ( .A1(n642), .A2(n641), .ZN(n650) );
  NAND2_X1 U721 ( .A1(n643), .A2(G80), .ZN(n644) );
  XNOR2_X1 U722 ( .A(n644), .B(KEYINPUT76), .ZN(n647) );
  NAND2_X1 U723 ( .A1(G93), .A2(n645), .ZN(n646) );
  NAND2_X1 U724 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U725 ( .A(KEYINPUT77), .B(n648), .Z(n649) );
  NOR2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U727 ( .A(KEYINPUT78), .B(n651), .Z(n822) );
  NAND2_X1 U728 ( .A1(n652), .A2(n822), .ZN(n653) );
  XNOR2_X1 U729 ( .A(n653), .B(KEYINPUT86), .ZN(n664) );
  XNOR2_X1 U730 ( .A(KEYINPUT19), .B(KEYINPUT84), .ZN(n655) );
  XNOR2_X1 U731 ( .A(G290), .B(KEYINPUT85), .ZN(n654) );
  XNOR2_X1 U732 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U733 ( .A(G299), .B(n656), .ZN(n658) );
  XNOR2_X1 U734 ( .A(n1005), .B(G166), .ZN(n657) );
  XNOR2_X1 U735 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U736 ( .A(n822), .B(n659), .ZN(n661) );
  XNOR2_X1 U737 ( .A(G305), .B(G288), .ZN(n660) );
  XNOR2_X1 U738 ( .A(n661), .B(n660), .ZN(n889) );
  NAND2_X1 U739 ( .A1(n890), .A2(G559), .ZN(n818) );
  XNOR2_X1 U740 ( .A(n889), .B(n818), .ZN(n662) );
  NAND2_X1 U741 ( .A1(G868), .A2(n662), .ZN(n663) );
  NAND2_X1 U742 ( .A1(n664), .A2(n663), .ZN(G295) );
  NAND2_X1 U743 ( .A1(G2084), .A2(G2078), .ZN(n665) );
  XOR2_X1 U744 ( .A(KEYINPUT20), .B(n665), .Z(n666) );
  NAND2_X1 U745 ( .A1(G2090), .A2(n666), .ZN(n668) );
  XOR2_X1 U746 ( .A(KEYINPUT21), .B(KEYINPUT87), .Z(n667) );
  XNOR2_X1 U747 ( .A(n668), .B(n667), .ZN(n669) );
  NAND2_X1 U748 ( .A1(G2072), .A2(n669), .ZN(G158) );
  XNOR2_X1 U749 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U750 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  NAND2_X1 U751 ( .A1(G132), .A2(G82), .ZN(n670) );
  XNOR2_X1 U752 ( .A(n670), .B(KEYINPUT22), .ZN(n671) );
  XNOR2_X1 U753 ( .A(n671), .B(KEYINPUT88), .ZN(n672) );
  NOR2_X1 U754 ( .A1(G218), .A2(n672), .ZN(n673) );
  NAND2_X1 U755 ( .A1(G96), .A2(n673), .ZN(n823) );
  NAND2_X1 U756 ( .A1(G2106), .A2(n823), .ZN(n674) );
  XNOR2_X1 U757 ( .A(n674), .B(KEYINPUT89), .ZN(n679) );
  NOR2_X1 U758 ( .A1(G237), .A2(G238), .ZN(n675) );
  NAND2_X1 U759 ( .A1(G120), .A2(n675), .ZN(n676) );
  NOR2_X1 U760 ( .A1(G235), .A2(n676), .ZN(n825) );
  NOR2_X1 U761 ( .A1(n677), .A2(n825), .ZN(n678) );
  NOR2_X1 U762 ( .A1(n679), .A2(n678), .ZN(G319) );
  INV_X1 U763 ( .A(G319), .ZN(n681) );
  NAND2_X1 U764 ( .A1(G483), .A2(G661), .ZN(n680) );
  NOR2_X1 U765 ( .A1(n681), .A2(n680), .ZN(n817) );
  NAND2_X1 U766 ( .A1(n817), .A2(G36), .ZN(G176) );
  INV_X1 U767 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U768 ( .A(G1981), .B(G305), .ZN(n1013) );
  AND2_X1 U769 ( .A1(G160), .A2(G40), .ZN(n682) );
  NOR2_X1 U770 ( .A1(G164), .A2(G1384), .ZN(n786) );
  NAND2_X1 U771 ( .A1(n698), .A2(G8), .ZN(n683) );
  INV_X1 U772 ( .A(n684), .ZN(n750) );
  NOR2_X1 U773 ( .A1(G2084), .A2(n735), .ZN(n688) );
  NAND2_X1 U774 ( .A1(G8), .A2(n688), .ZN(n732) );
  INV_X1 U775 ( .A(G1966), .ZN(n685) );
  XNOR2_X1 U776 ( .A(G2078), .B(KEYINPUT25), .ZN(n969) );
  NOR2_X1 U777 ( .A1(n735), .A2(n969), .ZN(n687) );
  AND2_X1 U778 ( .A1(n735), .A2(G1961), .ZN(n686) );
  NOR2_X1 U779 ( .A1(n687), .A2(n686), .ZN(n724) );
  NOR2_X1 U780 ( .A1(G171), .A2(n724), .ZN(n695) );
  NOR2_X1 U781 ( .A1(n730), .A2(n688), .ZN(n690) );
  XNOR2_X1 U782 ( .A(n690), .B(n689), .ZN(n691) );
  NAND2_X1 U783 ( .A1(n691), .A2(G8), .ZN(n692) );
  XNOR2_X1 U784 ( .A(KEYINPUT30), .B(n692), .ZN(n693) );
  NOR2_X1 U785 ( .A1(G168), .A2(n693), .ZN(n694) );
  XOR2_X1 U786 ( .A(KEYINPUT100), .B(KEYINPUT31), .Z(n696) );
  XNOR2_X1 U787 ( .A(n697), .B(n696), .ZN(n728) );
  INV_X1 U788 ( .A(n698), .ZN(n707) );
  NAND2_X1 U789 ( .A1(n707), .A2(G2072), .ZN(n699) );
  XOR2_X1 U790 ( .A(KEYINPUT27), .B(n699), .Z(n701) );
  NAND2_X1 U791 ( .A1(G1956), .A2(n735), .ZN(n700) );
  NAND2_X1 U792 ( .A1(n701), .A2(n700), .ZN(n719) );
  NOR2_X1 U793 ( .A1(n994), .A2(n719), .ZN(n702) );
  XNOR2_X1 U794 ( .A(KEYINPUT98), .B(n702), .ZN(n718) );
  XOR2_X1 U795 ( .A(G1996), .B(KEYINPUT95), .Z(n964) );
  NAND2_X1 U796 ( .A1(n707), .A2(n964), .ZN(n703) );
  XNOR2_X1 U797 ( .A(n703), .B(KEYINPUT26), .ZN(n705) );
  NAND2_X1 U798 ( .A1(G1341), .A2(n735), .ZN(n704) );
  NAND2_X1 U799 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U800 ( .A(KEYINPUT96), .B(n706), .ZN(n712) );
  NAND2_X1 U801 ( .A1(G1348), .A2(n735), .ZN(n709) );
  NAND2_X1 U802 ( .A1(n707), .A2(G2067), .ZN(n708) );
  NAND2_X1 U803 ( .A1(n709), .A2(n708), .ZN(n713) );
  NAND2_X1 U804 ( .A1(n1004), .A2(n713), .ZN(n710) );
  NAND2_X1 U805 ( .A1(n1005), .A2(n710), .ZN(n711) );
  NOR2_X1 U806 ( .A1(n712), .A2(n711), .ZN(n715) );
  NOR2_X1 U807 ( .A1(n713), .A2(n1004), .ZN(n714) );
  NOR2_X1 U808 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U809 ( .A(KEYINPUT97), .B(n716), .ZN(n717) );
  NOR2_X1 U810 ( .A1(n718), .A2(n717), .ZN(n722) );
  NAND2_X1 U811 ( .A1(n994), .A2(n719), .ZN(n720) );
  XOR2_X1 U812 ( .A(KEYINPUT28), .B(n720), .Z(n721) );
  XNOR2_X1 U813 ( .A(n723), .B(KEYINPUT29), .ZN(n726) );
  NAND2_X1 U814 ( .A1(n724), .A2(G171), .ZN(n725) );
  NAND2_X1 U815 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U816 ( .A1(n728), .A2(n727), .ZN(n734) );
  INV_X1 U817 ( .A(n734), .ZN(n729) );
  NOR2_X1 U818 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U819 ( .A1(n732), .A2(n731), .ZN(n745) );
  AND2_X1 U820 ( .A1(G286), .A2(G8), .ZN(n733) );
  NAND2_X1 U821 ( .A1(n734), .A2(n733), .ZN(n742) );
  INV_X1 U822 ( .A(G8), .ZN(n740) );
  NOR2_X1 U823 ( .A1(G1971), .A2(n750), .ZN(n737) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n735), .ZN(n736) );
  NOR2_X1 U825 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U826 ( .A1(n738), .A2(G303), .ZN(n739) );
  OR2_X1 U827 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U828 ( .A(n743), .B(KEYINPUT32), .ZN(n744) );
  NAND2_X1 U829 ( .A1(n745), .A2(n744), .ZN(n760) );
  NOR2_X1 U830 ( .A1(G1976), .A2(G288), .ZN(n753) );
  NOR2_X1 U831 ( .A1(G1971), .A2(G303), .ZN(n746) );
  NOR2_X1 U832 ( .A1(n753), .A2(n746), .ZN(n998) );
  XOR2_X1 U833 ( .A(n998), .B(KEYINPUT101), .Z(n747) );
  NAND2_X1 U834 ( .A1(n760), .A2(n747), .ZN(n748) );
  NAND2_X1 U835 ( .A1(G1976), .A2(G288), .ZN(n997) );
  NAND2_X1 U836 ( .A1(n748), .A2(n997), .ZN(n749) );
  NOR2_X1 U837 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U838 ( .A1(n751), .A2(KEYINPUT33), .ZN(n752) );
  NOR2_X1 U839 ( .A1(n1013), .A2(n752), .ZN(n756) );
  AND2_X1 U840 ( .A1(n753), .A2(KEYINPUT33), .ZN(n754) );
  NAND2_X1 U841 ( .A1(n754), .A2(n684), .ZN(n755) );
  AND2_X1 U842 ( .A1(n756), .A2(n755), .ZN(n767) );
  NOR2_X1 U843 ( .A1(G1981), .A2(G305), .ZN(n757) );
  XNOR2_X1 U844 ( .A(n757), .B(KEYINPUT94), .ZN(n758) );
  XNOR2_X1 U845 ( .A(n758), .B(KEYINPUT24), .ZN(n759) );
  AND2_X1 U846 ( .A1(n759), .A2(n684), .ZN(n766) );
  INV_X1 U847 ( .A(n760), .ZN(n763) );
  NAND2_X1 U848 ( .A1(G166), .A2(G8), .ZN(n761) );
  NOR2_X1 U849 ( .A1(G2090), .A2(n761), .ZN(n762) );
  NOR2_X1 U850 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U851 ( .A1(n684), .A2(n764), .ZN(n765) );
  NOR2_X1 U852 ( .A1(n767), .A2(n520), .ZN(n768) );
  INV_X1 U853 ( .A(n768), .ZN(n799) );
  XNOR2_X1 U854 ( .A(KEYINPUT92), .B(G1991), .ZN(n966) );
  NAND2_X1 U855 ( .A1(G95), .A2(n882), .ZN(n770) );
  NAND2_X1 U856 ( .A1(G131), .A2(n879), .ZN(n769) );
  NAND2_X1 U857 ( .A1(n770), .A2(n769), .ZN(n773) );
  NAND2_X1 U858 ( .A1(G119), .A2(n874), .ZN(n771) );
  XNOR2_X1 U859 ( .A(KEYINPUT91), .B(n771), .ZN(n772) );
  NOR2_X1 U860 ( .A1(n773), .A2(n772), .ZN(n775) );
  NAND2_X1 U861 ( .A1(G107), .A2(n875), .ZN(n774) );
  NAND2_X1 U862 ( .A1(n775), .A2(n774), .ZN(n866) );
  AND2_X1 U863 ( .A1(n966), .A2(n866), .ZN(n784) );
  NAND2_X1 U864 ( .A1(G129), .A2(n874), .ZN(n777) );
  NAND2_X1 U865 ( .A1(G141), .A2(n879), .ZN(n776) );
  NAND2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n780) );
  NAND2_X1 U867 ( .A1(n882), .A2(G105), .ZN(n778) );
  XOR2_X1 U868 ( .A(KEYINPUT38), .B(n778), .Z(n779) );
  NOR2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n782) );
  NAND2_X1 U870 ( .A1(G117), .A2(n875), .ZN(n781) );
  NAND2_X1 U871 ( .A1(n782), .A2(n781), .ZN(n861) );
  AND2_X1 U872 ( .A1(n861), .A2(G1996), .ZN(n783) );
  NOR2_X1 U873 ( .A1(n784), .A2(n783), .ZN(n930) );
  NAND2_X1 U874 ( .A1(G160), .A2(G40), .ZN(n785) );
  NOR2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n809) );
  INV_X1 U876 ( .A(n809), .ZN(n787) );
  NOR2_X1 U877 ( .A1(n930), .A2(n787), .ZN(n803) );
  XOR2_X1 U878 ( .A(G1986), .B(G290), .Z(n996) );
  XNOR2_X1 U879 ( .A(G2067), .B(KEYINPUT37), .ZN(n800) );
  NAND2_X1 U880 ( .A1(n874), .A2(G128), .ZN(n789) );
  NAND2_X1 U881 ( .A1(G116), .A2(n875), .ZN(n788) );
  NAND2_X1 U882 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U883 ( .A(n790), .B(KEYINPUT35), .ZN(n795) );
  NAND2_X1 U884 ( .A1(G104), .A2(n882), .ZN(n792) );
  NAND2_X1 U885 ( .A1(G140), .A2(n879), .ZN(n791) );
  NAND2_X1 U886 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U887 ( .A(KEYINPUT34), .B(n793), .Z(n794) );
  NAND2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U889 ( .A(n796), .B(KEYINPUT36), .Z(n871) );
  OR2_X1 U890 ( .A1(n800), .A2(n871), .ZN(n929) );
  NAND2_X1 U891 ( .A1(n996), .A2(n929), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n799), .A2(n798), .ZN(n812) );
  NAND2_X1 U893 ( .A1(n800), .A2(n871), .ZN(n918) );
  NOR2_X1 U894 ( .A1(G1996), .A2(n861), .ZN(n921) );
  NOR2_X1 U895 ( .A1(G1986), .A2(G290), .ZN(n801) );
  NOR2_X1 U896 ( .A1(n966), .A2(n866), .ZN(n926) );
  NOR2_X1 U897 ( .A1(n801), .A2(n926), .ZN(n802) );
  NOR2_X1 U898 ( .A1(n803), .A2(n802), .ZN(n804) );
  NOR2_X1 U899 ( .A1(n921), .A2(n804), .ZN(n805) );
  XNOR2_X1 U900 ( .A(KEYINPUT39), .B(n805), .ZN(n806) );
  XNOR2_X1 U901 ( .A(n806), .B(KEYINPUT102), .ZN(n807) );
  NAND2_X1 U902 ( .A1(n807), .A2(n929), .ZN(n808) );
  NAND2_X1 U903 ( .A1(n918), .A2(n808), .ZN(n810) );
  NAND2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U905 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U906 ( .A(n813), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U907 ( .A(G223), .ZN(n814) );
  NAND2_X1 U908 ( .A1(G2106), .A2(n814), .ZN(G217) );
  AND2_X1 U909 ( .A1(G15), .A2(G2), .ZN(n815) );
  NAND2_X1 U910 ( .A1(G661), .A2(n815), .ZN(G259) );
  NAND2_X1 U911 ( .A1(G3), .A2(G1), .ZN(n816) );
  NAND2_X1 U912 ( .A1(n817), .A2(n816), .ZN(G188) );
  XOR2_X1 U914 ( .A(n818), .B(n1005), .Z(n819) );
  NOR2_X1 U915 ( .A1(G860), .A2(n819), .ZN(n820) );
  XOR2_X1 U916 ( .A(KEYINPUT79), .B(n820), .Z(n821) );
  XOR2_X1 U917 ( .A(n822), .B(n821), .Z(G145) );
  INV_X1 U918 ( .A(G132), .ZN(G219) );
  INV_X1 U919 ( .A(G82), .ZN(G220) );
  INV_X1 U920 ( .A(n823), .ZN(n824) );
  NAND2_X1 U921 ( .A1(n825), .A2(n824), .ZN(G261) );
  INV_X1 U922 ( .A(G261), .ZN(G325) );
  XOR2_X1 U923 ( .A(G2100), .B(G2096), .Z(n827) );
  XNOR2_X1 U924 ( .A(KEYINPUT42), .B(G2678), .ZN(n826) );
  XNOR2_X1 U925 ( .A(n827), .B(n826), .ZN(n831) );
  XOR2_X1 U926 ( .A(KEYINPUT43), .B(G2090), .Z(n829) );
  XNOR2_X1 U927 ( .A(G2072), .B(G2067), .ZN(n828) );
  XNOR2_X1 U928 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U929 ( .A(n831), .B(n830), .Z(n833) );
  XNOR2_X1 U930 ( .A(G2084), .B(G2078), .ZN(n832) );
  XNOR2_X1 U931 ( .A(n833), .B(n832), .ZN(G227) );
  XOR2_X1 U932 ( .A(KEYINPUT107), .B(KEYINPUT41), .Z(n835) );
  XNOR2_X1 U933 ( .A(G2474), .B(KEYINPUT108), .ZN(n834) );
  XNOR2_X1 U934 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U935 ( .A(n836), .B(KEYINPUT105), .Z(n838) );
  XNOR2_X1 U936 ( .A(G1971), .B(G1986), .ZN(n837) );
  XNOR2_X1 U937 ( .A(n838), .B(n837), .ZN(n846) );
  XOR2_X1 U938 ( .A(G1976), .B(G1981), .Z(n840) );
  XNOR2_X1 U939 ( .A(G1966), .B(G1961), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U941 ( .A(KEYINPUT106), .B(G1991), .Z(n842) );
  XNOR2_X1 U942 ( .A(G1956), .B(G1996), .ZN(n841) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U944 ( .A(n844), .B(n843), .Z(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(G229) );
  NAND2_X1 U946 ( .A1(G124), .A2(n874), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n847), .B(KEYINPUT44), .ZN(n849) );
  NAND2_X1 U948 ( .A1(n882), .A2(G100), .ZN(n848) );
  NAND2_X1 U949 ( .A1(n849), .A2(n848), .ZN(n853) );
  NAND2_X1 U950 ( .A1(n879), .A2(G136), .ZN(n851) );
  NAND2_X1 U951 ( .A1(G112), .A2(n875), .ZN(n850) );
  NAND2_X1 U952 ( .A1(n851), .A2(n850), .ZN(n852) );
  NOR2_X1 U953 ( .A1(n853), .A2(n852), .ZN(G162) );
  NAND2_X1 U954 ( .A1(n874), .A2(G130), .ZN(n855) );
  NAND2_X1 U955 ( .A1(G118), .A2(n875), .ZN(n854) );
  NAND2_X1 U956 ( .A1(n855), .A2(n854), .ZN(n860) );
  NAND2_X1 U957 ( .A1(G106), .A2(n882), .ZN(n857) );
  NAND2_X1 U958 ( .A1(G142), .A2(n879), .ZN(n856) );
  NAND2_X1 U959 ( .A1(n857), .A2(n856), .ZN(n858) );
  XOR2_X1 U960 ( .A(n858), .B(KEYINPUT45), .Z(n859) );
  NOR2_X1 U961 ( .A1(n860), .A2(n859), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n862), .B(n861), .ZN(n870) );
  XOR2_X1 U963 ( .A(KEYINPUT46), .B(KEYINPUT109), .Z(n864) );
  XNOR2_X1 U964 ( .A(KEYINPUT111), .B(KEYINPUT48), .ZN(n863) );
  XNOR2_X1 U965 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U966 ( .A(n865), .B(n925), .Z(n868) );
  XOR2_X1 U967 ( .A(n866), .B(G162), .Z(n867) );
  XNOR2_X1 U968 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U969 ( .A(n870), .B(n869), .Z(n873) );
  XOR2_X1 U970 ( .A(G160), .B(n871), .Z(n872) );
  XNOR2_X1 U971 ( .A(n873), .B(n872), .ZN(n887) );
  NAND2_X1 U972 ( .A1(n874), .A2(G127), .ZN(n877) );
  NAND2_X1 U973 ( .A1(G115), .A2(n875), .ZN(n876) );
  NAND2_X1 U974 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U975 ( .A(n878), .B(KEYINPUT47), .ZN(n881) );
  NAND2_X1 U976 ( .A1(G139), .A2(n879), .ZN(n880) );
  NAND2_X1 U977 ( .A1(n881), .A2(n880), .ZN(n885) );
  NAND2_X1 U978 ( .A1(n882), .A2(G103), .ZN(n883) );
  XOR2_X1 U979 ( .A(KEYINPUT110), .B(n883), .Z(n884) );
  NOR2_X1 U980 ( .A1(n885), .A2(n884), .ZN(n912) );
  XOR2_X1 U981 ( .A(n912), .B(G164), .Z(n886) );
  XNOR2_X1 U982 ( .A(n887), .B(n886), .ZN(n888) );
  NOR2_X1 U983 ( .A1(G37), .A2(n888), .ZN(G395) );
  XOR2_X1 U984 ( .A(KEYINPUT112), .B(n889), .Z(n892) );
  XNOR2_X1 U985 ( .A(n890), .B(G286), .ZN(n891) );
  XNOR2_X1 U986 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U987 ( .A(G171), .B(n893), .ZN(n894) );
  NOR2_X1 U988 ( .A1(G37), .A2(n894), .ZN(G397) );
  XNOR2_X1 U989 ( .A(G2435), .B(G2427), .ZN(n904) );
  XOR2_X1 U990 ( .A(G2454), .B(G2430), .Z(n896) );
  XNOR2_X1 U991 ( .A(G2443), .B(G2451), .ZN(n895) );
  XNOR2_X1 U992 ( .A(n896), .B(n895), .ZN(n900) );
  XOR2_X1 U993 ( .A(G2446), .B(KEYINPUT103), .Z(n898) );
  XNOR2_X1 U994 ( .A(G1348), .B(G1341), .ZN(n897) );
  XNOR2_X1 U995 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U996 ( .A(n900), .B(n899), .Z(n902) );
  XNOR2_X1 U997 ( .A(KEYINPUT104), .B(G2438), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n905) );
  NAND2_X1 U1000 ( .A1(n905), .A2(G14), .ZN(n911) );
  NAND2_X1 U1001 ( .A1(G319), .A2(n911), .ZN(n908) );
  NOR2_X1 U1002 ( .A1(G227), .A2(G229), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(KEYINPUT49), .B(n906), .ZN(n907) );
  NOR2_X1 U1004 ( .A1(n908), .A2(n907), .ZN(n910) );
  NOR2_X1 U1005 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1006 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1007 ( .A(G225), .ZN(G308) );
  INV_X1 U1008 ( .A(G120), .ZN(G236) );
  INV_X1 U1009 ( .A(G96), .ZN(G221) );
  INV_X1 U1010 ( .A(n911), .ZN(G401) );
  XNOR2_X1 U1011 ( .A(KEYINPUT55), .B(KEYINPUT116), .ZN(n985) );
  XNOR2_X1 U1012 ( .A(G2072), .B(n912), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(n913), .B(KEYINPUT113), .ZN(n916) );
  XOR2_X1 U1014 ( .A(G2078), .B(G164), .Z(n914) );
  XNOR2_X1 U1015 ( .A(KEYINPUT114), .B(n914), .ZN(n915) );
  NOR2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(n917), .B(KEYINPUT50), .ZN(n919) );
  NAND2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n924) );
  XOR2_X1 U1019 ( .A(G2090), .B(G162), .Z(n920) );
  NOR2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(n922), .B(KEYINPUT51), .ZN(n923) );
  NOR2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n934) );
  XNOR2_X1 U1023 ( .A(G160), .B(G2084), .ZN(n928) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n932) );
  NAND2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1028 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1029 ( .A(KEYINPUT115), .B(n935), .ZN(n936) );
  XOR2_X1 U1030 ( .A(KEYINPUT52), .B(n936), .Z(n937) );
  NOR2_X1 U1031 ( .A1(n985), .A2(n937), .ZN(n938) );
  XNOR2_X1 U1032 ( .A(KEYINPUT117), .B(n938), .ZN(n939) );
  NAND2_X1 U1033 ( .A1(n939), .A2(G29), .ZN(n993) );
  XOR2_X1 U1034 ( .A(G1986), .B(G24), .Z(n943) );
  XNOR2_X1 U1035 ( .A(G1971), .B(G22), .ZN(n941) );
  XNOR2_X1 U1036 ( .A(G23), .B(G1976), .ZN(n940) );
  NOR2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n945) );
  XNOR2_X1 U1039 ( .A(KEYINPUT58), .B(KEYINPUT127), .ZN(n944) );
  XNOR2_X1 U1040 ( .A(n945), .B(n944), .ZN(n949) );
  XNOR2_X1 U1041 ( .A(G1966), .B(G21), .ZN(n947) );
  XNOR2_X1 U1042 ( .A(G1961), .B(G5), .ZN(n946) );
  NOR2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n961) );
  XNOR2_X1 U1045 ( .A(G1956), .B(G20), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(G6), .B(G1981), .ZN(n950) );
  NOR2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n958) );
  XOR2_X1 U1048 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n953) );
  XNOR2_X1 U1049 ( .A(KEYINPUT59), .B(G4), .ZN(n952) );
  XNOR2_X1 U1050 ( .A(n953), .B(n952), .ZN(n954) );
  XOR2_X1 U1051 ( .A(G1348), .B(n954), .Z(n956) );
  XNOR2_X1 U1052 ( .A(G19), .B(G1341), .ZN(n955) );
  NOR2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(KEYINPUT60), .B(n959), .ZN(n960) );
  NOR2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1057 ( .A(KEYINPUT61), .B(n962), .Z(n963) );
  NOR2_X1 U1058 ( .A1(G16), .A2(n963), .ZN(n991) );
  XOR2_X1 U1059 ( .A(G29), .B(KEYINPUT120), .Z(n987) );
  XOR2_X1 U1060 ( .A(n964), .B(G32), .Z(n965) );
  NAND2_X1 U1061 ( .A1(G28), .A2(n965), .ZN(n968) );
  XNOR2_X1 U1062 ( .A(G25), .B(n966), .ZN(n967) );
  NOR2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n977) );
  XOR2_X1 U1064 ( .A(n969), .B(G27), .Z(n975) );
  XNOR2_X1 U1065 ( .A(G2067), .B(G26), .ZN(n970) );
  XNOR2_X1 U1066 ( .A(n970), .B(KEYINPUT118), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(G33), .B(G2072), .ZN(n971) );
  NOR2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1069 ( .A(KEYINPUT119), .B(n973), .ZN(n974) );
  NOR2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(n978), .B(KEYINPUT53), .ZN(n981) );
  XOR2_X1 U1073 ( .A(G2084), .B(G34), .Z(n979) );
  XNOR2_X1 U1074 ( .A(KEYINPUT54), .B(n979), .ZN(n980) );
  NAND2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(G35), .B(G2090), .ZN(n982) );
  NOR2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1078 ( .A(n985), .B(n984), .ZN(n986) );
  NAND2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1080 ( .A1(G11), .A2(n988), .ZN(n989) );
  XOR2_X1 U1081 ( .A(KEYINPUT121), .B(n989), .Z(n990) );
  NOR2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n1022) );
  NAND2_X1 U1084 ( .A1(G303), .A2(G1971), .ZN(n1002) );
  XOR2_X1 U1085 ( .A(G1956), .B(n994), .Z(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n1000) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(n1003), .B(KEYINPUT123), .ZN(n1011) );
  XOR2_X1 U1091 ( .A(n1004), .B(G1348), .Z(n1007) );
  XNOR2_X1 U1092 ( .A(n1005), .B(G1341), .ZN(n1006) );
  NAND2_X1 U1093 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  XNOR2_X1 U1094 ( .A(G1961), .B(G301), .ZN(n1008) );
  NOR2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1096 ( .A1(n1011), .A2(n1010), .ZN(n1017) );
  XOR2_X1 U1097 ( .A(G168), .B(G1966), .Z(n1012) );
  NOR2_X1 U1098 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1099 ( .A(KEYINPUT122), .B(n1014), .Z(n1015) );
  XOR2_X1 U1100 ( .A(KEYINPUT57), .B(n1015), .Z(n1016) );
  NOR2_X1 U1101 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  XOR2_X1 U1102 ( .A(G16), .B(KEYINPUT56), .Z(n1018) );
  NOR2_X1 U1103 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1104 ( .A(n1020), .B(KEYINPUT124), .ZN(n1021) );
  NOR2_X1 U1105 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1106 ( .A(KEYINPUT62), .B(n1023), .ZN(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

