//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 0 1 1 0 1 0 1 0 0 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G210), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n189), .B(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT26), .B(G101), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n193), .B(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT28), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G143), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  OR2_X1    g016(.A1(KEYINPUT0), .A2(G128), .ZN(new_n203));
  NAND2_X1  g017(.A1(KEYINPUT0), .A2(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(G143), .B(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(new_n204), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  INV_X1    g024(.A(G137), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT64), .B1(new_n211), .B2(G134), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n213));
  INV_X1    g027(.A(G134), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(G137), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n211), .A2(KEYINPUT11), .A3(G134), .ZN(new_n217));
  AOI21_X1  g031(.A(KEYINPUT11), .B1(new_n211), .B2(G134), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n210), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT11), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n221), .B1(new_n214), .B2(G137), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n211), .A2(KEYINPUT11), .A3(G134), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n222), .A2(new_n212), .A3(new_n215), .A4(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(G131), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n209), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT65), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n216), .A2(new_n219), .A3(new_n210), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n214), .A2(G137), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n211), .A2(G134), .ZN(new_n230));
  OAI21_X1  g044(.A(G131), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G128), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT1), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n233), .B1(G143), .B2(new_n198), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n232), .B1(new_n234), .B2(KEYINPUT66), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n199), .A2(KEYINPUT1), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n207), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n207), .A2(new_n233), .A3(G128), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n228), .B(new_n231), .C1(new_n239), .C2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n224), .A2(G131), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n228), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT65), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n245), .A3(new_n209), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n227), .A2(new_n242), .A3(new_n246), .ZN(new_n247));
  XOR2_X1   g061(.A(G116), .B(G119), .Z(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT2), .B(G113), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XOR2_X1   g064(.A(KEYINPUT2), .B(G113), .Z(new_n251));
  XNOR2_X1  g065(.A(G116), .B(G119), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n250), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n248), .A2(KEYINPUT67), .A3(new_n249), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n247), .A2(new_n257), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n199), .A2(new_n201), .B1(new_n203), .B2(new_n204), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n199), .A2(new_n201), .A3(new_n204), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT68), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n206), .A2(new_n262), .A3(new_n208), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n261), .B(new_n263), .C1(new_n220), .C2(new_n225), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n242), .A2(new_n264), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n255), .A2(KEYINPUT69), .A3(new_n256), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT69), .B1(new_n255), .B2(new_n256), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n197), .B1(new_n258), .B2(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT28), .B1(new_n265), .B2(new_n268), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n196), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT30), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n247), .A2(new_n273), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n242), .A2(new_n264), .A3(KEYINPUT30), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n274), .A2(new_n257), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT31), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n277), .A2(new_n278), .A3(new_n269), .A4(new_n195), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n272), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n269), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n275), .B1(new_n273), .B2(new_n247), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n281), .B1(new_n282), .B2(new_n257), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n278), .B1(new_n283), .B2(new_n195), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n187), .B(new_n188), .C1(new_n280), .C2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT32), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n283), .A2(new_n195), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT31), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(new_n279), .A3(new_n272), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n290), .A2(KEYINPUT32), .A3(new_n187), .A4(new_n188), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT71), .B1(new_n283), .B2(new_n195), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n277), .A2(new_n269), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT71), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(new_n295), .A3(new_n196), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT29), .ZN(new_n297));
  INV_X1    g111(.A(new_n271), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n258), .A2(new_n269), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n195), .B(new_n298), .C1(new_n299), .C2(new_n197), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n293), .A2(new_n296), .A3(new_n297), .A4(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n242), .A2(new_n264), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n302), .B1(new_n266), .B2(new_n267), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n269), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n271), .B1(new_n304), .B2(KEYINPUT28), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n196), .A2(new_n297), .ZN(new_n306));
  AOI21_X1  g120(.A(G902), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n292), .B1(new_n308), .B2(G472), .ZN(new_n309));
  AOI211_X1 g123(.A(KEYINPUT72), .B(new_n187), .C1(new_n301), .C2(new_n307), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n287), .B(new_n291), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G125), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n312), .A2(KEYINPUT16), .A3(G140), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  AND2_X1   g128(.A1(G125), .A2(G140), .ZN(new_n315));
  NOR2_X1   g129(.A1(G125), .A2(G140), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT16), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n314), .A2(new_n317), .A3(G146), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT74), .ZN(new_n319));
  XNOR2_X1  g133(.A(G125), .B(G140), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n313), .B1(new_n320), .B2(KEYINPUT16), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(G146), .ZN(new_n323));
  NOR3_X1   g137(.A1(new_n321), .A2(KEYINPUT75), .A3(G146), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n314), .A2(new_n317), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n325), .B1(new_n326), .B2(new_n198), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n319), .B(new_n323), .C1(new_n324), .C2(new_n327), .ZN(new_n328));
  XOR2_X1   g142(.A(KEYINPUT24), .B(G110), .Z(new_n329));
  XNOR2_X1  g143(.A(G119), .B(G128), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT23), .B1(new_n232), .B2(G119), .ZN(new_n332));
  INV_X1    g146(.A(G119), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT73), .B1(new_n333), .B2(G128), .ZN(new_n334));
  XOR2_X1   g148(.A(new_n332), .B(new_n334), .Z(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G110), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n328), .A2(new_n331), .A3(new_n336), .ZN(new_n337));
  OAI22_X1  g151(.A1(new_n335), .A2(G110), .B1(new_n330), .B2(new_n329), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n320), .A2(new_n198), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n318), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT76), .B(KEYINPUT22), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(G137), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n343), .B(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n345), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n337), .A2(new_n340), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n188), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT25), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n346), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n348), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G217), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n354), .B1(G234), .B2(new_n188), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  OR2_X1    g170(.A1(new_n349), .A2(new_n355), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(G110), .B(G140), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n191), .A2(G227), .ZN(new_n361));
  XOR2_X1   g175(.A(new_n360), .B(new_n361), .Z(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT78), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n244), .B(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n199), .A2(KEYINPUT66), .A3(KEYINPUT1), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G128), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n234), .A2(KEYINPUT66), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n202), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n366), .B1(new_n370), .B2(new_n240), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT77), .ZN(new_n372));
  INV_X1    g186(.A(G107), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n373), .A3(G104), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(KEYINPUT3), .ZN(new_n375));
  INV_X1    g189(.A(G101), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n373), .A2(G104), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n372), .A2(new_n379), .A3(new_n373), .A4(G104), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n375), .A2(new_n376), .A3(new_n378), .A4(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G104), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n382), .A2(G107), .ZN(new_n383));
  OAI21_X1  g197(.A(G101), .B1(new_n377), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n207), .B1(G128), .B2(new_n236), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n381), .B(new_n384), .C1(new_n241), .C2(new_n387), .ZN(new_n388));
  AOI22_X1  g202(.A1(new_n371), .A2(new_n386), .B1(new_n388), .B2(new_n366), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n375), .A2(new_n378), .A3(new_n380), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G101), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(KEYINPUT4), .A3(new_n381), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n390), .A2(new_n393), .A3(G101), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n392), .A2(new_n261), .A3(new_n263), .A4(new_n394), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n365), .A2(new_n389), .A3(new_n395), .ZN(new_n396));
  AOI22_X1  g210(.A1(new_n389), .A2(new_n395), .B1(new_n243), .B2(new_n228), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n363), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT80), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI211_X1 g214(.A(KEYINPUT80), .B(new_n363), .C1(new_n396), .C2(new_n397), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n385), .A2(new_n370), .A3(new_n240), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n388), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n244), .ZN(new_n404));
  NOR2_X1   g218(.A1(KEYINPUT79), .A2(KEYINPUT12), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(KEYINPUT79), .A2(KEYINPUT12), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n403), .B(new_n244), .C1(KEYINPUT79), .C2(KEYINPUT12), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n365), .A2(new_n389), .A3(new_n395), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n410), .A3(new_n362), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n400), .A2(new_n401), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G469), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n413), .A3(new_n188), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n362), .B1(new_n409), .B2(new_n410), .ZN(new_n415));
  NOR3_X1   g229(.A1(new_n396), .A2(new_n397), .A3(new_n363), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(G469), .B1(new_n417), .B2(G902), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G221), .ZN(new_n420));
  XOR2_X1   g234(.A(KEYINPUT9), .B(G234), .Z(new_n421));
  AOI21_X1  g235(.A(new_n420), .B1(new_n421), .B2(new_n188), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(G214), .B1(G237), .B2(G902), .ZN(new_n425));
  INV_X1    g239(.A(G952), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n426), .A2(KEYINPUT90), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n426), .A2(KEYINPUT90), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n191), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(G234), .B2(G237), .ZN(new_n430));
  XOR2_X1   g244(.A(KEYINPUT21), .B(G898), .Z(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AOI211_X1 g246(.A(new_n188), .B(new_n191), .C1(G234), .C2(G237), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n430), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n370), .A2(new_n312), .A3(new_n240), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT84), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n206), .A2(G125), .A3(new_n208), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT84), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n370), .A2(new_n439), .A3(new_n312), .A4(new_n240), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n437), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n191), .A2(G224), .ZN(new_n442));
  XOR2_X1   g256(.A(new_n442), .B(KEYINPUT81), .Z(new_n443));
  OR2_X1    g257(.A1(KEYINPUT85), .A2(KEYINPUT7), .ZN(new_n444));
  NAND2_X1  g258(.A1(KEYINPUT85), .A2(KEYINPUT7), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT7), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT86), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n447), .B1(new_n443), .B2(new_n448), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n436), .A2(new_n438), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n443), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT86), .ZN(new_n452));
  AOI22_X1  g266(.A1(new_n441), .A2(new_n446), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n257), .A2(new_n392), .A3(new_n394), .ZN(new_n454));
  XNOR2_X1  g268(.A(G110), .B(G122), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n381), .A2(new_n253), .A3(new_n384), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT5), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n333), .A3(G116), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G113), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n252), .A2(KEYINPUT5), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n454), .A2(new_n455), .A3(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n455), .B(KEYINPUT8), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n460), .A2(KEYINPUT82), .B1(KEYINPUT5), .B2(new_n252), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(KEYINPUT82), .B2(new_n460), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n467), .A2(new_n456), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n462), .A2(new_n253), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n469), .A2(new_n385), .ZN(new_n470));
  OAI211_X1 g284(.A(KEYINPUT83), .B(new_n465), .C1(new_n468), .C2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT83), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n467), .A2(new_n456), .B1(new_n385), .B2(new_n469), .ZN(new_n473));
  INV_X1    g287(.A(new_n465), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n453), .A2(new_n464), .A3(new_n471), .A4(new_n475), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n476), .A2(new_n188), .ZN(new_n477));
  OAI21_X1  g291(.A(G210), .B1(G237), .B2(G902), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n454), .A2(new_n463), .ZN(new_n479));
  INV_X1    g293(.A(new_n455), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(KEYINPUT6), .A3(new_n464), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT6), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n479), .A2(new_n483), .A3(new_n480), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n436), .A2(new_n438), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(new_n451), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n477), .A2(new_n478), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n478), .B1(new_n477), .B2(new_n487), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n425), .B(new_n435), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n190), .A2(new_n191), .A3(G214), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(G143), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(KEYINPUT17), .A3(G131), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT87), .B1(new_n328), .B2(new_n496), .ZN(new_n497));
  OR2_X1    g311(.A1(new_n324), .A2(new_n327), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n319), .A2(new_n323), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT87), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n498), .A2(new_n499), .A3(new_n500), .A4(new_n495), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n494), .A2(G131), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n493), .A2(new_n210), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n497), .B(new_n501), .C1(KEYINPUT17), .C2(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(G113), .B(G122), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(new_n382), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT18), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n493), .B1(new_n508), .B2(new_n210), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n320), .B(new_n198), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n509), .B(new_n510), .C1(new_n502), .C2(new_n508), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n505), .A2(new_n507), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n507), .B1(new_n505), .B2(new_n511), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n188), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(G475), .ZN(new_n516));
  INV_X1    g330(.A(G116), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(G122), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT88), .B1(new_n518), .B2(KEYINPUT14), .ZN(new_n519));
  INV_X1    g333(.A(G122), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G116), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n518), .A2(KEYINPUT14), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT88), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT14), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n523), .A2(new_n524), .A3(new_n517), .A4(G122), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n519), .A2(new_n521), .A3(new_n522), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G107), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n521), .A2(new_n518), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n373), .ZN(new_n529));
  XNOR2_X1  g343(.A(G128), .B(G143), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n214), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n530), .A2(new_n214), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n527), .B(new_n529), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n528), .B(new_n373), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n530), .A2(KEYINPUT13), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n200), .A2(G128), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n536), .B(G134), .C1(KEYINPUT13), .C2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n535), .A2(new_n531), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n421), .A2(G217), .A3(new_n191), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n541), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n534), .A2(new_n539), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(G902), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT89), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT15), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n548), .A3(G478), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(G478), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n545), .A2(new_n546), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT20), .ZN(new_n554));
  INV_X1    g368(.A(new_n504), .ZN(new_n555));
  XOR2_X1   g369(.A(new_n320), .B(KEYINPUT19), .Z(new_n556));
  OAI21_X1  g370(.A(new_n318), .B1(new_n556), .B2(G146), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n511), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n507), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n512), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(G475), .A2(G902), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n554), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n562), .ZN(new_n564));
  AOI211_X1 g378(.A(KEYINPUT20), .B(new_n564), .C1(new_n512), .C2(new_n560), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n516), .B(new_n553), .C1(new_n563), .C2(new_n565), .ZN(new_n566));
  NOR3_X1   g380(.A1(new_n424), .A2(new_n491), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n311), .A2(new_n359), .A3(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(G101), .ZN(G3));
  INV_X1    g383(.A(KEYINPUT33), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT91), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n534), .A2(new_n539), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n571), .B1(new_n534), .B2(new_n539), .ZN(new_n574));
  OAI211_X1 g388(.A(KEYINPUT92), .B(new_n541), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n575), .A2(new_n544), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n540), .A2(KEYINPUT91), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n572), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n541), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT92), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n570), .B1(new_n576), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n542), .A2(new_n570), .A3(new_n544), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  OAI211_X1 g398(.A(G478), .B(new_n188), .C1(new_n582), .C2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n545), .A2(G478), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(KEYINPUT93), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n516), .B1(new_n563), .B2(new_n565), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(new_n491), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n424), .A2(new_n358), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n188), .B1(new_n280), .B2(new_n284), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(G472), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n285), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n592), .A2(new_n593), .A3(new_n597), .ZN(new_n598));
  XOR2_X1   g412(.A(KEYINPUT34), .B(G104), .Z(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(G6));
  NAND2_X1  g414(.A1(new_n561), .A2(new_n562), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT20), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n561), .A2(new_n554), .A3(new_n562), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(KEYINPUT94), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT94), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n565), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n604), .A2(new_n516), .A3(new_n552), .A4(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n607), .A2(new_n491), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n608), .A2(new_n597), .A3(new_n593), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT35), .B(G107), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G9));
  INV_X1    g425(.A(new_n355), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(new_n351), .B2(new_n352), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n345), .A2(KEYINPUT36), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n341), .B(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(new_n188), .A3(new_n612), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT95), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(KEYINPUT95), .B1(new_n613), .B2(new_n617), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n597), .A2(KEYINPUT96), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT96), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n619), .B1(new_n356), .B2(new_n616), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n613), .A2(new_n617), .A3(KEYINPUT95), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n624), .B1(new_n627), .B2(new_n596), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n623), .A2(new_n628), .A3(new_n567), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT37), .ZN(new_n630));
  XOR2_X1   g444(.A(new_n630), .B(G110), .Z(G12));
  INV_X1    g445(.A(new_n430), .ZN(new_n632));
  INV_X1    g446(.A(G900), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n433), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n607), .A2(new_n424), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n425), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n487), .A2(new_n188), .A3(new_n476), .ZN(new_n639));
  INV_X1    g453(.A(new_n478), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n638), .B1(new_n641), .B2(new_n488), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n627), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n311), .A2(new_n637), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G128), .ZN(G30));
  NAND2_X1  g460(.A1(new_n641), .A2(new_n488), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT38), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n638), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n195), .B1(new_n269), .B2(new_n303), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n651), .A2(KEYINPUT97), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(KEYINPUT97), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n288), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(G472), .B1(new_n654), .B2(G902), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n291), .A2(new_n287), .A3(new_n655), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n656), .A2(new_n618), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n590), .A2(new_n552), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n650), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT98), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n635), .B(KEYINPUT39), .Z(new_n663));
  OAI21_X1  g477(.A(KEYINPUT40), .B1(new_n424), .B2(new_n663), .ZN(new_n664));
  OR3_X1    g478(.A1(new_n424), .A2(KEYINPUT40), .A3(new_n663), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n662), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G143), .ZN(G45));
  INV_X1    g481(.A(KEYINPUT99), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n589), .A2(new_n590), .A3(new_n635), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n668), .B1(new_n669), .B2(new_n643), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n602), .A2(new_n603), .B1(G475), .B2(new_n515), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n575), .A2(new_n544), .ZN(new_n672));
  AOI21_X1  g486(.A(KEYINPUT92), .B1(new_n578), .B2(new_n541), .ZN(new_n673));
  OAI21_X1  g487(.A(KEYINPUT33), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(G902), .B1(new_n674), .B2(new_n583), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n587), .B1(new_n675), .B2(G478), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n677), .A2(KEYINPUT99), .A3(new_n642), .A4(new_n635), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n627), .A2(new_n424), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n311), .A2(new_n670), .A3(new_n678), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G146), .ZN(G48));
  NAND2_X1  g495(.A1(new_n412), .A2(new_n188), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(G469), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n683), .A2(new_n423), .A3(new_n414), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n311), .A2(new_n359), .A3(new_n592), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT41), .B(G113), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G15));
  NAND4_X1  g502(.A1(new_n311), .A2(new_n359), .A3(new_n608), .A4(new_n685), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G116), .ZN(G18));
  NOR3_X1   g504(.A1(new_n684), .A2(new_n566), .A3(new_n434), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n311), .A2(new_n644), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G119), .ZN(G21));
  NOR2_X1   g507(.A1(new_n658), .A2(new_n643), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n358), .B(KEYINPUT100), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n684), .A2(new_n434), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n279), .B1(new_n305), .B2(new_n195), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n187), .B(new_n188), .C1(new_n697), .C2(new_n284), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n595), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n694), .A2(new_n695), .A3(new_n696), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G122), .ZN(G24));
  INV_X1    g515(.A(new_n669), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n356), .A2(new_n616), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n595), .A2(new_n703), .A3(new_n698), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n702), .A2(new_n705), .A3(new_n642), .A4(new_n685), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT101), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n312), .ZN(G27));
  NOR4_X1   g522(.A1(new_n489), .A2(new_n490), .A3(new_n638), .A4(new_n422), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n396), .A2(new_n397), .ZN(new_n710));
  OAI21_X1  g524(.A(KEYINPUT103), .B1(new_n710), .B2(new_n363), .ZN(new_n711));
  INV_X1    g525(.A(new_n415), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT103), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n416), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n711), .A2(new_n712), .A3(G469), .A4(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(G469), .A2(G902), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT102), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n414), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n709), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n311), .A2(new_n359), .A3(new_n719), .A4(new_n702), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT42), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n308), .A2(G472), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(KEYINPUT72), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n308), .A2(new_n292), .A3(G472), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n291), .A2(KEYINPUT104), .ZN(new_n727));
  OR2_X1    g541(.A1(new_n291), .A2(KEYINPUT104), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n726), .A2(new_n287), .A3(new_n727), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n709), .A2(new_n718), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n730), .A2(new_n721), .A3(new_n669), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(new_n695), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n722), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G131), .ZN(G33));
  NOR2_X1   g548(.A1(new_n607), .A2(new_n636), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n311), .A2(new_n359), .A3(new_n719), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G134), .ZN(G36));
  NAND4_X1  g551(.A1(new_n711), .A2(new_n712), .A3(KEYINPUT45), .A4(new_n714), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT45), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n739), .B1(new_n415), .B2(new_n416), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n738), .A2(G469), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n717), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT46), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n741), .A2(KEYINPUT46), .A3(new_n717), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n744), .A2(new_n414), .A3(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n663), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n423), .A3(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT43), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n750), .B1(new_n590), .B2(new_n676), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n589), .A2(new_n671), .A3(KEYINPUT43), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n596), .A3(new_n703), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n748), .B1(new_n749), .B2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n753), .A2(KEYINPUT44), .A3(new_n596), .A4(new_n703), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n647), .A2(new_n638), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(KEYINPUT105), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G137), .ZN(G39));
  NAND2_X1  g575(.A1(new_n746), .A2(new_n423), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT47), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n746), .A2(KEYINPUT47), .A3(new_n423), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n669), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NOR4_X1   g580(.A1(new_n311), .A2(new_n359), .A3(new_n638), .A4(new_n647), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(KEYINPUT106), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G140), .ZN(G42));
  AND4_X1   g584(.A1(new_n686), .A2(new_n689), .A3(new_n692), .A4(new_n700), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n771), .A2(KEYINPUT53), .A3(new_n733), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n658), .A2(new_n643), .A3(new_n636), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n657), .A2(new_n423), .A3(new_n718), .A4(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n774), .A2(new_n680), .A3(new_n645), .A4(new_n706), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR4_X1   g591(.A1(new_n669), .A2(new_n704), .A3(new_n684), .A4(new_n643), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n622), .A2(new_n642), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n291), .A2(new_n287), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n779), .B1(new_n726), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n778), .B1(new_n781), .B2(new_n637), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n782), .A2(KEYINPUT52), .A3(new_n680), .A4(new_n774), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n777), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT108), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n785), .B1(new_n671), .B2(new_n676), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n589), .A2(new_n590), .A3(KEYINPUT108), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI211_X1 g602(.A(new_n638), .B(new_n434), .C1(new_n641), .C2(new_n488), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n788), .A2(new_n789), .A3(new_n597), .A4(new_n593), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n789), .A2(KEYINPUT109), .A3(new_n671), .A4(new_n552), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT109), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n516), .B(new_n552), .C1(new_n563), .C2(new_n565), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n792), .B1(new_n491), .B2(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n791), .A2(new_n794), .A3(new_n593), .A4(new_n597), .ZN(new_n795));
  AND4_X1   g609(.A1(new_n568), .A2(new_n629), .A3(new_n790), .A4(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n604), .A2(new_n516), .A3(new_n606), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n641), .A2(new_n425), .A3(new_n488), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n553), .A2(new_n635), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n311), .A2(new_n679), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT110), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n311), .A2(KEYINPUT110), .A3(new_n800), .A4(new_n679), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n719), .A2(new_n702), .A3(new_n705), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n736), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n796), .A2(new_n805), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n772), .A2(new_n784), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT112), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT112), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n772), .A2(new_n784), .A3(new_n809), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n777), .A2(new_n783), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n807), .B1(new_n803), .B2(new_n804), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n817), .A2(new_n733), .A3(new_n771), .A4(new_n796), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n815), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT111), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT111), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n821), .B(new_n815), .C1(new_n816), .C2(new_n818), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n814), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n796), .A2(new_n805), .A3(new_n808), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT113), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n817), .A2(new_n828), .A3(new_n796), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n827), .A2(new_n772), .A3(new_n829), .A4(new_n784), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n819), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  AOI22_X1  g646(.A1(new_n823), .A2(KEYINPUT54), .B1(new_n825), .B2(new_n832), .ZN(new_n833));
  AND4_X1   g647(.A1(new_n430), .A2(new_n753), .A3(new_n695), .A4(new_n699), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n834), .A2(new_n642), .A3(new_n685), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n834), .A2(new_n638), .A3(new_n649), .A4(new_n685), .ZN(new_n837));
  XOR2_X1   g651(.A(new_n837), .B(KEYINPUT50), .Z(new_n838));
  NAND2_X1  g652(.A1(new_n764), .A2(new_n765), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n683), .A2(new_n414), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n423), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n757), .B(new_n834), .C1(new_n839), .C2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n709), .A2(new_n430), .A3(new_n414), .A4(new_n683), .ZN(new_n843));
  OR3_X1    g657(.A1(new_n843), .A2(new_n358), .A3(new_n656), .ZN(new_n844));
  OR3_X1    g658(.A1(new_n844), .A2(new_n590), .A3(new_n589), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n843), .B1(new_n751), .B2(new_n752), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n705), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n838), .A2(new_n842), .A3(new_n845), .A4(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT51), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n429), .B1(new_n848), .B2(new_n849), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n844), .A2(new_n591), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n729), .A2(new_n695), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n846), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT48), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n850), .A2(new_n851), .A3(new_n852), .A4(new_n855), .ZN(new_n856));
  OAI22_X1  g670(.A1(new_n836), .A2(new_n856), .B1(G952), .B2(G953), .ZN(new_n857));
  OR3_X1    g671(.A1(new_n840), .A2(KEYINPUT107), .A3(KEYINPUT49), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n840), .B1(KEYINPUT107), .B2(KEYINPUT49), .ZN(new_n859));
  AOI211_X1 g673(.A(new_n638), .B(new_n422), .C1(KEYINPUT107), .C2(KEYINPUT49), .ZN(new_n860));
  AND4_X1   g674(.A1(new_n695), .A2(new_n858), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(new_n671), .A3(new_n589), .A4(new_n649), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n857), .B1(new_n656), .B2(new_n862), .ZN(G75));
  NOR2_X1   g677(.A1(new_n832), .A2(new_n188), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT56), .B1(new_n864), .B2(G210), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n482), .A2(new_n484), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n866), .B(new_n486), .Z(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT55), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  OR3_X1    g683(.A1(new_n865), .A2(KEYINPUT115), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n191), .A2(G952), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(new_n865), .B2(KEYINPUT115), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n869), .B1(new_n865), .B2(KEYINPUT115), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n870), .A2(new_n872), .A3(new_n873), .ZN(G51));
  NAND2_X1  g688(.A1(new_n831), .A2(new_n824), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n819), .A2(new_n830), .A3(new_n825), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n831), .A2(KEYINPUT116), .A3(new_n824), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n717), .B(KEYINPUT57), .Z(new_n880));
  NAND3_X1  g694(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n412), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n741), .B(KEYINPUT117), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n864), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n871), .B1(new_n882), .B2(new_n884), .ZN(G54));
  AND3_X1   g699(.A1(new_n864), .A2(KEYINPUT58), .A3(G475), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n886), .A2(new_n561), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n886), .A2(new_n561), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n887), .A2(new_n888), .A3(new_n871), .ZN(G60));
  NOR2_X1   g703(.A1(new_n582), .A2(new_n584), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n823), .A2(KEYINPUT54), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n877), .ZN(new_n893));
  XNOR2_X1  g707(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n894));
  NAND2_X1  g708(.A1(G478), .A2(G902), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n894), .B(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n891), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n878), .A2(new_n891), .A3(new_n879), .A4(new_n897), .ZN(new_n899));
  INV_X1    g713(.A(new_n871), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(KEYINPUT119), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n890), .B1(new_n833), .B2(new_n896), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT119), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n903), .A2(new_n904), .A3(new_n900), .A4(new_n899), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n902), .A2(new_n905), .ZN(G63));
  NAND2_X1  g720(.A1(G217), .A2(G902), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT120), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT60), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n831), .A2(new_n615), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n900), .ZN(new_n911));
  AOI22_X1  g725(.A1(new_n831), .A2(new_n909), .B1(new_n348), .B2(new_n346), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n911), .B1(new_n912), .B2(KEYINPUT122), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n913), .B(KEYINPUT61), .C1(KEYINPUT122), .C2(new_n912), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT61), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n915), .B1(new_n911), .B2(new_n912), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT121), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n914), .A2(new_n918), .A3(new_n919), .ZN(G66));
  AOI21_X1  g734(.A(new_n191), .B1(new_n431), .B2(G224), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n771), .A2(new_n796), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n921), .B1(new_n922), .B2(new_n191), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n866), .B1(G898), .B2(new_n191), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n923), .B(new_n924), .Z(G69));
  XOR2_X1   g739(.A(new_n282), .B(new_n556), .Z(new_n926));
  AOI22_X1  g740(.A1(new_n766), .A2(new_n767), .B1(new_n755), .B2(new_n758), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n786), .A2(new_n787), .A3(new_n793), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n424), .A2(new_n663), .A3(new_n798), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n311), .A2(new_n928), .A3(new_n359), .A4(new_n929), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT123), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n680), .A2(new_n645), .A3(new_n706), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n666), .A2(KEYINPUT62), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT62), .B1(new_n666), .B2(new_n932), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n927), .B(new_n931), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n926), .B1(new_n935), .B2(new_n191), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n932), .A2(new_n736), .ZN(new_n937));
  INV_X1    g751(.A(new_n748), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n853), .A2(new_n694), .A3(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n927), .A2(new_n937), .A3(new_n733), .A4(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n926), .B1(new_n940), .B2(G953), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(G900), .B2(G953), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n191), .B1(G227), .B2(G900), .ZN(new_n944));
  OAI22_X1  g758(.A1(new_n936), .A2(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n943), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT125), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n945), .B(new_n947), .ZN(G72));
  NAND2_X1  g762(.A1(G472), .A2(G902), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT63), .Z(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n935), .B2(new_n922), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n951), .A2(new_n294), .A3(new_n195), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n293), .A2(new_n296), .A3(new_n288), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n823), .A2(new_n953), .A3(new_n950), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n950), .B1(new_n940), .B2(new_n922), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n955), .A2(new_n283), .A3(new_n196), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n900), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(KEYINPUT126), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT126), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n956), .A2(new_n959), .A3(new_n900), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n952), .A2(new_n954), .A3(new_n958), .A4(new_n960), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT127), .ZN(G57));
endmodule


