//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 0 0 1 0 0 0 0 0 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n565, new_n566, new_n567,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n624, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1099, new_n1100;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT64), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  OR2_X1    g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NAND2_X1  g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G137), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  AND3_X1   g040(.A1(new_n465), .A2(KEYINPUT65), .A3(G101), .ZN(new_n466));
  AOI21_X1  g041(.A(KEYINPUT65), .B1(new_n465), .B2(G101), .ZN(new_n467));
  OAI22_X1  g042(.A1(new_n462), .A2(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n460), .A2(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n461), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OR2_X1    g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  OR2_X1    g048(.A1(G100), .A2(G2105), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n474), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n475));
  XOR2_X1   g050(.A(new_n475), .B(KEYINPUT67), .Z(new_n476));
  NAND2_X1  g051(.A1(new_n460), .A2(G2105), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT66), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  INV_X1    g054(.A(new_n462), .ZN(new_n480));
  AOI211_X1 g055(.A(new_n476), .B(new_n479), .C1(G136), .C2(new_n480), .ZN(G162));
  INV_X1    g056(.A(KEYINPUT71), .ZN(new_n482));
  INV_X1    g057(.A(G138), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  NOR2_X1   g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  AND2_X1   g061(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n484), .B(new_n485), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT70), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n461), .A2(G138), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(new_n458), .B2(new_n459), .ZN(new_n491));
  OAI21_X1  g066(.A(KEYINPUT4), .B1(new_n491), .B2(KEYINPUT68), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n484), .B(KEYINPUT68), .C1(new_n486), .C2(new_n487), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT69), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n484), .B1(new_n487), .B2(new_n486), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n485), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n498), .A2(new_n499), .A3(new_n493), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n489), .B1(new_n495), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n460), .A2(G126), .A3(G2105), .ZN(new_n502));
  OR2_X1    g077(.A1(G102), .A2(G2105), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n503), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n482), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n507));
  XNOR2_X1  g082(.A(new_n488), .B(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n496), .A2(new_n497), .ZN(new_n509));
  AND4_X1   g084(.A1(new_n499), .A2(new_n509), .A3(KEYINPUT4), .A4(new_n493), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n499), .B1(new_n498), .B2(new_n493), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n508), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n505), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(KEYINPUT71), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n506), .A2(new_n514), .ZN(G164));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT5), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n517), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n519), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n518), .A2(new_n520), .B1(new_n517), .B2(G543), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(KEYINPUT74), .A3(G62), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  XOR2_X1   g098(.A(new_n523), .B(KEYINPUT75), .Z(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g100(.A(KEYINPUT74), .B1(new_n521), .B2(G62), .ZN(new_n526));
  OAI21_X1  g101(.A(G651), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT72), .ZN(new_n528));
  INV_X1    g103(.A(G651), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n529), .B2(KEYINPUT6), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT6), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n531), .A2(KEYINPUT72), .A3(G651), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n530), .A2(new_n532), .B1(KEYINPUT6), .B2(new_n529), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n521), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n533), .A2(G543), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n535), .A2(G88), .B1(new_n536), .B2(G50), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n527), .A2(new_n537), .ZN(G303));
  INV_X1    g113(.A(G303), .ZN(G166));
  NAND2_X1  g114(.A1(new_n535), .A2(G89), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n536), .A2(G51), .ZN(new_n541));
  AND2_X1   g116(.A1(G63), .A2(G651), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT7), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n543), .A2(KEYINPUT7), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n521), .A2(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n540), .A2(new_n541), .A3(new_n546), .ZN(G286));
  INV_X1    g122(.A(G286), .ZN(G168));
  AOI22_X1  g123(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT76), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g126(.A(G651), .B1(new_n549), .B2(new_n550), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n535), .A2(G90), .B1(new_n536), .B2(G52), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(G301));
  INV_X1    g130(.A(G301), .ZN(G171));
  AOI22_X1  g131(.A1(new_n535), .A2(G81), .B1(new_n536), .B2(G43), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n557), .B(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n560), .A2(new_n529), .ZN(new_n561));
  AND2_X1   g136(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g139(.A(KEYINPUT78), .B(KEYINPUT8), .Z(new_n565));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n565), .B(new_n566), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n518), .A2(new_n520), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n517), .A2(G543), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n569), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT79), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n576));
  OAI211_X1 g151(.A(new_n576), .B(new_n569), .C1(new_n572), .C2(new_n573), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(G651), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(KEYINPUT80), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT80), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n575), .A2(new_n580), .A3(G651), .A4(new_n577), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n533), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G53), .ZN(new_n584));
  OR3_X1    g159(.A1(new_n583), .A2(KEYINPUT9), .A3(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT9), .B1(new_n583), .B2(new_n584), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n585), .A2(new_n586), .B1(G91), .B2(new_n535), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n582), .A2(new_n587), .ZN(G299));
  OAI21_X1  g163(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n589));
  INV_X1    g164(.A(G49), .ZN(new_n590));
  INV_X1    g165(.A(G87), .ZN(new_n591));
  OAI221_X1 g166(.A(new_n589), .B1(new_n583), .B2(new_n590), .C1(new_n591), .C2(new_n534), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT81), .ZN(G288));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT82), .ZN(new_n595));
  INV_X1    g170(.A(G61), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n572), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G651), .B1(new_n536), .B2(G48), .ZN(new_n598));
  INV_X1    g173(.A(G86), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(new_n534), .ZN(G305));
  INV_X1    g175(.A(G85), .ZN(new_n601));
  INV_X1    g176(.A(G47), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n534), .A2(new_n601), .B1(new_n583), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(new_n529), .ZN(new_n605));
  OR3_X1    g180(.A1(new_n603), .A2(new_n605), .A3(KEYINPUT83), .ZN(new_n606));
  OAI21_X1  g181(.A(KEYINPUT83), .B1(new_n603), .B2(new_n605), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(G290));
  NAND2_X1  g183(.A1(G301), .A2(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n535), .A2(G92), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT10), .Z(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n572), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n614), .A2(G651), .B1(new_n536), .B2(G54), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n609), .B1(new_n617), .B2(G868), .ZN(G284));
  OAI21_X1  g193(.A(new_n609), .B1(new_n617), .B2(G868), .ZN(G321));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  INV_X1    g195(.A(G299), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G297));
  OAI21_X1  g197(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G280));
  XNOR2_X1  g198(.A(KEYINPUT84), .B(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n617), .B1(G860), .B2(new_n624), .ZN(G148));
  NAND2_X1  g200(.A1(new_n617), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G868), .B2(new_n562), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g204(.A1(new_n460), .A2(new_n465), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n478), .A2(G123), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n480), .A2(G135), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n636), .A2(KEYINPUT85), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(KEYINPUT85), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(G111), .B2(new_n461), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n634), .B(new_n635), .C1(new_n637), .C2(new_n639), .ZN(new_n640));
  AOI22_X1  g215(.A1(new_n633), .A2(G2100), .B1(G2096), .B2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(G2100), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n632), .A2(new_n642), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n641), .B(new_n643), .C1(G2096), .C2(new_n640), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT86), .ZN(G156));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT89), .ZN(new_n647));
  XOR2_X1   g222(.A(KEYINPUT88), .B(G2438), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2430), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(new_n652), .A3(KEYINPUT14), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT90), .ZN(new_n654));
  XOR2_X1   g229(.A(G2451), .B(G2454), .Z(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n654), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT87), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1341), .B(G1348), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT91), .ZN(new_n663));
  INV_X1    g238(.A(G14), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n660), .B2(new_n661), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(G401));
  XNOR2_X1  g242(.A(G2072), .B(G2078), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT17), .Z(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(new_n670), .B2(new_n668), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT92), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n673), .A2(new_n670), .A3(new_n668), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT18), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n674), .A2(new_n670), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n679), .B1(new_n669), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(new_n642), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT93), .B(G2096), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(G1971), .B(G1976), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1956), .B(G2474), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1961), .B(G1966), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NOR3_X1   g266(.A1(new_n687), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n687), .A2(new_n690), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT20), .Z(new_n694));
  AOI211_X1 g269(.A(new_n692), .B(new_n694), .C1(new_n687), .C2(new_n691), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1981), .B(G1986), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(G229));
  MUX2_X1   g276(.A(G6), .B(G305), .S(G16), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT95), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT32), .B(G1981), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  MUX2_X1   g280(.A(G23), .B(new_n592), .S(G16), .Z(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT33), .B(G1976), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT97), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT96), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n706), .B(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G1971), .ZN(new_n711));
  NAND2_X1  g286(.A1(G166), .A2(G16), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G16), .B2(G22), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n710), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n711), .B2(new_n713), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n705), .A2(new_n715), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n716), .A2(KEYINPUT34), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(KEYINPUT34), .ZN(new_n718));
  INV_X1    g293(.A(G24), .ZN(new_n719));
  OR3_X1    g294(.A1(new_n719), .A2(KEYINPUT94), .A3(G16), .ZN(new_n720));
  OAI21_X1  g295(.A(KEYINPUT94), .B1(new_n719), .B2(G16), .ZN(new_n721));
  INV_X1    g296(.A(G290), .ZN(new_n722));
  INV_X1    g297(.A(G16), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n720), .B(new_n721), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G1986), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n478), .A2(G119), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n480), .A2(G131), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n461), .A2(G107), .ZN(new_n728));
  OAI21_X1  g303(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n726), .B(new_n727), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  MUX2_X1   g305(.A(G25), .B(new_n730), .S(G29), .Z(new_n731));
  XOR2_X1   g306(.A(KEYINPUT35), .B(G1991), .Z(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n731), .B(new_n733), .ZN(new_n734));
  NOR4_X1   g309(.A1(new_n717), .A2(new_n718), .A3(new_n725), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT98), .B(KEYINPUT36), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT102), .B(KEYINPUT23), .Z(new_n738));
  NAND2_X1  g313(.A1(new_n723), .A2(G20), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n621), .B2(new_n723), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT103), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1956), .ZN(new_n743));
  NAND2_X1  g318(.A1(G162), .A2(G29), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G29), .B2(G35), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT29), .B(G2090), .Z(new_n746));
  NOR2_X1   g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G29), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G26), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT28), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n478), .A2(G128), .ZN(new_n751));
  OAI21_X1  g326(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n752));
  INV_X1    g327(.A(G116), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(G2105), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n480), .B2(G140), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n750), .B1(new_n756), .B2(G29), .ZN(new_n757));
  INV_X1    g332(.A(G2067), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(G34), .ZN(new_n760));
  AOI21_X1  g335(.A(G29), .B1(new_n760), .B2(KEYINPUT24), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(KEYINPUT99), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(KEYINPUT99), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(KEYINPUT24), .B2(new_n760), .ZN(new_n764));
  OAI22_X1  g339(.A1(new_n472), .A2(new_n748), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G2084), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT25), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n460), .A2(G127), .ZN(new_n773));
  NAND2_X1  g348(.A1(G115), .A2(G2104), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n461), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AOI211_X1 g350(.A(new_n772), .B(new_n775), .C1(G139), .C2(new_n480), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n776), .A2(new_n748), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n748), .B2(G33), .ZN(new_n778));
  INV_X1    g353(.A(G2072), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n767), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n765), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n780), .B1(G2084), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT30), .B(G28), .ZN(new_n783));
  OR2_X1    g358(.A1(KEYINPUT31), .A2(G11), .ZN(new_n784));
  NAND2_X1  g359(.A1(KEYINPUT31), .A2(G11), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n783), .A2(new_n748), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI221_X1 g361(.A(new_n786), .B1(new_n640), .B2(new_n748), .C1(new_n778), .C2(new_n779), .ZN(new_n787));
  NOR4_X1   g362(.A1(new_n747), .A2(new_n759), .A3(new_n782), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n562), .A2(G16), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G16), .B2(G19), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n788), .B1(G1341), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n723), .A2(G21), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G168), .B2(new_n723), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1966), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n748), .A2(G32), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n478), .A2(G129), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n480), .A2(G141), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT100), .B(KEYINPUT26), .ZN(new_n799));
  NAND3_X1  g374(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G105), .B2(new_n465), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n797), .A2(new_n798), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n796), .B1(new_n803), .B2(G29), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT27), .B(G1996), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT101), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n745), .A2(new_n746), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n804), .B2(new_n806), .ZN(new_n808));
  NOR2_X1   g383(.A1(G4), .A2(G16), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n617), .B2(G16), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1348), .ZN(new_n811));
  NOR4_X1   g386(.A1(new_n792), .A2(new_n795), .A3(new_n808), .A4(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(G27), .A2(G29), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G164), .B2(G29), .ZN(new_n814));
  INV_X1    g389(.A(G2078), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n723), .A2(G5), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G171), .B2(new_n723), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(G1961), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n791), .B2(G1341), .ZN(new_n820));
  AND4_X1   g395(.A1(new_n743), .A2(new_n812), .A3(new_n816), .A4(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n735), .A2(KEYINPUT98), .A3(KEYINPUT36), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n737), .A2(new_n821), .A3(new_n822), .ZN(G150));
  INV_X1    g398(.A(G150), .ZN(G311));
  INV_X1    g399(.A(G93), .ZN(new_n825));
  INV_X1    g400(.A(G55), .ZN(new_n826));
  OAI22_X1  g401(.A1(new_n534), .A2(new_n825), .B1(new_n583), .B2(new_n826), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n828), .A2(new_n529), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT105), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G860), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT37), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n617), .A2(G559), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n562), .A2(new_n830), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n559), .A2(new_n561), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(new_n831), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n836), .B(new_n840), .Z(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  AND2_X1   g417(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n843));
  INV_X1    g418(.A(G860), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n842), .B2(KEYINPUT39), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n833), .B1(new_n843), .B2(new_n845), .ZN(G145));
  NAND2_X1  g421(.A1(new_n480), .A2(G142), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n461), .A2(G118), .ZN(new_n848));
  OAI21_X1  g423(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(G130), .B2(new_n478), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(new_n631), .Z(new_n852));
  XOR2_X1   g427(.A(new_n803), .B(new_n776), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n505), .B(KEYINPUT107), .Z(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(new_n512), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n756), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n730), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n854), .B(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(G162), .B(G160), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n640), .B(KEYINPUT106), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(G37), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n862), .B2(new_n859), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g440(.A(G290), .B(G305), .ZN(new_n866));
  XNOR2_X1  g441(.A(G303), .B(new_n592), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT108), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n868), .B1(new_n869), .B2(KEYINPUT42), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(KEYINPUT42), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n840), .B(new_n626), .ZN(new_n873));
  XNOR2_X1  g448(.A(G299), .B(new_n616), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(KEYINPUT41), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n875), .B1(new_n876), .B2(new_n873), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n872), .B(new_n877), .ZN(new_n878));
  MUX2_X1   g453(.A(new_n831), .B(new_n878), .S(G868), .Z(G295));
  MUX2_X1   g454(.A(new_n831), .B(new_n878), .S(G868), .Z(G331));
  XNOR2_X1  g455(.A(G301), .B(G168), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n840), .B(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(KEYINPUT109), .B1(new_n882), .B2(new_n874), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(new_n876), .B2(new_n882), .ZN(new_n884));
  AOI21_X1  g459(.A(G37), .B1(new_n884), .B2(new_n868), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(new_n868), .B2(new_n884), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT43), .ZN(new_n887));
  XNOR2_X1  g462(.A(KEYINPUT110), .B(KEYINPUT44), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(G397));
  XNOR2_X1  g464(.A(KEYINPUT111), .B(G1384), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n505), .B(KEYINPUT107), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n891), .B1(new_n501), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT112), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT45), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT112), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n896), .B(new_n891), .C1(new_n501), .C2(new_n892), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n894), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  XOR2_X1   g473(.A(KEYINPUT113), .B(G40), .Z(new_n899));
  OR2_X1    g474(.A1(new_n472), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n756), .A2(G2067), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n751), .A2(new_n758), .A3(new_n755), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT115), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n803), .B(G1996), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n907), .B1(new_n901), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n730), .A2(new_n733), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n902), .B1(new_n911), .B2(new_n904), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n902), .A2(G1996), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n913), .B(KEYINPUT46), .Z(new_n914));
  OAI21_X1  g489(.A(new_n901), .B1(new_n803), .B2(new_n905), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XOR2_X1   g491(.A(new_n916), .B(KEYINPUT47), .Z(new_n917));
  AND2_X1   g492(.A1(new_n730), .A2(new_n733), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n901), .B1(new_n918), .B2(new_n910), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n909), .A2(new_n919), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n902), .A2(G1986), .A3(G290), .ZN(new_n921));
  XOR2_X1   g496(.A(new_n921), .B(KEYINPUT48), .Z(new_n922));
  AOI211_X1 g497(.A(new_n912), .B(new_n917), .C1(new_n920), .C2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G1384), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n506), .A2(new_n514), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT50), .ZN(new_n926));
  AOI21_X1  g501(.A(G1384), .B1(new_n855), .B2(new_n512), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT50), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n900), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n924), .B1(new_n501), .B2(new_n892), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n900), .B1(new_n931), .B2(new_n895), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n506), .A2(new_n514), .A3(KEYINPUT45), .A4(new_n924), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI22_X1  g509(.A1(new_n930), .A2(G2084), .B1(new_n934), .B2(G1966), .ZN(new_n935));
  OAI21_X1  g510(.A(G8), .B1(new_n935), .B2(G286), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n936), .A2(KEYINPUT51), .ZN(new_n937));
  INV_X1    g512(.A(new_n900), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(new_n931), .B2(KEYINPUT50), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n939), .B1(KEYINPUT50), .B2(new_n925), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n932), .A2(new_n933), .ZN(new_n941));
  INV_X1    g516(.A(G1966), .ZN(new_n942));
  AOI22_X1  g517(.A1(new_n940), .A2(new_n766), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n943), .A2(G168), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT51), .B1(new_n936), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n937), .A2(new_n945), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n946), .A2(KEYINPUT62), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n946), .A2(KEYINPUT62), .ZN(new_n948));
  NOR2_X1   g523(.A1(G305), .A2(G1981), .ZN(new_n949));
  XNOR2_X1  g524(.A(KEYINPUT117), .B(G86), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n598), .B1(new_n534), .B2(new_n950), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n951), .A2(G1981), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT49), .ZN(new_n953));
  OR3_X1    g528(.A1(new_n949), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G8), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n955), .B1(new_n938), .B2(new_n927), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n953), .B1(new_n952), .B2(new_n949), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n954), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(G1976), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n592), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT116), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n956), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT52), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT52), .B1(G288), .B2(new_n959), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n964), .A2(new_n956), .A3(new_n961), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n958), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(G303), .A2(G8), .ZN(new_n967));
  XOR2_X1   g542(.A(new_n967), .B(KEYINPUT55), .Z(new_n968));
  NOR2_X1   g543(.A1(new_n930), .A2(G2090), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n925), .A2(new_n895), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n890), .B1(new_n855), .B2(new_n512), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n900), .B1(new_n971), .B2(KEYINPUT45), .ZN(new_n972));
  AOI21_X1  g547(.A(G1971), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  OAI211_X1 g548(.A(G8), .B(new_n968), .C1(new_n969), .C2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n973), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n900), .B1(new_n931), .B2(KEYINPUT50), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n506), .A2(new_n514), .A3(new_n928), .A4(new_n924), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OR2_X1    g553(.A1(new_n978), .A2(G2090), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n955), .B1(new_n975), .B2(new_n979), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n966), .B(new_n974), .C1(new_n968), .C2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT122), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n930), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1961), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n926), .A2(KEYINPUT122), .A3(new_n929), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n970), .A2(new_n815), .A3(new_n972), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(G2078), .ZN(new_n989));
  AOI22_X1  g564(.A1(new_n987), .A2(new_n988), .B1(new_n934), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n986), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT125), .B1(new_n991), .B2(G171), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT125), .ZN(new_n993));
  AOI211_X1 g568(.A(new_n993), .B(G301), .C1(new_n986), .C2(new_n990), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NOR4_X1   g570(.A1(new_n947), .A2(new_n948), .A3(new_n981), .A4(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(KEYINPUT118), .B(KEYINPUT63), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n943), .A2(new_n955), .A3(G286), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n997), .B1(new_n981), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT119), .ZN(new_n1001));
  OAI21_X1  g576(.A(G8), .B1(new_n969), .B2(new_n973), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n968), .B1(new_n1002), .B2(KEYINPUT120), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1003), .B1(KEYINPUT120), .B2(new_n1002), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n966), .A2(new_n974), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1004), .A2(KEYINPUT63), .A3(new_n1005), .A4(new_n998), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT119), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1007), .B(new_n997), .C1(new_n981), .C2(new_n999), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1001), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  AOI211_X1 g584(.A(G1976), .B(G288), .C1(new_n954), .C2(new_n957), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1010), .A2(new_n949), .ZN(new_n1011));
  INV_X1    g586(.A(new_n974), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n1011), .A2(new_n956), .B1(new_n1012), .B2(new_n966), .ZN(new_n1013));
  INV_X1    g588(.A(G1348), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n983), .A2(new_n1014), .A3(new_n985), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n938), .A2(new_n927), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1016), .A2(G2067), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1015), .A2(KEYINPUT60), .A3(new_n616), .A4(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1956), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n978), .A2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g596(.A(KEYINPUT56), .B(G2072), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n970), .A2(new_n972), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(G299), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1025), .B1(new_n582), .B2(new_n587), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1024), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1033), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(KEYINPUT61), .A3(new_n1034), .ZN(new_n1035));
  XOR2_X1   g610(.A(KEYINPUT58), .B(G1341), .Z(new_n1036));
  NAND2_X1  g611(.A1(new_n1016), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n970), .A2(new_n972), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1037), .B1(new_n1038), .B2(G1996), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n562), .ZN(new_n1040));
  NOR2_X1   g615(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  XOR2_X1   g617(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n1043));
  NAND3_X1  g618(.A1(new_n1039), .A2(new_n562), .A3(new_n1043), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1019), .A2(new_n1035), .A3(new_n1042), .A4(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT61), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1034), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1033), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1046), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT124), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT124), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1051), .B(new_n1046), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1045), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT60), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1015), .A2(KEYINPUT60), .A3(new_n1018), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(new_n617), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1054), .A2(new_n617), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n1032), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1053), .A2(new_n1058), .B1(new_n1034), .B2(new_n1060), .ZN(new_n1061));
  AOI211_X1 g636(.A(new_n988), .B(G2078), .C1(new_n971), .C2(KEYINPUT45), .ZN(new_n1062));
  NAND2_X1  g637(.A1(G160), .A2(G40), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT45), .B1(new_n893), .B2(KEYINPUT112), .ZN(new_n1064));
  AOI211_X1 g639(.A(KEYINPUT126), .B(new_n1063), .C1(new_n1064), .C2(new_n897), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT126), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1063), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1066), .B1(new_n898), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1062), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n987), .A2(new_n988), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n986), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(G171), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1072), .B(KEYINPUT54), .C1(G171), .C2(new_n991), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n981), .B1(new_n937), .B2(new_n945), .ZN(new_n1074));
  AND4_X1   g649(.A1(G301), .A2(new_n986), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n992), .A2(new_n994), .A3(new_n1075), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1073), .B(new_n1074), .C1(new_n1076), .C2(KEYINPUT54), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1009), .B(new_n1013), .C1(new_n1061), .C2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT127), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1045), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1080), .A2(new_n1081), .A3(new_n1058), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1060), .A2(new_n1034), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n1085));
  INV_X1    g660(.A(new_n995), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1085), .B1(new_n1086), .B2(new_n1075), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1074), .A2(new_n1073), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1084), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT127), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1089), .A2(new_n1090), .A3(new_n1009), .A4(new_n1013), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n996), .B1(new_n1079), .B2(new_n1091), .ZN(new_n1092));
  AND2_X1   g667(.A1(G290), .A2(G1986), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n921), .B1(new_n901), .B2(new_n1093), .ZN(new_n1094));
  XOR2_X1   g669(.A(new_n1094), .B(KEYINPUT114), .Z(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n920), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n923), .B1(new_n1092), .B2(new_n1096), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g672(.A(G319), .ZN(new_n1099));
  NOR3_X1   g673(.A1(G229), .A2(new_n1099), .A3(G227), .ZN(new_n1100));
  NAND4_X1  g674(.A1(new_n887), .A2(new_n666), .A3(new_n864), .A4(new_n1100), .ZN(G225));
  INV_X1    g675(.A(G225), .ZN(G308));
endmodule


