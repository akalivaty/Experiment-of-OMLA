

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579;

  NOR2_X1 U324 ( .A1(n540), .A2(n560), .ZN(n542) );
  XNOR2_X1 U325 ( .A(n511), .B(KEYINPUT48), .ZN(n535) );
  NOR2_X1 U326 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U327 ( .A(KEYINPUT89), .B(n405), .Z(n538) );
  XOR2_X1 U328 ( .A(KEYINPUT3), .B(G162GAT), .Z(n293) );
  XNOR2_X1 U329 ( .A(G155GAT), .B(G141GAT), .ZN(n292) );
  XNOR2_X1 U330 ( .A(n293), .B(n292), .ZN(n294) );
  XNOR2_X1 U331 ( .A(KEYINPUT2), .B(n294), .ZN(n395) );
  XOR2_X1 U332 ( .A(G127GAT), .B(G1GAT), .Z(n329) );
  XOR2_X1 U333 ( .A(G148GAT), .B(G120GAT), .Z(n443) );
  XOR2_X1 U334 ( .A(n329), .B(n443), .Z(n296) );
  XOR2_X1 U335 ( .A(G134GAT), .B(G29GAT), .Z(n320) );
  XOR2_X1 U336 ( .A(KEYINPUT0), .B(G113GAT), .Z(n371) );
  XNOR2_X1 U337 ( .A(n320), .B(n371), .ZN(n295) );
  XNOR2_X1 U338 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U339 ( .A(KEYINPUT4), .B(KEYINPUT88), .Z(n298) );
  NAND2_X1 U340 ( .A1(G225GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U341 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U342 ( .A(n300), .B(n299), .Z(n305) );
  XOR2_X1 U343 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n302) );
  XNOR2_X1 U344 ( .A(G85GAT), .B(G57GAT), .ZN(n301) );
  XNOR2_X1 U345 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U346 ( .A(n303), .B(KEYINPUT5), .ZN(n304) );
  XNOR2_X1 U347 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U348 ( .A(n395), .B(n306), .ZN(n405) );
  XOR2_X1 U349 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n308) );
  XNOR2_X1 U350 ( .A(G50GAT), .B(G43GAT), .ZN(n307) );
  XNOR2_X1 U351 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U352 ( .A(KEYINPUT69), .B(n309), .ZN(n432) );
  XOR2_X1 U353 ( .A(KEYINPUT9), .B(KEYINPUT65), .Z(n311) );
  XNOR2_X1 U354 ( .A(G162GAT), .B(KEYINPUT76), .ZN(n310) );
  XNOR2_X1 U355 ( .A(n311), .B(n310), .ZN(n324) );
  XOR2_X1 U356 ( .A(G92GAT), .B(G106GAT), .Z(n313) );
  XNOR2_X1 U357 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n312) );
  XNOR2_X1 U358 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U359 ( .A(G190GAT), .B(G36GAT), .Z(n344) );
  XOR2_X1 U360 ( .A(n314), .B(n344), .Z(n322) );
  XOR2_X1 U361 ( .A(G85GAT), .B(KEYINPUT74), .Z(n315) );
  XNOR2_X1 U362 ( .A(n315), .B(G99GAT), .ZN(n433) );
  INV_X1 U363 ( .A(n433), .ZN(n316) );
  XOR2_X1 U364 ( .A(n316), .B(KEYINPUT10), .Z(n318) );
  NAND2_X1 U365 ( .A1(G232GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U366 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U367 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U368 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U369 ( .A(n324), .B(n323), .Z(n325) );
  XNOR2_X1 U370 ( .A(n432), .B(n325), .ZN(n506) );
  INV_X1 U371 ( .A(n506), .ZN(n557) );
  XOR2_X1 U372 ( .A(KEYINPUT78), .B(G64GAT), .Z(n327) );
  XNOR2_X1 U373 ( .A(G155GAT), .B(G78GAT), .ZN(n326) );
  XNOR2_X1 U374 ( .A(n327), .B(n326), .ZN(n341) );
  XNOR2_X1 U375 ( .A(G22GAT), .B(G15GAT), .ZN(n328) );
  XNOR2_X1 U376 ( .A(n328), .B(KEYINPUT70), .ZN(n423) );
  XOR2_X1 U377 ( .A(n423), .B(n329), .Z(n331) );
  NAND2_X1 U378 ( .A1(G231GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U379 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U380 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n333) );
  XNOR2_X1 U381 ( .A(KEYINPUT77), .B(KEYINPUT12), .ZN(n332) );
  XNOR2_X1 U382 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U383 ( .A(n335), .B(n334), .Z(n339) );
  XNOR2_X1 U384 ( .A(G211GAT), .B(G183GAT), .ZN(n336) );
  XNOR2_X1 U385 ( .A(n336), .B(G8GAT), .ZN(n343) );
  XNOR2_X1 U386 ( .A(G57GAT), .B(G71GAT), .ZN(n337) );
  XNOR2_X1 U387 ( .A(n337), .B(KEYINPUT13), .ZN(n439) );
  XNOR2_X1 U388 ( .A(n343), .B(n439), .ZN(n338) );
  XNOR2_X1 U389 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U390 ( .A(n341), .B(n340), .ZN(n530) );
  NOR2_X1 U391 ( .A1(n506), .A2(n530), .ZN(n342) );
  XNOR2_X1 U392 ( .A(n342), .B(KEYINPUT16), .ZN(n413) );
  XOR2_X1 U393 ( .A(KEYINPUT91), .B(G204GAT), .Z(n346) );
  XNOR2_X1 U394 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U395 ( .A(n346), .B(n345), .ZN(n351) );
  XNOR2_X1 U396 ( .A(G92GAT), .B(G64GAT), .ZN(n347) );
  XNOR2_X1 U397 ( .A(n347), .B(G176GAT), .ZN(n438) );
  XOR2_X1 U398 ( .A(KEYINPUT90), .B(n438), .Z(n349) );
  NAND2_X1 U399 ( .A1(G226GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U400 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U401 ( .A(n351), .B(n350), .Z(n359) );
  XOR2_X1 U402 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n353) );
  XNOR2_X1 U403 ( .A(KEYINPUT18), .B(G169GAT), .ZN(n352) );
  XNOR2_X1 U404 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U405 ( .A(KEYINPUT81), .B(n354), .Z(n379) );
  XOR2_X1 U406 ( .A(KEYINPUT86), .B(G197GAT), .Z(n356) );
  XNOR2_X1 U407 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n355) );
  XNOR2_X1 U408 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U409 ( .A(KEYINPUT85), .B(n357), .Z(n392) );
  XNOR2_X1 U410 ( .A(n379), .B(n392), .ZN(n358) );
  XNOR2_X1 U411 ( .A(n359), .B(n358), .ZN(n536) );
  XOR2_X1 U412 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n361) );
  XNOR2_X1 U413 ( .A(G71GAT), .B(G15GAT), .ZN(n360) );
  XNOR2_X1 U414 ( .A(n361), .B(n360), .ZN(n365) );
  XOR2_X1 U415 ( .A(KEYINPUT64), .B(KEYINPUT79), .Z(n363) );
  XNOR2_X1 U416 ( .A(G183GAT), .B(KEYINPUT20), .ZN(n362) );
  XNOR2_X1 U417 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U418 ( .A(n365), .B(n364), .Z(n377) );
  XOR2_X1 U419 ( .A(G176GAT), .B(KEYINPUT80), .Z(n367) );
  XNOR2_X1 U420 ( .A(G120GAT), .B(G127GAT), .ZN(n366) );
  XNOR2_X1 U421 ( .A(n367), .B(n366), .ZN(n375) );
  XOR2_X1 U422 ( .A(G190GAT), .B(G99GAT), .Z(n369) );
  XNOR2_X1 U423 ( .A(G134GAT), .B(G43GAT), .ZN(n368) );
  XNOR2_X1 U424 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U425 ( .A(n371), .B(n370), .Z(n373) );
  NAND2_X1 U426 ( .A1(G227GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U427 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U428 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U429 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U430 ( .A(n379), .B(n378), .ZN(n500) );
  NOR2_X1 U431 ( .A1(n536), .A2(n500), .ZN(n380) );
  XNOR2_X1 U432 ( .A(KEYINPUT95), .B(n380), .ZN(n397) );
  XOR2_X1 U433 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n382) );
  XNOR2_X1 U434 ( .A(G50GAT), .B(G22GAT), .ZN(n381) );
  XNOR2_X1 U435 ( .A(n382), .B(n381), .ZN(n386) );
  XOR2_X1 U436 ( .A(KEYINPUT24), .B(KEYINPUT87), .Z(n384) );
  XNOR2_X1 U437 ( .A(G148GAT), .B(KEYINPUT84), .ZN(n383) );
  XNOR2_X1 U438 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U439 ( .A(n386), .B(n385), .Z(n394) );
  XOR2_X1 U440 ( .A(KEYINPUT73), .B(G204GAT), .Z(n388) );
  XNOR2_X1 U441 ( .A(G106GAT), .B(G78GAT), .ZN(n387) );
  XNOR2_X1 U442 ( .A(n388), .B(n387), .ZN(n434) );
  XOR2_X1 U443 ( .A(G211GAT), .B(n434), .Z(n390) );
  NAND2_X1 U444 ( .A1(G228GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U445 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U446 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U447 ( .A(n394), .B(n393), .ZN(n396) );
  XOR2_X1 U448 ( .A(n396), .B(n395), .Z(n540) );
  INV_X1 U449 ( .A(n540), .ZN(n409) );
  NAND2_X1 U450 ( .A1(n397), .A2(n409), .ZN(n398) );
  XNOR2_X1 U451 ( .A(n398), .B(KEYINPUT96), .ZN(n399) );
  XNOR2_X1 U452 ( .A(n399), .B(KEYINPUT25), .ZN(n403) );
  XNOR2_X1 U453 ( .A(n536), .B(KEYINPUT27), .ZN(n407) );
  NAND2_X1 U454 ( .A1(n540), .A2(n500), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n400), .B(KEYINPUT94), .ZN(n401) );
  XNOR2_X1 U456 ( .A(KEYINPUT26), .B(n401), .ZN(n561) );
  NOR2_X1 U457 ( .A1(n407), .A2(n561), .ZN(n402) );
  NOR2_X1 U458 ( .A1(n403), .A2(n402), .ZN(n404) );
  XNOR2_X1 U459 ( .A(n404), .B(KEYINPUT97), .ZN(n406) );
  NAND2_X1 U460 ( .A1(n406), .A2(n405), .ZN(n412) );
  NOR2_X1 U461 ( .A1(n407), .A2(n538), .ZN(n408) );
  XNOR2_X1 U462 ( .A(n408), .B(KEYINPUT92), .ZN(n523) );
  XNOR2_X1 U463 ( .A(n409), .B(KEYINPUT28), .ZN(n496) );
  NAND2_X1 U464 ( .A1(n523), .A2(n496), .ZN(n512) );
  XNOR2_X1 U465 ( .A(KEYINPUT93), .B(n512), .ZN(n410) );
  NAND2_X1 U466 ( .A1(n410), .A2(n500), .ZN(n411) );
  NAND2_X1 U467 ( .A1(n412), .A2(n411), .ZN(n458) );
  NAND2_X1 U468 ( .A1(n413), .A2(n458), .ZN(n414) );
  XOR2_X1 U469 ( .A(KEYINPUT98), .B(n414), .Z(n478) );
  XOR2_X1 U470 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n416) );
  XNOR2_X1 U471 ( .A(KEYINPUT68), .B(KEYINPUT66), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n430) );
  XOR2_X1 U473 ( .A(G197GAT), .B(G169GAT), .Z(n418) );
  XNOR2_X1 U474 ( .A(G141GAT), .B(G113GAT), .ZN(n417) );
  XNOR2_X1 U475 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U476 ( .A(KEYINPUT71), .B(KEYINPUT29), .Z(n420) );
  XNOR2_X1 U477 ( .A(G1GAT), .B(G8GAT), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U479 ( .A(n422), .B(n421), .Z(n428) );
  XOR2_X1 U480 ( .A(n423), .B(G36GAT), .Z(n425) );
  NAND2_X1 U481 ( .A1(G229GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U483 ( .A(G29GAT), .B(n426), .ZN(n427) );
  XNOR2_X1 U484 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U485 ( .A(n430), .B(n429), .Z(n431) );
  XNOR2_X1 U486 ( .A(n432), .B(n431), .ZN(n545) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n447) );
  XOR2_X1 U488 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n436) );
  NAND2_X1 U489 ( .A1(G230GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U491 ( .A(n437), .B(KEYINPUT32), .Z(n441) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U494 ( .A(n442), .B(KEYINPUT75), .Z(n445) );
  XNOR2_X1 U495 ( .A(n443), .B(KEYINPUT72), .ZN(n444) );
  XNOR2_X1 U496 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U497 ( .A(n447), .B(n446), .ZN(n568) );
  NOR2_X1 U498 ( .A1(n545), .A2(n568), .ZN(n463) );
  NAND2_X1 U499 ( .A1(n478), .A2(n463), .ZN(n448) );
  XOR2_X1 U500 ( .A(KEYINPUT99), .B(n448), .Z(n455) );
  NOR2_X1 U501 ( .A1(n538), .A2(n455), .ZN(n450) );
  XNOR2_X1 U502 ( .A(KEYINPUT100), .B(KEYINPUT34), .ZN(n449) );
  XNOR2_X1 U503 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U504 ( .A(G1GAT), .B(n451), .Z(G1324GAT) );
  NOR2_X1 U505 ( .A1(n536), .A2(n455), .ZN(n452) );
  XOR2_X1 U506 ( .A(G8GAT), .B(n452), .Z(G1325GAT) );
  NOR2_X1 U507 ( .A1(n500), .A2(n455), .ZN(n454) );
  XNOR2_X1 U508 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n453) );
  XNOR2_X1 U509 ( .A(n454), .B(n453), .ZN(G1326GAT) );
  NOR2_X1 U510 ( .A1(n496), .A2(n455), .ZN(n457) );
  XNOR2_X1 U511 ( .A(G22GAT), .B(KEYINPUT101), .ZN(n456) );
  XNOR2_X1 U512 ( .A(n457), .B(n456), .ZN(G1327GAT) );
  XNOR2_X1 U513 ( .A(KEYINPUT37), .B(KEYINPUT104), .ZN(n462) );
  NAND2_X1 U514 ( .A1(n530), .A2(n458), .ZN(n459) );
  XNOR2_X1 U515 ( .A(n459), .B(KEYINPUT103), .ZN(n460) );
  XNOR2_X1 U516 ( .A(n506), .B(KEYINPUT36), .ZN(n575) );
  NAND2_X1 U517 ( .A1(n460), .A2(n575), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n462), .B(n461), .ZN(n487) );
  NAND2_X1 U519 ( .A1(n487), .A2(n463), .ZN(n464) );
  XNOR2_X1 U520 ( .A(n464), .B(KEYINPUT38), .ZN(n475) );
  NOR2_X1 U521 ( .A1(n475), .A2(n538), .ZN(n468) );
  XOR2_X1 U522 ( .A(KEYINPUT102), .B(KEYINPUT39), .Z(n466) );
  XNOR2_X1 U523 ( .A(G29GAT), .B(KEYINPUT105), .ZN(n465) );
  XNOR2_X1 U524 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U525 ( .A(n468), .B(n467), .ZN(G1328GAT) );
  XNOR2_X1 U526 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n470) );
  NOR2_X1 U527 ( .A1(n536), .A2(n475), .ZN(n469) );
  XNOR2_X1 U528 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U529 ( .A(G36GAT), .B(n471), .ZN(G1329GAT) );
  NOR2_X1 U530 ( .A1(n475), .A2(n500), .ZN(n473) );
  XNOR2_X1 U531 ( .A(KEYINPUT40), .B(KEYINPUT108), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U533 ( .A(G43GAT), .B(n474), .Z(G1330GAT) );
  NOR2_X1 U534 ( .A1(n475), .A2(n496), .ZN(n477) );
  XNOR2_X1 U535 ( .A(G50GAT), .B(KEYINPUT109), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n477), .B(n476), .ZN(G1331GAT) );
  XNOR2_X1 U537 ( .A(KEYINPUT41), .B(n568), .ZN(n549) );
  INV_X1 U538 ( .A(n545), .ZN(n562) );
  NOR2_X1 U539 ( .A1(n549), .A2(n562), .ZN(n488) );
  NAND2_X1 U540 ( .A1(n488), .A2(n478), .ZN(n483) );
  NOR2_X1 U541 ( .A1(n538), .A2(n483), .ZN(n479) );
  XOR2_X1 U542 ( .A(G57GAT), .B(n479), .Z(n480) );
  XNOR2_X1 U543 ( .A(KEYINPUT42), .B(n480), .ZN(G1332GAT) );
  NOR2_X1 U544 ( .A1(n536), .A2(n483), .ZN(n481) );
  XOR2_X1 U545 ( .A(G64GAT), .B(n481), .Z(G1333GAT) );
  NOR2_X1 U546 ( .A1(n500), .A2(n483), .ZN(n482) );
  XOR2_X1 U547 ( .A(G71GAT), .B(n482), .Z(G1334GAT) );
  NOR2_X1 U548 ( .A1(n496), .A2(n483), .ZN(n485) );
  XNOR2_X1 U549 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n484) );
  XNOR2_X1 U550 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U551 ( .A(G78GAT), .B(n486), .ZN(G1335GAT) );
  NAND2_X1 U552 ( .A1(n488), .A2(n487), .ZN(n495) );
  NOR2_X1 U553 ( .A1(n538), .A2(n495), .ZN(n490) );
  XNOR2_X1 U554 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n489) );
  XNOR2_X1 U555 ( .A(n490), .B(n489), .ZN(G1336GAT) );
  NOR2_X1 U556 ( .A1(n536), .A2(n495), .ZN(n491) );
  XOR2_X1 U557 ( .A(KEYINPUT112), .B(n491), .Z(n492) );
  XNOR2_X1 U558 ( .A(G92GAT), .B(n492), .ZN(G1337GAT) );
  NOR2_X1 U559 ( .A1(n500), .A2(n495), .ZN(n494) );
  XNOR2_X1 U560 ( .A(G99GAT), .B(KEYINPUT113), .ZN(n493) );
  XNOR2_X1 U561 ( .A(n494), .B(n493), .ZN(G1338GAT) );
  NOR2_X1 U562 ( .A1(n496), .A2(n495), .ZN(n498) );
  XNOR2_X1 U563 ( .A(KEYINPUT114), .B(KEYINPUT44), .ZN(n497) );
  XNOR2_X1 U564 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U565 ( .A(G106GAT), .B(n499), .Z(G1339GAT) );
  INV_X1 U566 ( .A(n500), .ZN(n544) );
  INV_X1 U567 ( .A(n530), .ZN(n573) );
  NAND2_X1 U568 ( .A1(n575), .A2(n573), .ZN(n501) );
  XOR2_X1 U569 ( .A(KEYINPUT45), .B(n501), .Z(n502) );
  NAND2_X1 U570 ( .A1(n545), .A2(n502), .ZN(n503) );
  NOR2_X1 U571 ( .A1(n568), .A2(n503), .ZN(n510) );
  NOR2_X1 U572 ( .A1(n545), .A2(n549), .ZN(n504) );
  XNOR2_X1 U573 ( .A(n504), .B(KEYINPUT46), .ZN(n505) );
  NOR2_X1 U574 ( .A1(n506), .A2(n505), .ZN(n507) );
  XOR2_X1 U575 ( .A(KEYINPUT115), .B(n530), .Z(n552) );
  NAND2_X1 U576 ( .A1(n507), .A2(n552), .ZN(n508) );
  XNOR2_X1 U577 ( .A(n508), .B(KEYINPUT47), .ZN(n509) );
  NOR2_X1 U578 ( .A1(n510), .A2(n509), .ZN(n511) );
  NOR2_X1 U579 ( .A1(n512), .A2(n535), .ZN(n513) );
  NAND2_X1 U580 ( .A1(n544), .A2(n513), .ZN(n520) );
  NOR2_X1 U581 ( .A1(n545), .A2(n520), .ZN(n514) );
  XOR2_X1 U582 ( .A(G113GAT), .B(n514), .Z(G1340GAT) );
  NOR2_X1 U583 ( .A1(n549), .A2(n520), .ZN(n516) );
  XNOR2_X1 U584 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n515) );
  XNOR2_X1 U585 ( .A(n516), .B(n515), .ZN(G1341GAT) );
  NOR2_X1 U586 ( .A1(n552), .A2(n520), .ZN(n518) );
  XNOR2_X1 U587 ( .A(KEYINPUT50), .B(KEYINPUT116), .ZN(n517) );
  XNOR2_X1 U588 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U589 ( .A(G127GAT), .B(n519), .Z(G1342GAT) );
  NOR2_X1 U590 ( .A1(n557), .A2(n520), .ZN(n522) );
  XNOR2_X1 U591 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n521) );
  XNOR2_X1 U592 ( .A(n522), .B(n521), .ZN(G1343GAT) );
  NOR2_X1 U593 ( .A1(n561), .A2(n535), .ZN(n524) );
  NAND2_X1 U594 ( .A1(n524), .A2(n523), .ZN(n533) );
  NOR2_X1 U595 ( .A1(n545), .A2(n533), .ZN(n526) );
  XNOR2_X1 U596 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n525) );
  XNOR2_X1 U597 ( .A(n526), .B(n525), .ZN(G1344GAT) );
  NOR2_X1 U598 ( .A1(n549), .A2(n533), .ZN(n528) );
  XNOR2_X1 U599 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n527) );
  XNOR2_X1 U600 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U601 ( .A(G148GAT), .B(n529), .ZN(G1345GAT) );
  NOR2_X1 U602 ( .A1(n530), .A2(n533), .ZN(n531) );
  XOR2_X1 U603 ( .A(KEYINPUT118), .B(n531), .Z(n532) );
  XNOR2_X1 U604 ( .A(G155GAT), .B(n532), .ZN(G1346GAT) );
  NOR2_X1 U605 ( .A1(n557), .A2(n533), .ZN(n534) );
  XOR2_X1 U606 ( .A(G162GAT), .B(n534), .Z(G1347GAT) );
  NOR2_X1 U607 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U608 ( .A(n537), .B(KEYINPUT54), .ZN(n539) );
  NAND2_X1 U609 ( .A1(n539), .A2(n538), .ZN(n560) );
  XNOR2_X1 U610 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n541) );
  XNOR2_X1 U611 ( .A(n542), .B(n541), .ZN(n543) );
  NAND2_X1 U612 ( .A1(n544), .A2(n543), .ZN(n556) );
  NOR2_X1 U613 ( .A1(n545), .A2(n556), .ZN(n546) );
  XOR2_X1 U614 ( .A(G169GAT), .B(n546), .Z(G1348GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n548) );
  XNOR2_X1 U616 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n547) );
  XNOR2_X1 U617 ( .A(n548), .B(n547), .ZN(n551) );
  NOR2_X1 U618 ( .A1(n549), .A2(n556), .ZN(n550) );
  XOR2_X1 U619 ( .A(n551), .B(n550), .Z(G1349GAT) );
  NOR2_X1 U620 ( .A1(n552), .A2(n556), .ZN(n554) );
  XNOR2_X1 U621 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U623 ( .A(G183GAT), .B(n555), .ZN(G1350GAT) );
  XOR2_X1 U624 ( .A(G190GAT), .B(n558), .Z(n559) );
  XNOR2_X1 U625 ( .A(KEYINPUT58), .B(n559), .ZN(G1351GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n564) );
  NOR2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n576) );
  NAND2_X1 U628 ( .A1(n576), .A2(n562), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(n565) );
  XOR2_X1 U630 ( .A(n565), .B(KEYINPUT59), .Z(n567) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1352GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n570) );
  NAND2_X1 U634 ( .A1(n576), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n572) );
  XOR2_X1 U636 ( .A(G204GAT), .B(KEYINPUT125), .Z(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1353GAT) );
  NAND2_X1 U638 ( .A1(n576), .A2(n573), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n578) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n579), .ZN(G1355GAT) );
endmodule

