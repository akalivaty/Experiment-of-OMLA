//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n812, new_n813, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939;
  XNOR2_X1  g000(.A(G120gat), .B(G148gat), .ZN(new_n202));
  INV_X1    g001(.A(G176gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G204gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT104), .ZN(new_n208));
  NAND2_X1  g007(.A1(G71gat), .A2(G78gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT9), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT94), .ZN(new_n212));
  INV_X1    g011(.A(G64gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G57gat), .ZN(new_n214));
  INV_X1    g013(.A(G57gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G64gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT94), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n209), .A2(new_n218), .A3(new_n210), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n212), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G71gat), .B(G78gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n212), .A2(new_n217), .A3(new_n221), .A4(new_n219), .ZN(new_n224));
  INV_X1    g023(.A(G85gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT99), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT99), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G85gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G92gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(G85gat), .A2(G92gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT7), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT7), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n233), .A2(G85gat), .A3(G92gat), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n229), .A2(new_n230), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G99gat), .A2(G106gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT98), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT98), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(G99gat), .A3(G106gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n237), .A2(new_n239), .A3(KEYINPUT8), .ZN(new_n240));
  INV_X1    g039(.A(G99gat), .ZN(new_n241));
  INV_X1    g040(.A(G106gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(new_n236), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT102), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n243), .A2(KEYINPUT102), .A3(new_n236), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n235), .A2(new_n240), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n223), .B(new_n224), .C1(new_n248), .C2(KEYINPUT103), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT103), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n227), .A2(G85gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n225), .A2(KEYINPUT99), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n230), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n232), .A2(new_n234), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n240), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n246), .A2(new_n247), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n235), .A2(new_n244), .A3(new_n240), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n250), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n208), .B1(new_n249), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n223), .A2(new_n224), .ZN(new_n261));
  INV_X1    g060(.A(new_n244), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n255), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  AND4_X1   g063(.A1(new_n244), .A2(new_n253), .A3(new_n240), .A4(new_n254), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n261), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT103), .B1(new_n255), .B2(new_n256), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n267), .A2(new_n261), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT103), .B1(new_n248), .B2(new_n265), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(new_n269), .A3(KEYINPUT104), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n260), .A2(new_n266), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT105), .ZN(new_n272));
  NAND2_X1  g071(.A1(G230gat), .A2(G233gat), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n271), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT10), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n260), .A2(new_n276), .A3(new_n270), .A4(new_n266), .ZN(new_n277));
  INV_X1    g076(.A(new_n261), .ZN(new_n278));
  AND3_X1   g077(.A1(new_n263), .A2(KEYINPUT100), .A3(new_n258), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT100), .B1(new_n263), .B2(new_n258), .ZN(new_n280));
  OAI211_X1 g079(.A(KEYINPUT10), .B(new_n278), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n274), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n275), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n272), .B1(new_n271), .B2(new_n274), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n207), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NOR4_X1   g085(.A1(new_n275), .A2(new_n282), .A3(new_n284), .A4(new_n206), .ZN(new_n287));
  OR2_X1    g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n289));
  XNOR2_X1  g088(.A(G15gat), .B(G22gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT16), .ZN(new_n291));
  OR2_X1    g090(.A1(new_n291), .A2(G1gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(G1gat), .B2(new_n290), .ZN(new_n294));
  XOR2_X1   g093(.A(new_n294), .B(G8gat), .Z(new_n295));
  NAND2_X1  g094(.A1(new_n278), .A2(KEYINPUT21), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT96), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT97), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n297), .B1(new_n295), .B2(new_n296), .ZN(new_n301));
  NOR3_X1   g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n295), .A2(new_n296), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT96), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT97), .B1(new_n304), .B2(new_n298), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n289), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n278), .A2(KEYINPUT21), .ZN(new_n307));
  NAND2_X1  g106(.A1(G231gat), .A2(G233gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n308), .B(KEYINPUT95), .ZN(new_n309));
  XNOR2_X1  g108(.A(G183gat), .B(G211gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n307), .B(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G127gat), .B(G155gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n312), .B(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n300), .B1(new_n299), .B2(new_n301), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n304), .A2(KEYINPUT97), .A3(new_n298), .ZN(new_n316));
  INV_X1    g115(.A(new_n289), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  AND3_X1   g117(.A1(new_n306), .A2(new_n314), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n314), .B1(new_n306), .B2(new_n318), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(G190gat), .B(G218gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n279), .A2(new_n280), .ZN(new_n324));
  INV_X1    g123(.A(G29gat), .ZN(new_n325));
  INV_X1    g124(.A(G36gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n326), .A3(KEYINPUT89), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT89), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n328), .B1(G29gat), .B2(G36gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n329), .A3(KEYINPUT14), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT14), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n328), .B(new_n331), .C1(G29gat), .C2(G36gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(G29gat), .A2(G36gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT15), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n330), .A2(KEYINPUT15), .A3(new_n332), .A4(new_n333), .ZN(new_n337));
  XNOR2_X1  g136(.A(G43gat), .B(G50gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n330), .A2(new_n333), .ZN(new_n340));
  INV_X1    g139(.A(new_n338), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n340), .A2(KEYINPUT15), .A3(new_n332), .A4(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT17), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n339), .A2(KEYINPUT17), .A3(new_n342), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n324), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n343), .B1(new_n279), .B2(new_n280), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(G134gat), .ZN(new_n351));
  INV_X1    g150(.A(G134gat), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n347), .A2(new_n352), .A3(new_n348), .A4(new_n349), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n323), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n356), .B(G162gat), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n351), .A2(new_n353), .A3(new_n323), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n355), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n357), .ZN(new_n360));
  INV_X1    g159(.A(new_n358), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n360), .B1(new_n361), .B2(new_n354), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n321), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT101), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n321), .A2(KEYINPUT101), .A3(new_n362), .A4(new_n359), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT85), .ZN(new_n368));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n369), .B(KEYINPUT80), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G127gat), .B(G134gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT71), .ZN(new_n373));
  INV_X1    g172(.A(G113gat), .ZN(new_n374));
  INV_X1    g173(.A(G120gat), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT1), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n376), .B1(new_n374), .B2(new_n375), .ZN(new_n377));
  INV_X1    g176(.A(G127gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(G134gat), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n373), .B(new_n377), .C1(KEYINPUT71), .C2(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(KEYINPUT72), .B(G120gat), .Z(new_n381));
  OAI211_X1 g180(.A(new_n372), .B(new_n376), .C1(new_n381), .C2(new_n374), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  XOR2_X1   g182(.A(G141gat), .B(G148gat), .Z(new_n384));
  INV_X1    g183(.A(G155gat), .ZN(new_n385));
  INV_X1    g184(.A(G162gat), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT2), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G155gat), .B(G162gat), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n384), .A2(new_n389), .A3(new_n387), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n383), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n380), .A2(new_n391), .A3(new_n392), .A4(new_n382), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n371), .B1(new_n396), .B2(KEYINPUT5), .ZN(new_n397));
  OR3_X1    g196(.A1(new_n395), .A2(KEYINPUT83), .A3(KEYINPUT4), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n395), .A2(KEYINPUT4), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT84), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT84), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n395), .A2(new_n401), .A3(KEYINPUT4), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT83), .B1(new_n395), .B2(KEYINPUT4), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n398), .A2(new_n400), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  OR2_X1    g203(.A1(new_n393), .A2(KEYINPUT3), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n393), .A2(KEYINPUT3), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(new_n406), .A3(new_n383), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT5), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n397), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n395), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(KEYINPUT81), .A3(new_n412), .ZN(new_n413));
  AND2_X1   g212(.A1(new_n407), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n411), .A2(new_n412), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT81), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(new_n416), .A3(new_n399), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n414), .A2(KEYINPUT5), .A3(new_n417), .A4(new_n371), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n410), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n420));
  XNOR2_X1  g219(.A(G1gat), .B(G29gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G57gat), .B(G85gat), .ZN(new_n423));
  XOR2_X1   g222(.A(new_n422), .B(new_n423), .Z(new_n424));
  NAND2_X1  g223(.A1(new_n419), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT6), .ZN(new_n426));
  INV_X1    g225(.A(new_n424), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n410), .A2(new_n427), .A3(new_n418), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n425), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n428), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT6), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n368), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT85), .B1(new_n430), .B2(KEYINPUT6), .ZN(new_n433));
  XNOR2_X1  g232(.A(G211gat), .B(G218gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(KEYINPUT76), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT75), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n436), .A2(KEYINPUT22), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(KEYINPUT22), .ZN(new_n438));
  NAND2_X1  g237(.A1(G211gat), .A2(G218gat), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G197gat), .B(G204gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  XOR2_X1   g241(.A(new_n435), .B(new_n442), .Z(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(G183gat), .A2(G190gat), .ZN(new_n445));
  OR2_X1    g244(.A1(new_n445), .A2(KEYINPUT66), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT24), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(KEYINPUT66), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n445), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT24), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT67), .ZN(new_n452));
  OR2_X1    g251(.A1(G183gat), .A2(G190gat), .ZN(new_n453));
  OR3_X1    g252(.A1(new_n445), .A2(new_n447), .A3(KEYINPUT67), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n449), .A2(new_n452), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(G169gat), .A2(G176gat), .ZN(new_n456));
  OR3_X1    g255(.A1(new_n456), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n457));
  NAND2_X1  g256(.A1(G169gat), .A2(G176gat), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT64), .B1(new_n456), .B2(KEYINPUT23), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT23), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n456), .B(KEYINPUT65), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n455), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT25), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT26), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n458), .B1(new_n456), .B2(new_n465), .ZN(new_n466));
  OR2_X1    g265(.A1(new_n466), .A2(KEYINPUT70), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(KEYINPUT70), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n467), .B(new_n468), .C1(KEYINPUT26), .C2(new_n462), .ZN(new_n469));
  XNOR2_X1  g268(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n470));
  XOR2_X1   g269(.A(KEYINPUT27), .B(G183gat), .Z(new_n471));
  INV_X1    g270(.A(KEYINPUT68), .ZN(new_n472));
  AOI21_X1  g271(.A(G190gat), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT27), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT68), .B1(new_n474), .B2(G183gat), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n470), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT28), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n471), .A2(new_n477), .A3(G190gat), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n469), .B(new_n445), .C1(new_n476), .C2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n453), .A2(KEYINPUT24), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n445), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT25), .B1(new_n481), .B2(new_n451), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n456), .A2(KEYINPUT23), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n460), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n464), .A2(new_n479), .A3(new_n484), .ZN(new_n485));
  AND2_X1   g284(.A1(G226gat), .A2(G233gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT29), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n444), .B(new_n487), .C1(new_n489), .C2(new_n486), .ZN(new_n490));
  INV_X1    g289(.A(new_n487), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n486), .B1(new_n485), .B2(new_n488), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n443), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(G8gat), .B(G36gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n494), .B(new_n213), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(new_n230), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n490), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n498), .B(KEYINPUT78), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n432), .A2(new_n433), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT37), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n490), .A2(new_n493), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n496), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n501), .B1(new_n490), .B2(new_n493), .ZN(new_n504));
  OR3_X1    g303(.A1(new_n503), .A2(KEYINPUT38), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT77), .ZN(new_n506));
  INV_X1    g305(.A(new_n490), .ZN(new_n507));
  INV_X1    g306(.A(new_n493), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n490), .A2(new_n493), .A3(KEYINPUT77), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n501), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT38), .B1(new_n511), .B2(new_n503), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT86), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g313(.A(KEYINPUT86), .B(KEYINPUT38), .C1(new_n511), .C2(new_n503), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n500), .A2(new_n505), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(KEYINPUT31), .B(G50gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n443), .A2(KEYINPUT29), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n393), .B1(new_n518), .B2(KEYINPUT3), .ZN(new_n519));
  INV_X1    g318(.A(G78gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n405), .A2(new_n488), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n443), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n520), .B1(new_n519), .B2(new_n522), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n517), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n519), .A2(new_n522), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(G78gat), .ZN(new_n527));
  INV_X1    g326(.A(new_n517), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(G228gat), .A2(G233gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(G22gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(new_n242), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n525), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n533), .B1(new_n525), .B2(new_n530), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n371), .B1(new_n404), .B2(new_n407), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT39), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n396), .A2(new_n371), .ZN(new_n540));
  OR3_X1    g339(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n427), .B1(new_n538), .B2(new_n539), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(KEYINPUT40), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n428), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT79), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(new_n498), .B2(KEYINPUT78), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT30), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n498), .A2(new_n545), .A3(KEYINPUT30), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n498), .A2(KEYINPUT78), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n509), .A2(new_n510), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n496), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n544), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n541), .A2(new_n542), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n555), .A2(KEYINPUT40), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n537), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n485), .A2(new_n380), .A3(new_n382), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n464), .A2(new_n479), .A3(new_n383), .A4(new_n484), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n558), .A2(G227gat), .A3(G233gat), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT32), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT33), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G15gat), .B(G43gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(G71gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(new_n241), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n561), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n566), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n560), .B(KEYINPUT32), .C1(new_n562), .C2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n558), .A2(new_n559), .ZN(new_n571));
  NAND2_X1  g370(.A1(G227gat), .A2(G233gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT34), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT74), .ZN(new_n576));
  INV_X1    g375(.A(new_n574), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n577), .A2(new_n569), .A3(new_n567), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT74), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n570), .A2(new_n579), .A3(new_n574), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n576), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT36), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT73), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n577), .A2(new_n584), .A3(new_n570), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n577), .B1(new_n584), .B2(new_n570), .ZN(new_n586));
  OAI21_X1  g385(.A(KEYINPUT36), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g386(.A1(new_n516), .A2(new_n557), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n546), .A2(new_n547), .B1(KEYINPUT78), .B2(new_n498), .ZN(new_n589));
  AOI22_X1  g388(.A1(new_n589), .A2(new_n549), .B1(new_n552), .B2(new_n496), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n429), .A2(new_n431), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(new_n537), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT87), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n432), .A2(new_n433), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n551), .A2(new_n553), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n590), .B(KEYINPUT87), .C1(new_n432), .C2(new_n433), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n536), .A2(new_n576), .A3(new_n578), .A4(new_n580), .ZN(new_n599));
  NOR2_X1   g398(.A1(KEYINPUT88), .A2(KEYINPUT35), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(KEYINPUT88), .A2(KEYINPUT35), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n597), .A2(new_n598), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n536), .B1(new_n585), .B2(new_n586), .ZN(new_n604));
  OAI21_X1  g403(.A(KEYINPUT35), .B1(new_n592), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g404(.A1(new_n588), .A2(new_n593), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT18), .ZN(new_n607));
  AOI22_X1  g406(.A1(new_n607), .A2(KEYINPUT91), .B1(G229gat), .B2(G233gat), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n345), .A2(KEYINPUT90), .A3(new_n295), .A4(new_n346), .ZN(new_n609));
  AND3_X1   g408(.A1(new_n339), .A2(KEYINPUT17), .A3(new_n342), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT17), .B1(new_n339), .B2(new_n342), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n294), .B(G8gat), .ZN(new_n612));
  NOR3_X1   g411(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT90), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n614), .B1(new_n343), .B2(new_n612), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n608), .B(new_n609), .C1(new_n613), .C2(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n607), .A2(KEYINPUT91), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n295), .A2(new_n342), .A3(new_n339), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n343), .A2(new_n612), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n620), .A2(KEYINPUT92), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT92), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n343), .A2(new_n623), .A3(new_n612), .ZN(new_n624));
  NAND2_X1  g423(.A1(G229gat), .A2(G233gat), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n625), .B(KEYINPUT13), .Z(new_n626));
  NAND3_X1  g425(.A1(new_n622), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n345), .A2(new_n295), .A3(new_n346), .ZN(new_n628));
  INV_X1    g427(.A(new_n615), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n630), .A2(new_n617), .A3(new_n608), .A4(new_n609), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n619), .A2(new_n627), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G113gat), .B(G141gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G197gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT11), .ZN(new_n635));
  INV_X1    g434(.A(G169gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT12), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n632), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n619), .A2(new_n638), .A3(new_n627), .A4(new_n631), .ZN(new_n641));
  AND2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(KEYINPUT93), .B1(new_n606), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n603), .A2(new_n605), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n516), .A2(new_n557), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n583), .A2(new_n587), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(new_n593), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT93), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n640), .A2(new_n641), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  AOI211_X1 g450(.A(new_n288), .B(new_n367), .C1(new_n643), .C2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n591), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT106), .B(G1gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(G1324gat));
  XOR2_X1   g455(.A(KEYINPUT42), .B(G8gat), .Z(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n652), .A2(new_n596), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n658), .B1(new_n659), .B2(new_n291), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n652), .A2(KEYINPUT16), .A3(new_n596), .A4(new_n657), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n660), .A2(new_n661), .A3(new_n663), .ZN(G1325gat));
  INV_X1    g463(.A(new_n581), .ZN(new_n665));
  AOI21_X1  g464(.A(G15gat), .B1(new_n652), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n646), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(G15gat), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n666), .B1(new_n652), .B2(new_n669), .ZN(G1326gat));
  NAND2_X1  g469(.A1(new_n652), .A2(new_n537), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT43), .B(G22gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1327gat));
  NOR2_X1   g472(.A1(new_n288), .A2(new_n321), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n675), .B1(new_n643), .B2(new_n651), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n362), .A2(new_n359), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n676), .A2(new_n325), .A3(new_n653), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT45), .ZN(new_n679));
  INV_X1    g478(.A(new_n677), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n680), .B1(new_n644), .B2(new_n647), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT44), .B1(new_n606), .B2(new_n680), .ZN(new_n684));
  AOI211_X1 g483(.A(new_n642), .B(new_n675), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n685), .A2(KEYINPUT107), .A3(new_n653), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT107), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n681), .A2(new_n682), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n606), .A2(KEYINPUT44), .A3(new_n680), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n650), .B(new_n674), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n687), .B1(new_n690), .B2(new_n591), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n686), .A2(new_n691), .A3(G29gat), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n679), .A2(new_n692), .ZN(G1328gat));
  AND2_X1   g492(.A1(new_n676), .A2(new_n677), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n694), .A2(new_n326), .A3(new_n596), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT46), .ZN(new_n696));
  OAI21_X1  g495(.A(G36gat), .B1(new_n690), .B2(new_n590), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n694), .A2(new_n698), .A3(new_n326), .A4(new_n596), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n696), .A2(new_n697), .A3(new_n699), .ZN(G1329gat));
  OAI21_X1  g499(.A(G43gat), .B1(new_n690), .B2(new_n646), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n581), .A2(G43gat), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n676), .A2(new_n677), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT47), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n701), .B(new_n703), .C1(new_n705), .C2(KEYINPUT47), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(G1330gat));
  OAI21_X1  g508(.A(G50gat), .B1(new_n690), .B2(new_n536), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n536), .A2(G50gat), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n676), .A2(new_n677), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT48), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  OAI211_X1 g515(.A(new_n710), .B(new_n712), .C1(new_n714), .C2(KEYINPUT48), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(G1331gat));
  NOR2_X1   g517(.A1(new_n367), .A2(new_n650), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n648), .A2(new_n719), .A3(new_n288), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n653), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n596), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n724));
  XOR2_X1   g523(.A(KEYINPUT49), .B(G64gat), .Z(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(new_n723), .B2(new_n725), .ZN(G1333gat));
  AOI21_X1  g525(.A(G71gat), .B1(new_n720), .B2(new_n665), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT110), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n648), .A2(new_n719), .A3(G71gat), .A4(new_n288), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n729), .B2(new_n646), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n720), .A2(KEYINPUT110), .A3(G71gat), .A4(new_n667), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n727), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  XOR2_X1   g531(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1334gat));
  NAND2_X1  g533(.A1(new_n720), .A2(new_n537), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G78gat), .ZN(G1335gat));
  INV_X1    g535(.A(new_n321), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n642), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT112), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n288), .B(new_n739), .C1(new_n688), .C2(new_n689), .ZN(new_n740));
  OR3_X1    g539(.A1(new_n740), .A2(KEYINPUT113), .A3(new_n591), .ZN(new_n741));
  INV_X1    g540(.A(new_n229), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT113), .B1(new_n740), .B2(new_n591), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n681), .A2(new_n745), .A3(new_n739), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n745), .B1(new_n681), .B2(new_n739), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n748), .A2(new_n653), .A3(new_n229), .A4(new_n288), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n744), .A2(new_n749), .ZN(G1336gat));
  INV_X1    g549(.A(new_n288), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n590), .A2(G92gat), .A3(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753));
  AOI22_X1  g552(.A1(new_n748), .A2(new_n752), .B1(KEYINPUT115), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(G92gat), .B1(new_n740), .B2(new_n590), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n754), .B(new_n755), .C1(KEYINPUT115), .C2(new_n753), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n681), .A2(new_n739), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT114), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n746), .B2(new_n747), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(KEYINPUT114), .A3(new_n745), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n759), .A2(new_n760), .A3(new_n752), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n755), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n756), .B1(new_n762), .B2(new_n753), .ZN(G1337gat));
  OAI21_X1  g562(.A(G99gat), .B1(new_n740), .B2(new_n646), .ZN(new_n764));
  INV_X1    g563(.A(new_n748), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n665), .A2(new_n241), .A3(new_n288), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(G1338gat));
  OAI21_X1  g566(.A(G106gat), .B1(new_n740), .B2(new_n536), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n537), .A2(new_n242), .A3(new_n288), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n768), .B(new_n769), .C1(new_n765), .C2(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(KEYINPUT116), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n759), .A2(new_n760), .A3(new_n772), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n768), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n771), .B1(new_n774), .B2(new_n769), .ZN(G1339gat));
  NAND4_X1  g574(.A1(new_n365), .A2(new_n751), .A3(new_n642), .A4(new_n366), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT117), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n277), .A2(new_n281), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n273), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n277), .A2(new_n274), .A3(new_n281), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n780), .A2(KEYINPUT54), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n207), .B1(new_n282), .B2(new_n783), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n782), .A2(KEYINPUT55), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT55), .B1(new_n782), .B2(new_n784), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n785), .A2(new_n786), .A3(new_n287), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n625), .B1(new_n630), .B2(new_n609), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n626), .B1(new_n622), .B2(new_n624), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n637), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n641), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n787), .A2(new_n677), .A3(new_n791), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n787), .A2(new_n650), .B1(new_n288), .B2(new_n791), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n792), .B1(new_n793), .B2(new_n677), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n737), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n776), .A2(new_n777), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n778), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n596), .A2(new_n591), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n599), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(G113gat), .B1(new_n802), .B2(new_n642), .ZN(new_n803));
  INV_X1    g602(.A(new_n604), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n799), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n805), .A2(new_n374), .A3(new_n650), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n803), .A2(new_n806), .ZN(G1340gat));
  AOI21_X1  g606(.A(new_n375), .B1(new_n801), .B2(new_n288), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(KEYINPUT118), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n805), .A2(new_n381), .A3(new_n288), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(G1341gat));
  AOI21_X1  g610(.A(G127gat), .B1(new_n805), .B2(new_n321), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n737), .A2(new_n378), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n812), .B1(new_n801), .B2(new_n813), .ZN(G1342gat));
  NAND3_X1  g613(.A1(new_n805), .A2(new_n352), .A3(new_n677), .ZN(new_n815));
  XOR2_X1   g614(.A(new_n815), .B(KEYINPUT56), .Z(new_n816));
  OAI21_X1  g615(.A(G134gat), .B1(new_n802), .B2(new_n680), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(G1343gat));
  NAND2_X1  g617(.A1(new_n646), .A2(new_n798), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n797), .A2(new_n537), .A3(new_n820), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n821), .A2(G141gat), .A3(new_n642), .ZN(new_n822));
  OAI21_X1  g621(.A(KEYINPUT119), .B1(new_n793), .B2(new_n677), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n641), .B(new_n790), .C1(new_n286), .C2(new_n287), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n781), .A2(KEYINPUT54), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n826), .A2(new_n282), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n282), .A2(new_n783), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n206), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n825), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n287), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n782), .A2(KEYINPUT55), .A3(new_n784), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n824), .B1(new_n833), .B2(new_n642), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT119), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n835), .A3(new_n680), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n823), .A2(new_n792), .A3(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n837), .A2(new_n838), .A3(new_n737), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n837), .B2(new_n737), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n778), .A2(new_n796), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT57), .B1(new_n842), .B2(new_n536), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n797), .A2(new_n537), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n820), .B1(new_n844), .B2(KEYINPUT57), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n843), .A2(new_n650), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n822), .B1(new_n847), .B2(G141gat), .ZN(new_n848));
  NAND2_X1  g647(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n849));
  XOR2_X1   g648(.A(new_n849), .B(KEYINPUT122), .Z(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n848), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n822), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n834), .A2(new_n835), .A3(new_n680), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n835), .B1(new_n834), .B2(new_n680), .ZN(new_n857));
  INV_X1    g656(.A(new_n792), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT120), .B1(new_n859), .B2(new_n321), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n776), .B(KEYINPUT117), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n837), .A2(new_n838), .A3(new_n737), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n855), .B1(new_n863), .B2(new_n537), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n864), .A2(new_n642), .A3(new_n845), .ZN(new_n865));
  INV_X1    g664(.A(G141gat), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n854), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n852), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n850), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n869), .ZN(G1344gat));
  NOR2_X1   g669(.A1(new_n864), .A2(new_n845), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(new_n872), .A3(new_n288), .ZN(new_n873));
  INV_X1    g672(.A(new_n821), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n872), .B1(new_n874), .B2(new_n288), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n875), .A2(G148gat), .ZN(new_n876));
  AOI211_X1 g675(.A(KEYINPUT57), .B(new_n536), .C1(new_n795), .C2(new_n776), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n877), .B1(new_n844), .B2(KEYINPUT57), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n288), .ZN(new_n879));
  OAI211_X1 g678(.A(KEYINPUT59), .B(G148gat), .C1(new_n879), .C2(new_n819), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n873), .A2(new_n876), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT123), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT123), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n873), .A2(new_n883), .A3(new_n876), .A4(new_n880), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(G1345gat));
  AOI21_X1  g684(.A(G155gat), .B1(new_n874), .B2(new_n321), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n737), .A2(new_n385), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n871), .B2(new_n887), .ZN(G1346gat));
  NAND3_X1  g687(.A1(new_n874), .A2(new_n386), .A3(new_n677), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n864), .A2(new_n680), .A3(new_n845), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n890), .B2(new_n386), .ZN(G1347gat));
  NOR2_X1   g690(.A1(new_n590), .A2(new_n653), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n797), .A2(new_n892), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n893), .A2(new_n804), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n636), .A3(new_n650), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n800), .ZN(new_n896));
  OAI21_X1  g695(.A(G169gat), .B1(new_n896), .B2(new_n642), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  XOR2_X1   g697(.A(new_n898), .B(KEYINPUT124), .Z(G1348gat));
  AOI21_X1  g698(.A(G176gat), .B1(new_n894), .B2(new_n288), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n896), .A2(new_n203), .A3(new_n751), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n900), .A2(new_n901), .ZN(G1349gat));
  NOR2_X1   g701(.A1(new_n737), .A2(new_n471), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n894), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(G183gat), .B1(new_n896), .B2(new_n737), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n906), .B1(KEYINPUT125), .B2(KEYINPUT60), .ZN(new_n907));
  NAND2_X1  g706(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n908));
  XOR2_X1   g707(.A(new_n908), .B(KEYINPUT126), .Z(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n907), .B(new_n910), .ZN(G1350gat));
  OAI21_X1  g710(.A(G190gat), .B1(new_n896), .B2(new_n680), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT61), .ZN(new_n913));
  INV_X1    g712(.A(G190gat), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n894), .A2(new_n914), .A3(new_n677), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(G1351gat));
  NAND2_X1  g715(.A1(new_n646), .A2(new_n892), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n878), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n919), .A2(new_n642), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n920), .A2(KEYINPUT127), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(KEYINPUT127), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n921), .A2(G197gat), .A3(new_n922), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n844), .A2(new_n917), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n642), .A2(G197gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(G1352gat));
  NAND3_X1  g726(.A1(new_n924), .A2(new_n205), .A3(new_n288), .ZN(new_n928));
  XOR2_X1   g727(.A(new_n928), .B(KEYINPUT62), .Z(new_n929));
  OAI21_X1  g728(.A(G204gat), .B1(new_n879), .B2(new_n917), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1353gat));
  OR3_X1    g730(.A1(new_n925), .A2(G211gat), .A3(new_n737), .ZN(new_n932));
  INV_X1    g731(.A(new_n919), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(new_n321), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n934), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n935));
  AOI21_X1  g734(.A(KEYINPUT63), .B1(new_n934), .B2(G211gat), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(G1354gat));
  AOI21_X1  g736(.A(G218gat), .B1(new_n924), .B2(new_n677), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n677), .A2(G218gat), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n933), .B2(new_n939), .ZN(G1355gat));
endmodule


