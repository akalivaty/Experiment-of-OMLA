//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 1 1 1 0 1 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT2), .ZN(new_n203));
  INV_X1    g002(.A(G148gat), .ZN(new_n204));
  INV_X1    g003(.A(G141gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT77), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT77), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G141gat), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n204), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n205), .A2(G148gat), .ZN(new_n210));
  OAI211_X1 g009(.A(KEYINPUT78), .B(new_n203), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G155gat), .B(G162gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT78), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n214), .B(new_n203), .C1(new_n209), .C2(new_n210), .ZN(new_n215));
  XNOR2_X1  g014(.A(G141gat), .B(G148gat), .ZN(new_n216));
  NOR3_X1   g015(.A1(new_n212), .A2(new_n216), .A3(KEYINPUT2), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n213), .A2(new_n218), .A3(KEYINPUT3), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT79), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n213), .A2(new_n218), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n213), .A2(new_n218), .A3(KEYINPUT79), .A4(KEYINPUT3), .ZN(new_n225));
  INV_X1    g024(.A(G120gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G113gat), .ZN(new_n227));
  INV_X1    g026(.A(G113gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G120gat), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT1), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G127gat), .B(G134gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT69), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT68), .B(G113gat), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n234), .B(new_n227), .C1(new_n235), .C2(new_n226), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n231), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n240), .A2(G113gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n228), .A2(KEYINPUT68), .ZN(new_n242));
  OAI21_X1  g041(.A(G120gat), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n234), .B1(new_n243), .B2(new_n227), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n233), .B1(new_n239), .B2(new_n244), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n221), .A2(new_n224), .A3(new_n225), .A4(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G225gat), .A2(G233gat), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n212), .A2(new_n211), .B1(new_n215), .B2(new_n217), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT4), .B1(new_n248), .B2(new_n245), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n231), .A2(new_n237), .ZN(new_n250));
  INV_X1    g049(.A(new_n227), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n228), .A2(KEYINPUT68), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n240), .A2(G113gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n251), .B1(new_n254), .B2(G120gat), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n250), .B1(new_n255), .B2(new_n234), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n243), .A2(new_n227), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT69), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n232), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(new_n222), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n249), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n247), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n259), .A2(new_n222), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n248), .A2(new_n245), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT5), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n246), .A2(new_n262), .A3(KEYINPUT5), .A4(new_n247), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G1gat), .B(G29gat), .ZN(new_n272));
  INV_X1    g071(.A(G85gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT0), .B(G57gat), .ZN(new_n275));
  XOR2_X1   g074(.A(new_n274), .B(new_n275), .Z(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n271), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT84), .ZN(new_n279));
  AOI211_X1 g078(.A(KEYINPUT39), .B(new_n247), .C1(new_n246), .C2(new_n262), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n279), .B1(new_n280), .B2(new_n276), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n246), .A2(new_n262), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(new_n264), .ZN(new_n283));
  OAI211_X1 g082(.A(KEYINPUT84), .B(new_n277), .C1(new_n283), .C2(KEYINPUT39), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT39), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n265), .A2(new_n266), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n285), .B1(new_n286), .B2(new_n247), .ZN(new_n287));
  AOI22_X1  g086(.A1(new_n281), .A2(new_n284), .B1(new_n283), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n278), .B1(new_n288), .B2(KEYINPUT40), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT40), .ZN(new_n290));
  AND2_X1   g089(.A1(new_n281), .A2(new_n284), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n283), .A2(new_n287), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G190gat), .ZN(new_n294));
  AND2_X1   g093(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT28), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT27), .B(G183gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n300), .A2(KEYINPUT28), .A3(new_n294), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT26), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NOR3_X1   g104(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G169gat), .ZN(new_n310));
  INV_X1    g109(.A(G176gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n309), .B1(KEYINPUT26), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G183gat), .A2(G190gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n302), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT67), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT24), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n315), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(G183gat), .A2(G190gat), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT67), .B1(G183gat), .B2(G190gat), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n319), .B(new_n321), .C1(new_n318), .C2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT23), .B1(new_n305), .B2(new_n306), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT23), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n309), .B1(new_n325), .B2(new_n312), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n323), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT25), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n320), .B(KEYINPUT65), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n315), .B(KEYINPUT24), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT25), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n310), .A2(new_n311), .A3(KEYINPUT23), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n325), .B1(G169gat), .B2(G176gat), .ZN(new_n334));
  AND4_X1   g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .A4(new_n308), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n316), .A2(new_n328), .A3(new_n336), .ZN(new_n337));
  XOR2_X1   g136(.A(KEYINPUT73), .B(KEYINPUT29), .Z(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n340));
  INV_X1    g139(.A(G226gat), .ZN(new_n341));
  INV_X1    g140(.A(G233gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n339), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(G211gat), .ZN(new_n346));
  INV_X1    g145(.A(G218gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(G211gat), .A2(G218gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G197gat), .B(G204gat), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT22), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  AND3_X1   g152(.A1(new_n350), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n350), .B1(new_n353), .B2(new_n351), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n337), .A2(new_n343), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT74), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n343), .B1(new_n337), .B2(new_n338), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n345), .B(new_n356), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  AND2_X1   g159(.A1(G197gat), .A2(G204gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(G197gat), .A2(G204gat), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n349), .B(new_n348), .C1(new_n363), .C2(new_n352), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n350), .A2(new_n351), .A3(new_n353), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n327), .A2(KEYINPUT25), .B1(new_n331), .B2(new_n335), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT29), .B1(new_n367), .B2(new_n316), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n357), .B(new_n366), .C1(new_n368), .C2(new_n343), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n360), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT75), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT75), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n360), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G8gat), .B(G36gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(G64gat), .B(G92gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n371), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  XOR2_X1   g177(.A(new_n376), .B(KEYINPUT76), .Z(new_n379));
  INV_X1    g178(.A(new_n373), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n372), .B1(new_n360), .B2(new_n369), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n378), .A2(new_n382), .A3(KEYINPUT30), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT30), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n371), .A2(new_n384), .A3(new_n373), .A4(new_n377), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n289), .A2(new_n293), .A3(new_n383), .A4(new_n385), .ZN(new_n386));
  XOR2_X1   g185(.A(G78gat), .B(G106gat), .Z(new_n387));
  AOI21_X1  g186(.A(KEYINPUT3), .B1(new_n366), .B2(new_n338), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT82), .B1(new_n222), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n338), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n223), .B1(new_n356), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT82), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n392), .A3(new_n248), .ZN(new_n393));
  NAND2_X1  g192(.A1(G228gat), .A2(G233gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n389), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n366), .B1(new_n224), .B2(new_n338), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT3), .B1(new_n213), .B2(new_n218), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n356), .B1(new_n398), .B2(new_n390), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n223), .B1(new_n356), .B2(KEYINPUT29), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n248), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n394), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n397), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n399), .A2(new_n401), .ZN(new_n406));
  INV_X1    g205(.A(new_n394), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n399), .A2(new_n394), .A3(new_n389), .A4(new_n393), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n403), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n387), .B1(new_n405), .B2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G22gat), .B(G50gat), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n404), .B1(new_n397), .B2(new_n402), .ZN(new_n413));
  INV_X1    g212(.A(new_n387), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n408), .A2(new_n409), .A3(new_n403), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n411), .A2(new_n412), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n412), .B1(new_n411), .B2(new_n416), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n269), .A2(KEYINPUT6), .A3(new_n276), .A4(new_n270), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(KEYINPUT81), .ZN(new_n421));
  INV_X1    g220(.A(new_n278), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT6), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n271), .A2(new_n277), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT37), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n371), .A2(new_n426), .A3(new_n373), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT37), .B1(new_n380), .B2(new_n381), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n427), .A2(new_n428), .A3(new_n376), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT38), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n421), .B(new_n425), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n427), .ZN(new_n432));
  OR2_X1    g231(.A1(new_n358), .A2(new_n359), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n433), .A2(new_n366), .A3(new_n345), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n357), .B1(new_n368), .B2(new_n343), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT37), .B1(new_n435), .B2(new_n366), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n438), .A2(new_n430), .A3(new_n379), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT85), .B1(new_n432), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n439), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT85), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(new_n442), .A3(new_n427), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n440), .A2(new_n443), .A3(new_n378), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n386), .B(new_n419), .C1(new_n431), .C2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT32), .ZN(new_n446));
  XNOR2_X1  g245(.A(G15gat), .B(G43gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(G99gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(KEYINPUT70), .B(G71gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n448), .B(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n446), .B1(new_n451), .B2(KEYINPUT33), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n337), .A2(new_n259), .ZN(new_n453));
  NAND2_X1  g252(.A1(G227gat), .A2(G233gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(KEYINPUT64), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n367), .A2(new_n245), .A3(new_n316), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n453), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n446), .A2(KEYINPUT33), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT71), .B1(new_n460), .B2(new_n451), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT71), .ZN(new_n462));
  AOI211_X1 g261(.A(new_n462), .B(new_n450), .C1(new_n457), .C2(new_n459), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n458), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT34), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n453), .A2(new_n456), .ZN(new_n466));
  INV_X1    g265(.A(new_n455), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI211_X1 g267(.A(KEYINPUT34), .B(new_n455), .C1(new_n453), .C2(new_n456), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n464), .A2(new_n471), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n470), .B(new_n458), .C1(new_n461), .C2(new_n463), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT72), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT36), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(KEYINPUT72), .A2(KEYINPUT36), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n474), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n472), .A2(new_n473), .A3(new_n475), .A4(new_n476), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n424), .A2(KEYINPUT80), .A3(new_n423), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT80), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n276), .B1(new_n269), .B2(new_n270), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n483), .B1(new_n484), .B2(KEYINPUT6), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n482), .A2(new_n422), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n421), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n383), .A2(new_n385), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n419), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n481), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n445), .A2(new_n491), .ZN(new_n492));
  NOR3_X1   g291(.A1(new_n417), .A2(new_n474), .A3(new_n418), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT35), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n425), .A2(new_n421), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n493), .A2(new_n494), .A3(new_n488), .A4(new_n495), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n486), .A2(new_n421), .B1(new_n383), .B2(new_n385), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n494), .B1(new_n497), .B2(new_n493), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n496), .B1(new_n498), .B2(KEYINPUT86), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT86), .ZN(new_n500));
  AOI211_X1 g299(.A(new_n500), .B(new_n494), .C1(new_n497), .C2(new_n493), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n492), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  OR3_X1    g301(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(G29gat), .A2(G36gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G43gat), .B(G50gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT15), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n505), .A2(KEYINPUT89), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT89), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n503), .A2(new_n513), .A3(new_n504), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT15), .ZN(new_n516));
  INV_X1    g315(.A(G50gat), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n517), .A2(G43gat), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n517), .A2(G43gat), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n516), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n506), .B(KEYINPUT90), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(new_n509), .A3(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n511), .B1(new_n515), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT17), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G15gat), .B(G22gat), .ZN(new_n526));
  INV_X1    g325(.A(G1gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT16), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(G1gat), .B2(new_n526), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(G8gat), .ZN(new_n531));
  INV_X1    g330(.A(G8gat), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n529), .B(new_n532), .C1(G1gat), .C2(new_n526), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  OAI211_X1 g334(.A(KEYINPUT17), .B(new_n511), .C1(new_n515), .C2(new_n522), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n525), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(G229gat), .A2(G233gat), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n523), .A2(new_n534), .A3(KEYINPUT91), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT91), .B1(new_n523), .B2(new_n534), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n537), .B(new_n538), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT18), .ZN(new_n542));
  OAI22_X1  g341(.A1(new_n539), .A2(new_n540), .B1(new_n523), .B2(new_n534), .ZN(new_n543));
  XOR2_X1   g342(.A(KEYINPUT92), .B(KEYINPUT13), .Z(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(new_n538), .ZN(new_n545));
  AOI22_X1  g344(.A1(new_n541), .A2(new_n542), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n539), .A2(new_n540), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n547), .A2(KEYINPUT18), .A3(new_n538), .A4(new_n537), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT12), .ZN(new_n549));
  XNOR2_X1  g348(.A(G169gat), .B(G197gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(new_n205), .ZN(new_n551));
  XOR2_X1   g350(.A(KEYINPUT87), .B(KEYINPUT11), .Z(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT88), .B(G113gat), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n553), .A2(new_n555), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n549), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n558), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n560), .A2(new_n556), .A3(KEYINPUT12), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n546), .A2(new_n548), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n562), .B1(new_n546), .B2(new_n548), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567));
  INV_X1    g366(.A(G92gat), .ZN(new_n568));
  AOI22_X1  g367(.A1(KEYINPUT8), .A2(new_n567), .B1(new_n273), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT98), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT7), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n570), .B(new_n571), .C1(new_n273), .C2(new_n568), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n570), .A2(new_n571), .ZN(new_n573));
  OAI211_X1 g372(.A(G85gat), .B(G92gat), .C1(KEYINPUT98), .C2(KEYINPUT7), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n569), .B(new_n572), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G99gat), .B(G106gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n573), .A2(new_n574), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n579), .A2(new_n576), .A3(new_n572), .A4(new_n569), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n525), .A2(new_n536), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT99), .ZN(new_n583));
  INV_X1    g382(.A(new_n581), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(new_n523), .ZN(new_n585));
  AND2_X1   g384(.A1(G232gat), .A2(G233gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT41), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n583), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n587), .ZN(new_n589));
  AOI211_X1 g388(.A(KEYINPUT99), .B(new_n589), .C1(new_n584), .C2(new_n523), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n582), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G190gat), .B(G218gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n586), .A2(KEYINPUT41), .ZN(new_n594));
  XNOR2_X1  g393(.A(G134gat), .B(G162gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n596), .A2(KEYINPUT100), .ZN(new_n597));
  INV_X1    g396(.A(new_n592), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n582), .B(new_n598), .C1(new_n588), .C2(new_n590), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n593), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n596), .B(KEYINPUT100), .Z(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n602), .B1(new_n593), .B2(new_n599), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G183gat), .B(G211gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n605), .B(new_n606), .Z(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT95), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT93), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n612), .B1(G71gat), .B2(G78gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(G57gat), .B(G64gat), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G71gat), .B(G78gat), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT9), .ZN(new_n620));
  INV_X1    g419(.A(G71gat), .ZN(new_n621));
  INV_X1    g420(.A(G78gat), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OR2_X1    g422(.A1(G57gat), .A2(G64gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(G57gat), .A2(G64gat), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n617), .B1(new_n626), .B2(new_n613), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT94), .ZN(new_n628));
  NOR3_X1   g427(.A1(new_n619), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n616), .A2(new_n618), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n626), .A2(new_n617), .A3(new_n613), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT94), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n611), .B1(new_n629), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n628), .B1(new_n619), .B2(new_n627), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n630), .A2(KEYINPUT94), .A3(new_n631), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(KEYINPUT95), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n633), .A2(KEYINPUT21), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(G231gat), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(new_n342), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n637), .A2(new_n535), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n640), .B1(new_n637), .B2(new_n535), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n610), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n637), .A2(new_n535), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n639), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n637), .A2(new_n535), .A3(new_n640), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(new_n609), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT21), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n648), .B1(new_n629), .B2(new_n632), .ZN(new_n649));
  XOR2_X1   g448(.A(G127gat), .B(G155gat), .Z(new_n650));
  XOR2_X1   g449(.A(new_n649), .B(new_n650), .Z(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n643), .A2(new_n647), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n652), .B1(new_n643), .B2(new_n647), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n608), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n643), .A2(new_n647), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n651), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n643), .A2(new_n647), .A3(new_n652), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(new_n607), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n604), .B1(new_n655), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(G230gat), .A2(G233gat), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT10), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n581), .A2(new_n662), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n633), .A2(new_n636), .A3(new_n663), .ZN(new_n664));
  AOI22_X1  g463(.A1(new_n634), .A2(new_n635), .B1(new_n580), .B2(new_n578), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n619), .A2(new_n627), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n666), .A2(new_n581), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n665), .A2(KEYINPUT10), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n661), .B1(new_n664), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n581), .B1(new_n629), .B2(new_n632), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n666), .A2(new_n581), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n661), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  XOR2_X1   g472(.A(G176gat), .B(G204gat), .Z(new_n674));
  XNOR2_X1  g473(.A(G120gat), .B(G148gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n669), .A2(new_n673), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n678), .B1(new_n669), .B2(new_n673), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AND4_X1   g481(.A1(new_n502), .A2(new_n566), .A3(new_n660), .A4(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n487), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(G1gat), .ZN(G1324gat));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n687));
  INV_X1    g486(.A(new_n488), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT103), .B(KEYINPUT16), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G8gat), .ZN(new_n692));
  AOI21_X1  g491(.A(KEYINPUT42), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n690), .A2(new_n692), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n689), .A2(G8gat), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT42), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n687), .B(new_n694), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n698), .B1(new_n695), .B2(new_n696), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT104), .B1(new_n700), .B2(new_n693), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(G1325gat));
  INV_X1    g501(.A(new_n474), .ZN(new_n703));
  AOI21_X1  g502(.A(G15gat), .B1(new_n683), .B2(new_n703), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n481), .A2(G15gat), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n704), .B1(new_n683), .B2(new_n705), .ZN(G1326gat));
  NAND2_X1  g505(.A1(new_n683), .A2(new_n490), .ZN(new_n707));
  XNOR2_X1  g506(.A(KEYINPUT43), .B(G22gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1327gat));
  AND2_X1   g508(.A1(new_n502), .A2(new_n604), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n655), .A2(new_n659), .ZN(new_n711));
  INV_X1    g510(.A(new_n682), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n711), .A2(new_n712), .A3(new_n565), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(G29gat), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n714), .A2(new_n715), .A3(new_n684), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT45), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718));
  AND3_X1   g517(.A1(new_n502), .A2(new_n718), .A3(new_n604), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n718), .B1(new_n502), .B2(new_n604), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n713), .ZN(new_n722));
  OAI21_X1  g521(.A(G29gat), .B1(new_n722), .B2(new_n487), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n717), .A2(new_n723), .ZN(G1328gat));
  INV_X1    g523(.A(G36gat), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n714), .A2(new_n725), .A3(new_n688), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(KEYINPUT46), .Z(new_n727));
  OAI21_X1  g526(.A(G36gat), .B1(new_n722), .B2(new_n488), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(G1329gat));
  OAI211_X1 g528(.A(new_n481), .B(new_n713), .C1(new_n719), .C2(new_n720), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G43gat), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT105), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n730), .A2(new_n733), .A3(G43gat), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n474), .A2(G43gat), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n710), .A2(new_n713), .A3(new_n735), .ZN(new_n736));
  AND3_X1   g535(.A1(new_n732), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT106), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n736), .A2(KEYINPUT47), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n738), .B1(new_n731), .B2(new_n739), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n731), .A2(new_n739), .A3(new_n738), .ZN(new_n741));
  OAI22_X1  g540(.A1(new_n737), .A2(KEYINPUT47), .B1(new_n740), .B2(new_n741), .ZN(G1330gat));
  OAI21_X1  g541(.A(G50gat), .B1(new_n722), .B2(new_n419), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n714), .A2(new_n517), .A3(new_n490), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT48), .B1(new_n744), .B2(KEYINPUT107), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n743), .B(new_n744), .C1(KEYINPUT107), .C2(KEYINPUT48), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(G1331gat));
  INV_X1    g548(.A(new_n711), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n712), .A2(new_n565), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n750), .A2(new_n604), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n502), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n684), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g555(.A1(new_n753), .A2(new_n488), .ZN(new_n757));
  NOR2_X1   g556(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n758));
  AND2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n757), .B2(new_n758), .ZN(G1333gat));
  INV_X1    g560(.A(new_n481), .ZN(new_n762));
  OAI21_X1  g561(.A(G71gat), .B1(new_n753), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n703), .A2(new_n621), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n763), .B1(new_n753), .B2(new_n764), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g565(.A1(new_n753), .A2(new_n419), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(new_n622), .ZN(G1335gat));
  NOR2_X1   g567(.A1(new_n711), .A2(new_n751), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n721), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(G85gat), .B1(new_n770), .B2(new_n487), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n502), .A2(new_n772), .A3(new_n604), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n711), .A2(new_n566), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n772), .B1(new_n502), .B2(new_n604), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT51), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n502), .A2(new_n604), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT108), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n779), .A2(new_n780), .A3(new_n773), .A4(new_n774), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n487), .A2(G85gat), .A3(new_n682), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n777), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n771), .A2(new_n783), .ZN(G1336gat));
  NAND3_X1  g583(.A1(new_n721), .A2(new_n688), .A3(new_n769), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G92gat), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n488), .A2(G92gat), .A3(new_n682), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n777), .A2(new_n781), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n786), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(new_n775), .B2(new_n776), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n780), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n791), .B(KEYINPUT51), .C1(new_n775), .C2(new_n776), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n793), .A2(new_n794), .A3(new_n788), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n795), .A2(new_n786), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n790), .B1(new_n796), .B2(new_n787), .ZN(G1337gat));
  OAI21_X1  g596(.A(G99gat), .B1(new_n770), .B2(new_n762), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n474), .A2(G99gat), .A3(new_n682), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n777), .A2(new_n781), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(G1338gat));
  OAI211_X1 g600(.A(new_n490), .B(new_n769), .C1(new_n719), .C2(new_n720), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT53), .B1(new_n802), .B2(G106gat), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n419), .A2(G106gat), .A3(new_n682), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n777), .A2(new_n781), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT110), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT110), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n803), .A2(new_n805), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n793), .A2(new_n794), .A3(new_n804), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n802), .A2(G106gat), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT53), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n810), .A2(new_n814), .ZN(G1339gat));
  INV_X1    g614(.A(new_n604), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n670), .A2(new_n671), .A3(new_n662), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n633), .A2(new_n636), .A3(new_n663), .ZN(new_n818));
  INV_X1    g617(.A(new_n661), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n669), .A2(KEYINPUT54), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n819), .B1(new_n817), .B2(new_n818), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n678), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n821), .A2(new_n824), .A3(KEYINPUT55), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n825), .A2(new_n679), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n821), .A2(new_n824), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n826), .A2(KEYINPUT111), .A3(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT111), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n825), .A2(new_n679), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT55), .B1(new_n821), .B2(new_n824), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n565), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n538), .B1(new_n547), .B2(new_n537), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n543), .A2(new_n545), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n560), .B(new_n556), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n546), .A2(new_n548), .A3(new_n562), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n682), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n816), .B1(new_n835), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n830), .A2(new_n834), .ZN(new_n843));
  INV_X1    g642(.A(new_n840), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(new_n604), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n711), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n711), .A2(new_n565), .A3(new_n816), .A4(new_n682), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n849), .A2(new_n493), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n688), .A2(new_n487), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n566), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(G113gat), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n855), .B1(new_n235), .B2(new_n854), .ZN(G1340gat));
  OAI22_X1  g655(.A1(new_n852), .A2(new_n682), .B1(KEYINPUT112), .B2(G120gat), .ZN(new_n857));
  NAND2_X1  g656(.A1(KEYINPUT112), .A2(G120gat), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT113), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n857), .B(new_n859), .ZN(G1341gat));
  NAND2_X1  g659(.A1(new_n853), .A2(new_n711), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n861), .B(G127gat), .ZN(G1342gat));
  NOR2_X1   g661(.A1(new_n852), .A2(new_n816), .ZN(new_n863));
  INV_X1    g662(.A(G134gat), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n865), .A2(KEYINPUT56), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(KEYINPUT56), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n866), .B(new_n867), .C1(new_n864), .C2(new_n863), .ZN(G1343gat));
  INV_X1    g667(.A(KEYINPUT58), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n851), .A2(new_n762), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n849), .A2(new_n490), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n565), .A2(G141gat), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n869), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n206), .A2(new_n208), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n849), .A2(new_n877), .A3(new_n490), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n825), .B(new_n679), .C1(new_n563), .C2(new_n564), .ZN(new_n879));
  AOI21_X1  g678(.A(KEYINPUT114), .B1(new_n827), .B2(new_n828), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT114), .ZN(new_n881));
  AOI211_X1 g680(.A(new_n881), .B(KEYINPUT55), .C1(new_n821), .C2(new_n824), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n816), .B1(new_n883), .B2(new_n841), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n711), .B1(new_n845), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n490), .B1(new_n885), .B2(new_n848), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n870), .B1(new_n886), .B2(KEYINPUT57), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n878), .A2(new_n566), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n875), .B1(new_n876), .B2(new_n888), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT116), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n878), .A2(KEYINPUT115), .A3(new_n887), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT115), .B1(new_n878), .B2(new_n887), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n566), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n872), .ZN(new_n894));
  AOI22_X1  g693(.A1(new_n893), .A2(new_n876), .B1(new_n894), .B2(new_n873), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n890), .B1(new_n895), .B2(new_n869), .ZN(G1344gat));
  NAND3_X1  g695(.A1(new_n894), .A2(new_n204), .A3(new_n712), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(G148gat), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n891), .A2(new_n892), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(new_n712), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n847), .A2(KEYINPUT117), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT117), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n660), .A2(new_n903), .A3(new_n565), .A4(new_n682), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n604), .A2(new_n829), .A3(new_n679), .A4(new_n825), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT118), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n826), .A2(KEYINPUT118), .A3(new_n604), .A4(new_n829), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n844), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n711), .B1(new_n884), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n490), .B1(new_n905), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(KEYINPUT119), .A3(new_n877), .ZN(new_n913));
  OAI211_X1 g712(.A(KEYINPUT57), .B(new_n490), .C1(new_n846), .C2(new_n848), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(KEYINPUT119), .B1(new_n912), .B2(new_n877), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n917), .A2(new_n712), .A3(new_n871), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n898), .B1(new_n918), .B2(G148gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n897), .B1(new_n901), .B2(new_n919), .ZN(G1345gat));
  AOI21_X1  g719(.A(G155gat), .B1(new_n894), .B2(new_n711), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n711), .A2(G155gat), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n921), .B1(new_n900), .B2(new_n922), .ZN(G1346gat));
  NAND2_X1  g722(.A1(new_n900), .A2(new_n604), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G162gat), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n816), .A2(G162gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n872), .B2(new_n926), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n684), .A2(new_n488), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n493), .B(new_n928), .C1(new_n846), .C2(new_n848), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT120), .ZN(new_n930));
  OAI21_X1  g729(.A(G169gat), .B1(new_n930), .B2(new_n565), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT121), .ZN(new_n932));
  INV_X1    g731(.A(new_n929), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n310), .A3(new_n566), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1348gat));
  OR3_X1    g734(.A1(new_n930), .A2(new_n311), .A3(new_n682), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n936), .A2(KEYINPUT123), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(KEYINPUT123), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n311), .B1(new_n929), .B2(new_n682), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT122), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n937), .A2(new_n938), .A3(new_n940), .ZN(G1349gat));
  OAI21_X1  g740(.A(G183gat), .B1(new_n930), .B2(new_n750), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n933), .A2(new_n300), .A3(new_n711), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g744(.A1(new_n933), .A2(new_n294), .A3(new_n604), .ZN(new_n946));
  OAI21_X1  g745(.A(G190gat), .B1(new_n930), .B2(new_n816), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT124), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT61), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n949), .B1(KEYINPUT61), .B2(new_n947), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n948), .B1(new_n947), .B2(KEYINPUT61), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n946), .B1(new_n950), .B2(new_n951), .ZN(G1351gat));
  NAND2_X1  g751(.A1(new_n928), .A2(new_n762), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n917), .A2(new_n566), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(G197gat), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n849), .A2(new_n490), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(new_n954), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n565), .A2(G197gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(G1352gat));
  NAND3_X1  g759(.A1(new_n917), .A2(new_n712), .A3(new_n954), .ZN(new_n961));
  XOR2_X1   g760(.A(KEYINPUT125), .B(G204gat), .Z(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(new_n958), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n682), .A2(new_n962), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(KEYINPUT62), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT62), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n964), .A2(new_n968), .A3(new_n965), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT126), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  OAI211_X1 g771(.A(new_n963), .B(new_n967), .C1(new_n971), .C2(new_n972), .ZN(G1353gat));
  NAND3_X1  g772(.A1(new_n964), .A2(new_n346), .A3(new_n711), .ZN(new_n974));
  OAI211_X1 g773(.A(new_n711), .B(new_n954), .C1(new_n915), .C2(new_n916), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n975), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n976));
  AOI21_X1  g775(.A(KEYINPUT63), .B1(new_n975), .B2(G211gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n978), .A2(KEYINPUT127), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT127), .ZN(new_n980));
  OAI211_X1 g779(.A(new_n980), .B(new_n974), .C1(new_n976), .C2(new_n977), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n979), .A2(new_n981), .ZN(G1354gat));
  NAND4_X1  g781(.A1(new_n917), .A2(G218gat), .A3(new_n604), .A4(new_n954), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n347), .B1(new_n958), .B2(new_n816), .ZN(new_n984));
  AND2_X1   g783(.A1(new_n983), .A2(new_n984), .ZN(G1355gat));
endmodule


