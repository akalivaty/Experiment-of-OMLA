//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 0 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012;
  INV_X1    g000(.A(G211gat), .ZN(new_n202));
  INV_X1    g001(.A(G218gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G211gat), .A2(G218gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT74), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT74), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n204), .A2(new_n208), .A3(new_n205), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT73), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G197gat), .B(G204gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n211), .A2(new_n212), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n210), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n211), .B(KEYINPUT73), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n218), .A2(new_n214), .A3(new_n207), .A4(new_n209), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT75), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n217), .A2(new_n219), .A3(KEYINPUT75), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT2), .ZN(new_n225));
  INV_X1    g024(.A(G141gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G148gat), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n226), .A2(G148gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n225), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G155gat), .B(G162gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G155gat), .ZN(new_n234));
  INV_X1    g033(.A(G162gat), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT2), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT80), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n236), .B(new_n237), .ZN(new_n238));
  OR2_X1    g037(.A1(KEYINPUT79), .A2(G148gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(KEYINPUT79), .A2(G148gat), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n226), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n231), .B1(new_n241), .B2(new_n228), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n233), .B1(new_n238), .B2(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n243), .A2(KEYINPUT3), .ZN(new_n244));
  XOR2_X1   g043(.A(KEYINPUT76), .B(KEYINPUT29), .Z(new_n245));
  OAI21_X1  g044(.A(new_n224), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n245), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n243), .A2(new_n247), .A3(new_n219), .A4(new_n217), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n243), .A2(KEYINPUT3), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT88), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n248), .A2(KEYINPUT88), .A3(new_n249), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n246), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(G228gat), .A2(G233gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G22gat), .ZN(new_n257));
  INV_X1    g056(.A(new_n255), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n259), .B1(new_n220), .B2(KEYINPUT29), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n243), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n246), .A2(new_n258), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n256), .A2(new_n257), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT89), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n256), .A2(new_n262), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G22gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT89), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n256), .A2(new_n267), .A3(new_n257), .A4(new_n262), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n264), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(G78gat), .B(G106gat), .Z(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(G50gat), .ZN(new_n271));
  XOR2_X1   g070(.A(KEYINPUT87), .B(KEYINPUT31), .Z(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT91), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n273), .B1(new_n263), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT90), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n277), .B(G22gat), .C1(new_n265), .C2(new_n275), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(G22gat), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n256), .A2(KEYINPUT91), .A3(new_n262), .A4(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n276), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n274), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G183gat), .A2(G190gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n284));
  INV_X1    g083(.A(G169gat), .ZN(new_n285));
  INV_X1    g084(.A(G176gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT26), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT26), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n283), .B1(new_n289), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT66), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g095(.A(KEYINPUT66), .B(new_n283), .C1(new_n289), .C2(new_n293), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT27), .B(G183gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT28), .B1(new_n300), .B2(G190gat), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT28), .ZN(new_n302));
  INV_X1    g101(.A(G190gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n299), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n283), .A2(KEYINPUT24), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT24), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n307), .B1(G183gat), .B2(G190gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n306), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT23), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT64), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT64), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT23), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n291), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n291), .A2(KEYINPUT23), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n311), .A2(new_n318), .A3(new_n319), .A4(new_n290), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT25), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n307), .A2(G183gat), .A3(G190gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n283), .A2(KEYINPUT24), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n323), .B1(new_n324), .B2(new_n309), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n291), .B1(new_n313), .B2(new_n315), .ZN(new_n326));
  INV_X1    g125(.A(new_n290), .ZN(new_n327));
  NOR3_X1   g126(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n287), .A2(new_n288), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n321), .B1(new_n329), .B2(KEYINPUT23), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n298), .A2(new_n305), .B1(new_n322), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G127gat), .B(G134gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G113gat), .B(G120gat), .ZN(new_n335));
  NOR3_X1   g134(.A1(new_n334), .A2(KEYINPUT1), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT1), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT67), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n337), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(G120gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G113gat), .ZN(new_n341));
  INV_X1    g140(.A(G113gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G120gat), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n343), .A3(new_n338), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n334), .B1(new_n339), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT68), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n342), .A2(G120gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n340), .A2(G113gat), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT67), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n350), .A2(new_n337), .A3(new_n344), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT68), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(new_n352), .A3(new_n334), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n336), .B1(new_n347), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT69), .B1(new_n332), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n332), .A2(new_n354), .ZN(new_n356));
  INV_X1    g155(.A(new_n336), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n343), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT1), .B1(new_n358), .B2(KEYINPUT67), .ZN(new_n359));
  AOI211_X1 g158(.A(KEYINPUT68), .B(new_n333), .C1(new_n359), .C2(new_n344), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n352), .B1(new_n351), .B2(new_n334), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n357), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT69), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n321), .A2(new_n320), .B1(new_n328), .B2(new_n330), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n301), .A2(new_n304), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n365), .B1(new_n296), .B2(new_n297), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n362), .B(new_n363), .C1(new_n364), .C2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n355), .A2(new_n356), .A3(new_n367), .ZN(new_n368));
  AND2_X1   g167(.A1(G227gat), .A2(G233gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  XOR2_X1   g169(.A(new_n370), .B(KEYINPUT34), .Z(new_n371));
  INV_X1    g170(.A(KEYINPUT32), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n372), .B1(new_n368), .B2(new_n369), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT33), .B1(new_n368), .B2(new_n369), .ZN(new_n374));
  XNOR2_X1  g173(.A(G15gat), .B(G43gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n375), .B(G71gat), .ZN(new_n376));
  INV_X1    g175(.A(G99gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NOR3_X1   g178(.A1(new_n373), .A2(new_n374), .A3(new_n379), .ZN(new_n380));
  AOI221_X4 g179(.A(new_n372), .B1(KEYINPUT33), .B2(new_n378), .C1(new_n368), .C2(new_n369), .ZN(new_n381));
  NOR3_X1   g180(.A1(new_n380), .A2(KEYINPUT70), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT70), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n369), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT32), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT33), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n387), .A3(new_n378), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n373), .B1(new_n374), .B2(new_n379), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n383), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n371), .B1(new_n382), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT71), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n388), .A2(new_n389), .ZN(new_n394));
  OR2_X1    g193(.A1(new_n394), .A2(new_n371), .ZN(new_n395));
  OAI211_X1 g194(.A(KEYINPUT71), .B(new_n371), .C1(new_n382), .C2(new_n390), .ZN(new_n396));
  AND4_X1   g195(.A1(new_n282), .A2(new_n393), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G1gat), .B(G29gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n398), .B(G85gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT0), .B(G57gat), .ZN(new_n400));
  XOR2_X1   g199(.A(new_n399), .B(new_n400), .Z(new_n401));
  XNOR2_X1  g200(.A(KEYINPUT79), .B(G148gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(G141gat), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n232), .B1(new_n403), .B2(new_n227), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n236), .B(KEYINPUT80), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n404), .A2(new_n405), .B1(new_n232), .B2(new_n230), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n259), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n362), .A2(new_n407), .A3(new_n249), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT81), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT81), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n362), .A2(new_n407), .A3(new_n410), .A4(new_n249), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n406), .B(new_n357), .C1(new_n360), .C2(new_n361), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT4), .ZN(new_n414));
  NAND2_X1  g213(.A1(G225gat), .A2(G233gat), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n416), .A2(KEYINPUT5), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n412), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT82), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n419), .B1(new_n413), .B2(KEYINPUT4), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n413), .A2(KEYINPUT4), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT4), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n354), .A2(KEYINPUT82), .A3(new_n422), .A4(new_n406), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n412), .A2(new_n424), .A3(new_n415), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n362), .A2(new_n243), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT83), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n427), .A3(new_n413), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n362), .A2(KEYINPUT83), .A3(new_n243), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n416), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT5), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n401), .B(new_n418), .C1(new_n425), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT84), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT6), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n412), .A2(new_n424), .A3(new_n415), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n435), .A2(KEYINPUT5), .A3(new_n430), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT84), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n436), .A2(new_n437), .A3(new_n401), .A4(new_n418), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n433), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT85), .ZN(new_n440));
  AOI211_X1 g239(.A(new_n440), .B(new_n401), .C1(new_n436), .C2(new_n418), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n418), .B1(new_n425), .B2(new_n431), .ZN(new_n442));
  INV_X1    g241(.A(new_n401), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT85), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT86), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n439), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n430), .A2(KEYINPUT5), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n412), .A2(new_n414), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n448), .A2(new_n435), .B1(new_n449), .B2(new_n417), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n440), .B1(new_n450), .B2(new_n401), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n442), .A2(KEYINPUT85), .A3(new_n443), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n433), .A2(new_n434), .A3(new_n438), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT86), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n450), .A2(new_n401), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT6), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n447), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(G8gat), .B(G36gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(G64gat), .B(G92gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n459), .B(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(G226gat), .A2(G233gat), .ZN(new_n462));
  INV_X1    g261(.A(new_n288), .ZN(new_n463));
  NOR3_X1   g262(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n292), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n293), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT66), .B1(new_n467), .B2(new_n283), .ZN(new_n468));
  INV_X1    g267(.A(new_n297), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n305), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n322), .A2(new_n331), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n462), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n247), .B1(new_n366), .B2(new_n364), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n472), .B1(new_n462), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT77), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n222), .A2(new_n223), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n462), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n478), .B1(new_n366), .B2(new_n364), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n245), .B1(new_n470), .B2(new_n471), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n479), .B1(new_n480), .B2(new_n478), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT77), .B1(new_n481), .B2(new_n224), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT29), .B1(new_n470), .B2(new_n471), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n479), .B(new_n476), .C1(new_n484), .C2(new_n478), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT78), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n461), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n485), .B(KEYINPUT78), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n475), .B1(new_n474), .B2(new_n476), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n481), .A2(KEYINPUT77), .A3(new_n224), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n461), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n489), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n488), .A2(KEYINPUT30), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT30), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n489), .A2(new_n492), .A3(new_n496), .A4(new_n493), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n397), .A2(KEYINPUT35), .A3(new_n458), .A4(new_n498), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n495), .A2(new_n497), .A3(KEYINPUT93), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT93), .B1(new_n495), .B2(new_n497), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n394), .B(new_n371), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n442), .A2(new_n443), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n433), .A2(new_n505), .A3(new_n434), .A4(new_n438), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n457), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n502), .A2(new_n282), .A3(new_n504), .A4(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT35), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n506), .A2(new_n457), .A3(new_n494), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT37), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n489), .A2(new_n492), .A3(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n479), .B(new_n224), .C1(new_n484), .C2(new_n478), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n514), .B(KEYINPUT37), .C1(new_n474), .C2(new_n224), .ZN(new_n515));
  XOR2_X1   g314(.A(KEYINPUT95), .B(KEYINPUT38), .Z(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  AND4_X1   g316(.A1(new_n461), .A2(new_n513), .A3(new_n515), .A4(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT96), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT37), .B1(new_n483), .B2(new_n487), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n521), .A2(new_n461), .A3(new_n513), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n518), .A2(new_n519), .B1(new_n522), .B2(new_n516), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n511), .A2(new_n520), .A3(new_n523), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n428), .A2(new_n429), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT39), .B1(new_n525), .B2(new_n416), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n412), .A2(new_n414), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n526), .B1(new_n416), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT94), .B(KEYINPUT39), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n527), .A2(new_n416), .A3(new_n529), .ZN(new_n530));
  NOR3_X1   g329(.A1(new_n528), .A2(new_n443), .A3(new_n530), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n531), .A2(KEYINPUT40), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n456), .B1(new_n531), .B2(KEYINPUT40), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n532), .B(new_n533), .C1(new_n500), .C2(new_n501), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n524), .A2(new_n534), .A3(new_n282), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n393), .A2(KEYINPUT36), .A3(new_n395), .A4(new_n396), .ZN(new_n536));
  XNOR2_X1  g335(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n503), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n282), .B(KEYINPUT92), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n541), .B1(new_n458), .B2(new_n498), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n499), .B(new_n510), .C1(new_n540), .C2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT18), .ZN(new_n544));
  XOR2_X1   g343(.A(G43gat), .B(G50gat), .Z(new_n545));
  INV_X1    g344(.A(KEYINPUT97), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G43gat), .B(G50gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT97), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n547), .A2(KEYINPUT15), .A3(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(KEYINPUT98), .B(KEYINPUT15), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n545), .A2(new_n551), .B1(G29gat), .B2(G36gat), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NOR3_X1   g353(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT99), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n550), .B(new_n552), .C1(new_n554), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G29gat), .A2(G36gat), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n558), .B1(new_n554), .B2(new_n555), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n547), .A2(new_n559), .A3(KEYINPUT15), .A4(new_n549), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT17), .ZN(new_n562));
  XNOR2_X1  g361(.A(G15gat), .B(G22gat), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT16), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n564), .A2(G1gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(G1gat), .B2(new_n563), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n567), .A2(G8gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(G8gat), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n562), .A2(new_n570), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n557), .A2(new_n560), .ZN(new_n572));
  OR2_X1    g371(.A1(new_n572), .A2(new_n570), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G229gat), .A2(G233gat), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n544), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n572), .A2(new_n570), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n575), .B(KEYINPUT13), .Z(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n571), .A2(KEYINPUT18), .A3(new_n573), .A4(new_n575), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n577), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G113gat), .B(G141gat), .ZN(new_n584));
  INV_X1    g383(.A(G197gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT11), .B(G169gat), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n586), .B(new_n587), .Z(new_n588));
  XOR2_X1   g387(.A(new_n588), .B(KEYINPUT12), .Z(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n583), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n583), .A2(new_n590), .ZN(new_n592));
  AND3_X1   g391(.A1(new_n591), .A2(KEYINPUT100), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT100), .B1(new_n591), .B2(new_n592), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(G99gat), .A2(G106gat), .ZN(new_n597));
  INV_X1    g396(.A(G85gat), .ZN(new_n598));
  INV_X1    g397(.A(G92gat), .ZN(new_n599));
  AOI22_X1  g398(.A1(KEYINPUT8), .A2(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT103), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G85gat), .A2(G92gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT7), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G99gat), .B(G106gat), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n596), .B1(new_n607), .B2(new_n572), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT104), .ZN(new_n609));
  XNOR2_X1  g408(.A(G190gat), .B(G218gat), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n610), .B(KEYINPUT105), .Z(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n562), .A2(new_n607), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n609), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT106), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n609), .A2(new_n613), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT107), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n617), .A2(new_n618), .A3(new_n611), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n609), .A2(new_n613), .ZN(new_n620));
  OAI21_X1  g419(.A(KEYINPUT107), .B1(new_n620), .B2(new_n612), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n616), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G134gat), .B(G162gat), .Z(new_n623));
  AOI21_X1  g422(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT102), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n621), .A2(new_n619), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n625), .B1(new_n620), .B2(new_n612), .ZN(new_n628));
  AOI22_X1  g427(.A1(new_n622), .A2(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G127gat), .B(G155gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G211gat), .ZN(new_n631));
  INV_X1    g430(.A(G231gat), .ZN(new_n632));
  INV_X1    g431(.A(G233gat), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(G71gat), .A2(G78gat), .ZN(new_n636));
  OR2_X1    g435(.A1(G71gat), .A2(G78gat), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT9), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(G64gat), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT101), .ZN(new_n641));
  INV_X1    g440(.A(G57gat), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(KEYINPUT101), .A2(G57gat), .A3(G64gat), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n639), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(KEYINPUT9), .B1(new_n642), .B2(new_n640), .ZN(new_n646));
  NOR2_X1   g445(.A1(G57gat), .A2(G64gat), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n636), .B(new_n637), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(KEYINPUT21), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n570), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(G183gat), .ZN(new_n653));
  INV_X1    g452(.A(G183gat), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n570), .A2(new_n654), .A3(new_n651), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n650), .A2(KEYINPUT21), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n657), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n659), .B1(new_n653), .B2(new_n655), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n635), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n658), .A2(new_n635), .A3(new_n660), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n631), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n658), .A2(new_n660), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n634), .ZN(new_n667));
  INV_X1    g466(.A(new_n631), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(new_n661), .A3(new_n668), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n664), .A2(new_n665), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n665), .B1(new_n664), .B2(new_n669), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(G230gat), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n633), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n649), .B(KEYINPUT108), .Z(new_n675));
  NOR2_X1   g474(.A1(new_n649), .A2(KEYINPUT108), .ZN(new_n676));
  MUX2_X1   g475(.A(new_n675), .B(new_n676), .S(new_n607), .Z(new_n677));
  INV_X1    g476(.A(KEYINPUT10), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OR3_X1    g478(.A1(new_n607), .A2(new_n678), .A3(new_n649), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n674), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n674), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n677), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(G120gat), .B(G148gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(G176gat), .B(G204gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n682), .A2(new_n684), .A3(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n684), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n687), .B1(new_n690), .B2(new_n681), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n629), .A2(new_n672), .A3(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n543), .A2(new_n595), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT109), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT109), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n543), .A2(new_n697), .A3(new_n595), .A4(new_n694), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n458), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(G1gat), .ZN(G1324gat));
  INV_X1    g501(.A(new_n502), .ZN(new_n703));
  INV_X1    g502(.A(G8gat), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n564), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n699), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n564), .A2(new_n704), .ZN(new_n708));
  OR3_X1    g507(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n699), .ZN(new_n710));
  OAI21_X1  g509(.A(G8gat), .B1(new_n710), .B2(new_n502), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n707), .B1(new_n706), .B2(new_n708), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n709), .A2(new_n711), .A3(new_n712), .ZN(G1325gat));
  AOI21_X1  g512(.A(G15gat), .B1(new_n699), .B2(new_n504), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n710), .A2(new_n539), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n714), .B1(new_n715), .B2(G15gat), .ZN(G1326gat));
  XNOR2_X1  g515(.A(KEYINPUT110), .B(KEYINPUT43), .ZN(new_n717));
  INV_X1    g516(.A(new_n541), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n257), .B1(new_n699), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  AOI211_X1 g519(.A(G22gat), .B(new_n541), .C1(new_n696), .C2(new_n698), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n717), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n717), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n719), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n723), .A2(new_n725), .ZN(G1327gat));
  INV_X1    g525(.A(KEYINPUT113), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n622), .A2(new_n626), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n627), .A2(new_n628), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n629), .A2(new_n727), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n543), .A2(new_n736), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n458), .A2(KEYINPUT35), .A3(new_n498), .ZN(new_n738));
  AOI22_X1  g537(.A1(new_n738), .A2(new_n397), .B1(new_n509), .B2(new_n508), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n458), .A2(new_n498), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n718), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n741), .A2(new_n539), .A3(new_n535), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n629), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n737), .B1(new_n743), .B2(new_n734), .ZN(new_n744));
  XOR2_X1   g543(.A(new_n692), .B(KEYINPUT111), .Z(new_n745));
  NAND2_X1  g544(.A1(new_n591), .A2(new_n592), .ZN(new_n746));
  INV_X1    g545(.A(new_n672), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  XOR2_X1   g547(.A(new_n748), .B(KEYINPUT112), .Z(new_n749));
  NAND3_X1  g548(.A1(new_n744), .A2(new_n700), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G29gat), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT45), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n672), .A2(new_n692), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n743), .A2(new_n595), .A3(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(new_n458), .ZN(new_n755));
  INV_X1    g554(.A(G29gat), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n752), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NOR4_X1   g556(.A1(new_n754), .A2(KEYINPUT45), .A3(G29gat), .A4(new_n458), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n751), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT114), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n751), .B(KEYINPUT114), .C1(new_n757), .C2(new_n758), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(G1328gat));
  NOR3_X1   g562(.A1(new_n754), .A2(G36gat), .A3(new_n502), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT46), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n744), .A2(new_n703), .A3(new_n749), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G36gat), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n764), .A2(new_n765), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n766), .A2(new_n768), .A3(new_n769), .ZN(G1329gat));
  INV_X1    g569(.A(new_n539), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n744), .A2(new_n771), .A3(new_n749), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n744), .A2(KEYINPUT115), .A3(new_n771), .A4(new_n749), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n774), .A2(new_n775), .A3(G43gat), .ZN(new_n776));
  OR3_X1    g575(.A1(new_n754), .A2(G43gat), .A3(new_n503), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n776), .A2(KEYINPUT47), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n772), .A2(G43gat), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n777), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT47), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n778), .A2(new_n782), .ZN(G1330gat));
  INV_X1    g582(.A(new_n282), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n744), .A2(new_n784), .A3(new_n749), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n754), .A2(G50gat), .ZN(new_n786));
  AOI22_X1  g585(.A1(new_n785), .A2(G50gat), .B1(new_n786), .B2(new_n718), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT48), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n744), .A2(new_n718), .A3(new_n749), .ZN(new_n789));
  AOI22_X1  g588(.A1(new_n789), .A2(G50gat), .B1(new_n786), .B2(new_n718), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(KEYINPUT48), .B2(new_n790), .ZN(G1331gat));
  INV_X1    g590(.A(new_n745), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n728), .A2(new_n729), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n793), .A2(new_n747), .A3(new_n746), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n543), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n700), .ZN(new_n796));
  XOR2_X1   g595(.A(KEYINPUT116), .B(G57gat), .Z(new_n797));
  XNOR2_X1  g596(.A(new_n796), .B(new_n797), .ZN(G1332gat));
  NAND2_X1  g597(.A1(new_n795), .A2(new_n703), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n799), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n800));
  XOR2_X1   g599(.A(KEYINPUT49), .B(G64gat), .Z(new_n801));
  OAI21_X1  g600(.A(new_n800), .B1(new_n799), .B2(new_n801), .ZN(G1333gat));
  NAND3_X1  g601(.A1(new_n795), .A2(G71gat), .A3(new_n771), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n795), .A2(new_n504), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n804), .B2(G71gat), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g605(.A1(new_n795), .A2(new_n718), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g607(.A1(new_n672), .A2(new_n746), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n543), .A2(new_n793), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n812), .A2(KEYINPUT117), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n743), .A2(KEYINPUT51), .A3(new_n809), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n812), .A2(KEYINPUT117), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n458), .A2(G85gat), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n813), .A2(new_n692), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n672), .A2(new_n746), .A3(new_n693), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n744), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n700), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n817), .B1(new_n821), .B2(new_n598), .ZN(G1336gat));
  NAND2_X1  g621(.A1(new_n813), .A2(new_n815), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n792), .A2(new_n599), .A3(new_n703), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n744), .A2(new_n703), .A3(new_n818), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n826), .B1(new_n828), .B2(new_n599), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n824), .B1(new_n812), .B2(new_n814), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n830), .B1(G92gat), .B2(new_n827), .ZN(new_n831));
  OAI22_X1  g630(.A1(new_n825), .A2(new_n829), .B1(new_n826), .B2(new_n831), .ZN(G1337gat));
  NOR2_X1   g631(.A1(new_n503), .A2(G99gat), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n813), .A2(new_n692), .A3(new_n815), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n771), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n834), .B1(new_n836), .B2(new_n377), .ZN(G1338gat));
  NOR3_X1   g636(.A1(new_n745), .A2(G106gat), .A3(new_n282), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n813), .A2(new_n815), .A3(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n744), .A2(new_n784), .A3(new_n818), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(G106gat), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n839), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n734), .B1(new_n543), .B2(new_n793), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n735), .B1(new_n739), .B2(new_n742), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n718), .B(new_n818), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(G106gat), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n810), .A2(new_n811), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT51), .B1(new_n743), .B2(new_n809), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n838), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT118), .B1(new_n851), .B2(KEYINPUT53), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n853));
  AOI211_X1 g652(.A(new_n853), .B(new_n840), .C1(new_n847), .C2(new_n850), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n843), .B1(new_n852), .B2(new_n854), .ZN(G1339gat));
  INV_X1    g654(.A(new_n746), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n694), .A2(KEYINPUT119), .A3(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n629), .A2(new_n672), .A3(new_n693), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(new_n859), .B2(new_n746), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT55), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n679), .A2(new_n674), .A3(new_n680), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(KEYINPUT54), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(new_n681), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n679), .A2(new_n680), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n867), .A3(new_n683), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n687), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n862), .B1(new_n865), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n688), .B1(new_n681), .B2(new_n867), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n871), .B(KEYINPUT55), .C1(new_n681), .C2(new_n864), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n870), .A2(new_n689), .A3(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n588), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n574), .A2(new_n576), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n876), .B(KEYINPUT120), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n579), .A2(new_n580), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n879), .A2(KEYINPUT121), .A3(new_n591), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT121), .B1(new_n879), .B2(new_n591), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n728), .A2(new_n727), .A3(new_n729), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n874), .B(new_n882), .C1(new_n883), .C2(new_n730), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n879), .A2(new_n591), .ZN(new_n885));
  OAI22_X1  g684(.A1(new_n873), .A2(new_n856), .B1(new_n693), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n731), .A2(new_n886), .A3(new_n732), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n861), .B1(new_n888), .B2(new_n672), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n541), .A3(new_n504), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n703), .A2(new_n458), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n595), .ZN(new_n895));
  OAI21_X1  g694(.A(G113gat), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n889), .A2(new_n397), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(new_n892), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n342), .A3(new_n746), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n896), .A2(new_n899), .ZN(G1340gat));
  OAI21_X1  g699(.A(G120gat), .B1(new_n894), .B2(new_n745), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n898), .A2(new_n340), .A3(new_n692), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1341gat));
  NAND3_X1  g702(.A1(new_n893), .A2(G127gat), .A3(new_n672), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n904), .A2(KEYINPUT122), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n904), .A2(KEYINPUT122), .ZN(new_n906));
  AOI21_X1  g705(.A(G127gat), .B1(new_n898), .B2(new_n672), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(G1342gat));
  OAI21_X1  g707(.A(G134gat), .B1(new_n894), .B2(new_n629), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n703), .A2(G134gat), .A3(new_n629), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n889), .A2(new_n700), .A3(new_n397), .A4(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(KEYINPUT56), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n911), .A2(KEYINPUT56), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n909), .A2(new_n912), .A3(new_n913), .ZN(G1343gat));
  INV_X1    g713(.A(KEYINPUT57), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n889), .A2(new_n915), .A3(new_n784), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n873), .A2(new_n593), .A3(new_n594), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n885), .A2(new_n693), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n629), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n672), .B1(new_n884), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n857), .A2(new_n860), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n718), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT57), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n891), .A2(new_n539), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n916), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n226), .B1(new_n926), .B2(new_n595), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n672), .B1(new_n884), .B2(new_n887), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n784), .B1(new_n928), .B2(new_n921), .ZN(new_n929));
  NOR4_X1   g728(.A1(new_n929), .A2(new_n924), .A3(G141gat), .A4(new_n895), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n930), .A2(KEYINPUT58), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n916), .A2(new_n923), .A3(new_n746), .A4(new_n925), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n930), .B1(new_n932), .B2(G141gat), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT58), .ZN(new_n934));
  OAI22_X1  g733(.A1(new_n927), .A2(new_n931), .B1(new_n933), .B2(new_n934), .ZN(G1344gat));
  AOI211_X1 g734(.A(KEYINPUT59), .B(new_n402), .C1(new_n926), .C2(new_n692), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT59), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n874), .A2(new_n793), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(KEYINPUT123), .B1(new_n629), .B2(new_n873), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n939), .A2(new_n940), .A3(new_n882), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n941), .A2(new_n919), .ZN(new_n942));
  OAI22_X1  g741(.A1(new_n942), .A2(new_n672), .B1(new_n595), .B2(new_n859), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n541), .A2(KEYINPUT57), .ZN(new_n944));
  AOI22_X1  g743(.A1(new_n943), .A2(new_n944), .B1(new_n929), .B2(KEYINPUT57), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(new_n692), .A3(new_n925), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n937), .B1(new_n946), .B2(G148gat), .ZN(new_n947));
  INV_X1    g746(.A(new_n929), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(new_n925), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n692), .A2(new_n402), .ZN(new_n950));
  OAI22_X1  g749(.A1(new_n936), .A2(new_n947), .B1(new_n949), .B2(new_n950), .ZN(G1345gat));
  NOR2_X1   g750(.A1(new_n747), .A2(new_n234), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n948), .A2(new_n672), .A3(new_n925), .ZN(new_n953));
  AOI22_X1  g752(.A1(new_n926), .A2(new_n952), .B1(new_n234), .B2(new_n953), .ZN(G1346gat));
  AOI21_X1  g753(.A(new_n235), .B1(new_n926), .B2(new_n733), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n700), .A2(new_n235), .A3(new_n502), .A4(new_n793), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n929), .A2(new_n771), .A3(new_n956), .ZN(new_n957));
  OR2_X1    g756(.A1(new_n955), .A2(new_n957), .ZN(G1347gat));
  NOR2_X1   g757(.A1(new_n700), .A2(new_n502), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  NOR4_X1   g759(.A1(new_n890), .A2(new_n285), .A3(new_n895), .A4(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n897), .A2(new_n856), .A3(new_n960), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n962), .B(KEYINPUT124), .C1(G169gat), .C2(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT124), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n963), .A2(G169gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n965), .B1(new_n966), .B2(new_n961), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n964), .A2(new_n967), .ZN(G1348gat));
  NOR2_X1   g767(.A1(new_n897), .A2(new_n960), .ZN(new_n969));
  AOI21_X1  g768(.A(G176gat), .B1(new_n969), .B2(new_n692), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n890), .A2(new_n960), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n745), .A2(new_n286), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(G1349gat));
  NAND3_X1  g772(.A1(new_n969), .A2(new_n299), .A3(new_n672), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n890), .A2(new_n747), .A3(new_n960), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n974), .B1(new_n975), .B2(new_n654), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(KEYINPUT60), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT60), .ZN(new_n978));
  OAI211_X1 g777(.A(new_n974), .B(new_n978), .C1(new_n654), .C2(new_n975), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(new_n979), .ZN(G1350gat));
  NAND3_X1  g779(.A1(new_n969), .A2(new_n303), .A3(new_n733), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT61), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n971), .A2(new_n793), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n982), .B1(new_n983), .B2(G190gat), .ZN(new_n984));
  AOI211_X1 g783(.A(KEYINPUT61), .B(new_n303), .C1(new_n971), .C2(new_n793), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n981), .B1(new_n984), .B2(new_n985), .ZN(G1351gat));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n987), .B1(new_n959), .B2(new_n539), .ZN(new_n988));
  NOR3_X1   g787(.A1(new_n960), .A2(KEYINPUT126), .A3(new_n771), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n945), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g789(.A(G197gat), .B1(new_n990), .B2(new_n895), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n539), .A2(new_n703), .A3(new_n784), .ZN(new_n992));
  XOR2_X1   g791(.A(new_n992), .B(KEYINPUT125), .Z(new_n993));
  NAND3_X1  g792(.A1(new_n993), .A2(new_n458), .A3(new_n889), .ZN(new_n994));
  INV_X1    g793(.A(new_n994), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n995), .A2(new_n585), .A3(new_n746), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n991), .A2(new_n996), .ZN(G1352gat));
  NOR3_X1   g796(.A1(new_n994), .A2(G204gat), .A3(new_n693), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT62), .ZN(new_n999));
  OR2_X1    g798(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g799(.A(G204gat), .B1(new_n990), .B2(new_n745), .ZN(new_n1001));
  INV_X1    g800(.A(KEYINPUT127), .ZN(new_n1002));
  AND3_X1   g801(.A1(new_n998), .A2(new_n1002), .A3(new_n999), .ZN(new_n1003));
  AOI21_X1  g802(.A(new_n1002), .B1(new_n998), .B2(new_n999), .ZN(new_n1004));
  OAI211_X1 g803(.A(new_n1000), .B(new_n1001), .C1(new_n1003), .C2(new_n1004), .ZN(G1353gat));
  NAND3_X1  g804(.A1(new_n995), .A2(new_n202), .A3(new_n672), .ZN(new_n1006));
  OAI211_X1 g805(.A(new_n945), .B(new_n672), .C1(new_n988), .C2(new_n989), .ZN(new_n1007));
  AND3_X1   g806(.A1(new_n1007), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1008));
  AOI21_X1  g807(.A(KEYINPUT63), .B1(new_n1007), .B2(G211gat), .ZN(new_n1009));
  OAI21_X1  g808(.A(new_n1006), .B1(new_n1008), .B2(new_n1009), .ZN(G1354gat));
  OAI21_X1  g809(.A(G218gat), .B1(new_n990), .B2(new_n629), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n995), .A2(new_n203), .A3(new_n733), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1011), .A2(new_n1012), .ZN(G1355gat));
endmodule


