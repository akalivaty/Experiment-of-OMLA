//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  AND3_X1   g0012(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n213));
  AOI21_X1  g0013(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n214));
  OAI21_X1  g0014(.A(G20), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT66), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT65), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n209), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n212), .B1(new_n215), .B2(new_n216), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XOR2_X1   g0026(.A(G250), .B(G257), .Z(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT67), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G264), .B(G270), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n230), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G87), .B(G97), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT68), .ZN(new_n237));
  XOR2_X1   g0037(.A(G107), .B(G116), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT69), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n202), .A2(G68), .ZN(new_n241));
  INV_X1    g0041(.A(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n240), .B(new_n246), .ZN(G351));
  NAND2_X1  g0047(.A1(G33), .A2(G41), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n248), .B1(new_n213), .B2(new_n214), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G223), .ZN(new_n251));
  AND2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  OAI21_X1  g0055(.A(KEYINPUT71), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OR2_X1    g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT71), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(new_n260), .A3(G1698), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n251), .B1(new_n256), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(G1698), .B1(new_n257), .B2(new_n258), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G222), .ZN(new_n264));
  INV_X1    g0064(.A(G77), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n264), .B1(new_n265), .B2(new_n259), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n250), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G41), .ZN(new_n268));
  INV_X1    g0068(.A(G45), .ZN(new_n269));
  AOI21_X1  g0069(.A(G1), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n248), .A2(G1), .A3(G13), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(new_n271), .A3(G274), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n274));
  AOI21_X1  g0074(.A(KEYINPUT70), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n271), .A2(KEYINPUT70), .A3(new_n274), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n273), .B1(new_n278), .B2(G226), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n267), .A2(G190), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n267), .A2(new_n279), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G200), .ZN(new_n282));
  INV_X1    g0082(.A(G58), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT8), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT8), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G58), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G33), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(G20), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n287), .A2(new_n289), .B1(G150), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n203), .A2(G20), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G1), .A2(G13), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT64), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n297));
  NAND3_X1  g0097(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G13), .ZN(new_n300));
  NOR3_X1   g0100(.A1(new_n300), .A2(new_n207), .A3(G1), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n293), .A2(new_n299), .B1(new_n202), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT9), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n299), .A2(new_n301), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n206), .A2(G20), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n304), .A2(G50), .A3(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n302), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n303), .B1(new_n302), .B2(new_n306), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n280), .B(new_n282), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT10), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT75), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT74), .B1(new_n308), .B2(new_n309), .ZN(new_n313));
  INV_X1    g0113(.A(new_n309), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT74), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n314), .A2(new_n315), .A3(new_n307), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT10), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n282), .A2(new_n318), .A3(new_n280), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n312), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n317), .A2(new_n319), .A3(new_n312), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n311), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n302), .A2(new_n306), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G169), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(new_n281), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(G179), .B2(new_n281), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT16), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n257), .A2(new_n207), .A3(new_n258), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT7), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n257), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n258), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n242), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n283), .A2(new_n242), .ZN(new_n335));
  OAI21_X1  g0135(.A(G20), .B1(new_n335), .B2(new_n201), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n290), .A2(G159), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n329), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT7), .B1(new_n254), .B2(new_n207), .ZN(new_n340));
  NOR4_X1   g0140(.A1(new_n252), .A2(new_n253), .A3(new_n331), .A4(G20), .ZN(new_n341));
  OAI21_X1  g0141(.A(G68), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n338), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(KEYINPUT16), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n339), .A2(new_n344), .A3(new_n299), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n287), .A2(new_n305), .ZN(new_n346));
  INV_X1    g0146(.A(new_n287), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n304), .A2(new_n346), .B1(new_n301), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT81), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT18), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n345), .A2(KEYINPUT81), .A3(new_n348), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n251), .A2(new_n255), .ZN(new_n354));
  INV_X1    g0154(.A(G226), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G1698), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n354), .B(new_n356), .C1(new_n252), .C2(new_n253), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G33), .A2(G87), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n250), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n271), .A2(G232), .A3(new_n274), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n272), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G179), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n360), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n249), .B1(new_n358), .B2(new_n357), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n272), .A2(new_n361), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n364), .B(KEYINPUT82), .C1(new_n367), .C2(G169), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT82), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(new_n369), .A3(new_n363), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n351), .A2(new_n352), .A3(new_n353), .A4(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G200), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(new_n360), .B2(new_n362), .ZN(new_n374));
  INV_X1    g0174(.A(G190), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n365), .A2(new_n366), .A3(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n345), .A2(new_n377), .A3(new_n348), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT17), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n345), .A2(new_n377), .A3(KEYINPUT17), .A4(new_n348), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n351), .A2(new_n353), .A3(new_n371), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n382), .B1(KEYINPUT18), .B2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n323), .A2(new_n328), .A3(new_n372), .A4(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G33), .A2(G97), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT76), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT76), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n388), .A2(G33), .A3(G97), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(G226), .A2(G1698), .ZN(new_n391));
  INV_X1    g0191(.A(G232), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n391), .B1(new_n392), .B2(G1698), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n390), .B1(new_n259), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n272), .B1(new_n394), .B2(new_n249), .ZN(new_n395));
  INV_X1    g0195(.A(G238), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n276), .B2(new_n277), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT13), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT77), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n387), .A2(new_n389), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n355), .A2(new_n255), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n392), .A2(G1698), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n401), .B(new_n402), .C1(new_n252), .C2(new_n253), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n273), .B1(new_n404), .B2(new_n250), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT13), .ZN(new_n406));
  INV_X1    g0206(.A(new_n277), .ZN(new_n407));
  OAI21_X1  g0207(.A(G238), .B1(new_n407), .B2(new_n275), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n405), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n398), .A2(new_n399), .A3(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n405), .A2(new_n408), .A3(KEYINPUT77), .A4(new_n406), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(G169), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT14), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n413), .A2(KEYINPUT80), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n410), .A2(G169), .A3(new_n411), .A4(new_n414), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n398), .A2(new_n409), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n419), .A2(new_n363), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n301), .A2(new_n242), .ZN(new_n423));
  XNOR2_X1  g0223(.A(new_n423), .B(KEYINPUT12), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n304), .A2(G68), .A3(new_n305), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT79), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n290), .A2(G50), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT78), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n289), .A2(G77), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(new_n207), .B2(G68), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n299), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT11), .ZN(new_n434));
  OR2_X1    g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n424), .A2(new_n425), .A3(KEYINPUT79), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n433), .A2(new_n434), .ZN(new_n437));
  AND4_X1   g0237(.A1(new_n428), .A2(new_n435), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n422), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n410), .A2(G200), .A3(new_n411), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n438), .B(new_n441), .C1(new_n419), .C2(new_n375), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n396), .B1(new_n256), .B2(new_n261), .ZN(new_n443));
  INV_X1    g0243(.A(new_n263), .ZN(new_n444));
  INV_X1    g0244(.A(G107), .ZN(new_n445));
  OAI22_X1  g0245(.A1(new_n444), .A2(new_n392), .B1(new_n445), .B2(new_n259), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n250), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n273), .B1(new_n278), .B2(G244), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n363), .ZN(new_n451));
  XNOR2_X1  g0251(.A(KEYINPUT15), .B(G87), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n289), .ZN(new_n454));
  INV_X1    g0254(.A(new_n290), .ZN(new_n455));
  OAI221_X1 g0255(.A(new_n454), .B1(new_n207), .B2(new_n265), .C1(new_n455), .C2(new_n347), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n456), .A2(new_n299), .B1(new_n265), .B2(new_n301), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n304), .A2(G77), .A3(new_n305), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n449), .A2(new_n326), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n451), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n373), .B1(new_n447), .B2(new_n448), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT73), .ZN(new_n463));
  OR3_X1    g0263(.A1(new_n459), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n450), .A2(KEYINPUT72), .A3(G190), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n463), .B1(new_n459), .B2(new_n462), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT72), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n449), .B2(new_n375), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n464), .A2(new_n465), .A3(new_n466), .A4(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n440), .A2(new_n442), .A3(new_n461), .A4(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n385), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n206), .A2(G33), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n304), .A2(G116), .A3(new_n472), .ZN(new_n473));
  OR2_X1    g0273(.A1(KEYINPUT85), .A2(G116), .ZN(new_n474));
  NAND2_X1  g0274(.A1(KEYINPUT85), .A2(G116), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n301), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n474), .A2(G20), .A3(new_n475), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G283), .ZN(new_n480));
  INV_X1    g0280(.A(G97), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n480), .B(new_n207), .C1(G33), .C2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n299), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT20), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n483), .A2(new_n484), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n473), .B(new_n478), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n259), .A2(G264), .A3(G1698), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n259), .A2(G257), .A3(new_n255), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n254), .A2(G303), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n250), .ZN(new_n492));
  XNOR2_X1  g0292(.A(KEYINPUT5), .B(G41), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n206), .A2(G45), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n271), .A2(G274), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT86), .ZN(new_n500));
  INV_X1    g0300(.A(new_n271), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n501), .B1(new_n495), .B2(new_n493), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n500), .B1(new_n502), .B2(G270), .ZN(new_n503));
  AND4_X1   g0303(.A1(new_n500), .A2(new_n496), .A3(G270), .A4(new_n271), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n492), .B(new_n499), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n505), .A2(KEYINPUT21), .A3(G169), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n505), .A2(new_n363), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n487), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n487), .B1(new_n505), .B2(G200), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n375), .B2(new_n505), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n505), .A2(new_n487), .A3(G169), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT87), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT21), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n512), .B1(new_n511), .B2(new_n513), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n508), .B(new_n510), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n207), .B(G87), .C1(new_n252), .C2(new_n253), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT22), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT22), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n259), .A2(new_n520), .A3(new_n207), .A4(G87), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n288), .B1(new_n474), .B2(new_n475), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT23), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(new_n207), .B2(G107), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n445), .A2(KEYINPUT23), .A3(G20), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n523), .A2(new_n207), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(KEYINPUT24), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT24), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n530), .B1(new_n522), .B2(new_n527), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n299), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n259), .A2(G257), .A3(G1698), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G294), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT88), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n263), .A2(new_n537), .A3(G250), .ZN(new_n538));
  OAI211_X1 g0338(.A(G250), .B(new_n255), .C1(new_n252), .C2(new_n253), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT88), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n250), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n498), .B1(G264), .B2(new_n502), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(G190), .A3(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n544), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n249), .B1(new_n536), .B2(new_n541), .ZN(new_n547));
  OAI21_X1  g0347(.A(G200), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT25), .ZN(new_n549));
  INV_X1    g0349(.A(new_n301), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n550), .B2(G107), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n301), .A2(KEYINPUT25), .A3(new_n445), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n304), .A2(new_n472), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n553), .B1(new_n554), .B2(new_n445), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n532), .A2(new_n545), .A3(new_n548), .A4(new_n556), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n532), .A2(new_n556), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n543), .A2(new_n363), .A3(new_n544), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n546), .A2(new_n547), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n559), .B1(new_n560), .B2(G169), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n557), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n301), .A2(new_n481), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n554), .B2(new_n481), .ZN(new_n564));
  OAI21_X1  g0364(.A(G107), .B1(new_n340), .B2(new_n341), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n290), .A2(G77), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT83), .ZN(new_n567));
  XNOR2_X1  g0367(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT6), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n569), .A2(new_n481), .A3(G107), .ZN(new_n570));
  XNOR2_X1  g0370(.A(G97), .B(G107), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n570), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n565), .B(new_n568), .C1(new_n207), .C2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n564), .B1(new_n573), .B2(new_n299), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n496), .A2(G257), .A3(new_n271), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n263), .A2(KEYINPUT4), .A3(G244), .ZN(new_n576));
  OAI211_X1 g0376(.A(G244), .B(new_n255), .C1(new_n252), .C2(new_n253), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT4), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n259), .A2(G250), .A3(G1698), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n576), .A2(new_n579), .A3(new_n480), .A4(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n575), .B1(new_n581), .B2(new_n250), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n582), .A2(G190), .A3(new_n499), .ZN(new_n583));
  AOI211_X1 g0383(.A(new_n498), .B(new_n575), .C1(new_n581), .C2(new_n250), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n574), .B(new_n583), .C1(new_n373), .C2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n564), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n568), .B1(new_n207), .B2(new_n572), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n445), .B1(new_n332), .B2(new_n333), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n299), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n582), .A2(new_n363), .A3(new_n499), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n590), .B(new_n591), .C1(G169), .C2(new_n584), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n585), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT19), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n207), .B1(new_n400), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(G87), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n596), .A2(new_n481), .A3(new_n445), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(KEYINPUT19), .B1(new_n289), .B2(G97), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n254), .A2(G20), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n599), .B1(new_n600), .B2(G68), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n213), .A2(new_n214), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n598), .A2(new_n601), .B1(new_n602), .B2(new_n298), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n452), .A2(new_n301), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n554), .A2(new_n452), .ZN(new_n606));
  NOR3_X1   g0406(.A1(new_n603), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n259), .A2(G244), .A3(G1698), .ZN(new_n608));
  INV_X1    g0408(.A(new_n523), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n608), .B(new_n609), .C1(new_n444), .C2(new_n396), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n250), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT84), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n494), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n206), .A2(KEYINPUT84), .A3(G45), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n613), .A2(G250), .A3(new_n271), .A4(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n497), .B2(new_n494), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n326), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n616), .B1(new_n610), .B2(new_n250), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n363), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n598), .A2(new_n601), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n299), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n611), .A2(G190), .A3(new_n617), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n554), .A2(new_n596), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n624), .A2(new_n625), .A3(new_n604), .A4(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n620), .A2(new_n373), .ZN(new_n629));
  OAI22_X1  g0429(.A1(new_n607), .A2(new_n622), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n562), .A2(new_n593), .A3(new_n630), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n471), .A2(new_n517), .A3(new_n631), .ZN(G372));
  INV_X1    g0432(.A(new_n328), .ZN(new_n633));
  OR3_X1    g0433(.A1(new_n317), .A2(new_n312), .A3(new_n319), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n634), .A2(new_n320), .B1(KEYINPUT10), .B2(new_n310), .ZN(new_n635));
  INV_X1    g0435(.A(new_n382), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n420), .B1(new_n416), .B2(new_n417), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n637), .A2(new_n438), .ZN(new_n638));
  INV_X1    g0438(.A(new_n461), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n639), .A2(new_n442), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n636), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n349), .A2(new_n371), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT18), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n349), .A2(new_n371), .A3(new_n352), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT90), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n635), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n641), .A2(KEYINPUT90), .A3(new_n645), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n633), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n471), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT26), .B1(new_n630), .B2(new_n592), .ZN(new_n652));
  INV_X1    g0452(.A(new_n592), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n624), .A2(new_n604), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n619), .B(new_n621), .C1(new_n655), .C2(new_n606), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n603), .A2(new_n605), .A3(new_n626), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n618), .A2(KEYINPUT89), .A3(G200), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT89), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n620), .B2(new_n373), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n657), .A2(new_n625), .A3(new_n658), .A4(new_n660), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n653), .A2(new_n654), .A3(new_n656), .A4(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n652), .A2(new_n662), .A3(new_n656), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n532), .A2(new_n556), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n664), .B(new_n559), .C1(G169), .C2(new_n560), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n665), .B(new_n508), .C1(new_n514), .C2(new_n515), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n658), .A2(new_n660), .ZN(new_n667));
  OAI22_X1  g0467(.A1(new_n667), .A2(new_n628), .B1(new_n622), .B2(new_n607), .ZN(new_n668));
  INV_X1    g0468(.A(new_n557), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n593), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n663), .B1(new_n666), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n650), .B1(new_n651), .B2(new_n671), .ZN(G369));
  OR2_X1    g0472(.A1(new_n514), .A2(new_n515), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n508), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT91), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n674), .A2(new_n487), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n487), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n517), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT92), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT92), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n683), .A2(new_n688), .A3(new_n685), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(G330), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n682), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n558), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT93), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n562), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(KEYINPUT93), .B1(new_n558), .B2(new_n693), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(KEYINPUT94), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(KEYINPUT94), .B1(new_n696), .B2(new_n697), .ZN(new_n700));
  OAI22_X1  g0500(.A1(new_n699), .A2(new_n700), .B1(new_n665), .B2(new_n693), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n692), .A2(new_n701), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n665), .A2(new_n682), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n696), .A2(new_n697), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT94), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n682), .B1(new_n673), .B2(new_n508), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(new_n698), .A3(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n702), .A2(new_n703), .A3(new_n708), .ZN(G399));
  NAND2_X1  g0509(.A1(new_n210), .A2(new_n268), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n597), .A2(G116), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(G1), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n216), .B2(new_n710), .ZN(new_n713));
  XOR2_X1   g0513(.A(new_n713), .B(KEYINPUT28), .Z(new_n714));
  INV_X1    g0514(.A(KEYINPUT95), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n652), .A2(new_n662), .A3(new_n656), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n670), .A2(new_n666), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n682), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n715), .B1(new_n718), .B2(KEYINPUT29), .ZN(new_n719));
  OAI21_X1  g0519(.A(KEYINPUT26), .B1(new_n668), .B2(new_n592), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n656), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n630), .A2(KEYINPUT26), .A3(new_n592), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n682), .B1(new_n723), .B2(new_n717), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT29), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT29), .ZN(new_n726));
  OAI211_X1 g0526(.A(KEYINPUT95), .B(new_n726), .C1(new_n671), .C2(new_n682), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n719), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n631), .A2(new_n517), .A3(new_n693), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n503), .A2(new_n504), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n731), .A2(G179), .A3(new_n492), .A4(new_n499), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n543), .A2(new_n582), .A3(new_n620), .A4(new_n544), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n730), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n582), .A2(new_n620), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n507), .A2(new_n735), .A3(KEYINPUT30), .A4(new_n560), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n543), .A2(new_n544), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n582), .A2(new_n499), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n620), .A2(G179), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n737), .A2(new_n738), .A3(new_n739), .A4(new_n505), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n734), .A2(new_n736), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n682), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT31), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n741), .A2(KEYINPUT31), .A3(new_n682), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n729), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G330), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n728), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n714), .B1(new_n748), .B2(new_n206), .ZN(new_n749));
  XOR2_X1   g0549(.A(new_n749), .B(KEYINPUT96), .Z(G364));
  INV_X1    g0550(.A(new_n690), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G330), .ZN(new_n752));
  INV_X1    g0552(.A(new_n710), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n300), .A2(G20), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n206), .B1(new_n754), .B2(G45), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n690), .A2(new_n691), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n752), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n602), .B1(G20), .B2(new_n326), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n210), .A2(new_n259), .ZN(new_n767));
  INV_X1    g0567(.A(G355), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n767), .A2(new_n768), .B1(G116), .B2(new_n210), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n210), .A2(new_n254), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT97), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n216), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n772), .B1(new_n269), .B2(new_n773), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n246), .A2(new_n269), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n769), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n375), .A2(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(new_n363), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G97), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT100), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n207), .A2(new_n363), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G200), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n781), .B1(new_n783), .B2(G190), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n783), .A2(new_n781), .A3(G190), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n780), .B1(new_n787), .B2(new_n242), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT101), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n783), .A2(new_n375), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n254), .B1(new_n790), .B2(G50), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n782), .B(KEYINPUT98), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G190), .A2(G200), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n792), .A2(new_n777), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n791), .B1(new_n794), .B2(new_n265), .C1(new_n283), .C2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n207), .A2(G179), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n797), .A2(new_n375), .A3(G200), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n445), .ZN(new_n799));
  XOR2_X1   g0599(.A(KEYINPUT99), .B(G159), .Z(new_n800));
  NAND2_X1  g0600(.A1(new_n797), .A2(new_n793), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT32), .Z(new_n803));
  NAND3_X1  g0603(.A1(new_n797), .A2(G190), .A3(G200), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n596), .ZN(new_n805));
  NOR4_X1   g0605(.A1(new_n796), .A2(new_n799), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n801), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n259), .B1(new_n807), .B2(G329), .ZN(new_n808));
  INV_X1    g0608(.A(G294), .ZN(new_n809));
  INV_X1    g0609(.A(new_n779), .ZN(new_n810));
  INV_X1    g0610(.A(G322), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n808), .B1(new_n809), .B2(new_n810), .C1(new_n795), .C2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n794), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n812), .B1(G311), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n790), .ZN(new_n815));
  INV_X1    g0615(.A(G326), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G283), .ZN(new_n818));
  INV_X1    g0618(.A(G303), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n818), .A2(new_n798), .B1(new_n804), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n787), .ZN(new_n821));
  XNOR2_X1  g0621(.A(KEYINPUT33), .B(G317), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n817), .B(new_n820), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n789), .A2(new_n806), .B1(new_n814), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n761), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n757), .B1(new_n766), .B2(new_n776), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT102), .Z(new_n827));
  INV_X1    g0627(.A(new_n764), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n827), .B1(new_n751), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n760), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(G396));
  NAND2_X1  g0631(.A1(new_n682), .A2(new_n459), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n639), .B1(new_n469), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n461), .A2(new_n682), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n718), .B(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n757), .B1(new_n836), .B2(new_n747), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n747), .B2(new_n836), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n761), .A2(new_n762), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n758), .B1(new_n839), .B2(new_n265), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n259), .B1(new_n807), .B2(G311), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n780), .B(new_n841), .C1(new_n795), .C2(new_n809), .ZN(new_n842));
  INV_X1    g0642(.A(new_n798), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n790), .A2(G303), .B1(new_n843), .B2(G87), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n844), .B1(new_n445), .B2(new_n804), .C1(new_n787), .C2(new_n818), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n842), .B(new_n845), .C1(new_n476), .C2(new_n813), .ZN(new_n846));
  INV_X1    g0646(.A(new_n795), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n847), .A2(G143), .B1(G137), .B2(new_n790), .ZN(new_n848));
  INV_X1    g0648(.A(G150), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n848), .B1(new_n849), .B2(new_n787), .C1(new_n794), .C2(new_n800), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT34), .ZN(new_n851));
  INV_X1    g0651(.A(G132), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n259), .B1(new_n801), .B2(new_n852), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n810), .A2(new_n283), .B1(new_n804), .B2(new_n202), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n853), .B(new_n854), .C1(G68), .C2(new_n843), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n846), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n840), .B1(new_n856), .B2(new_n825), .C1(new_n835), .C2(new_n763), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n838), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(G384));
  AND3_X1   g0659(.A1(new_n345), .A2(KEYINPUT106), .A3(new_n348), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT106), .B1(new_n345), .B2(new_n348), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n371), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n680), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n860), .B2(new_n861), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n862), .A2(new_n864), .A3(new_n378), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT37), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT37), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n378), .A2(new_n867), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n345), .A2(KEYINPUT81), .A3(new_n348), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT81), .B1(new_n345), .B2(new_n348), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n868), .B1(new_n871), .B2(new_n371), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n351), .A2(new_n353), .A3(new_n863), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n866), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n383), .A2(KEYINPUT18), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(new_n372), .A3(new_n636), .ZN(new_n877));
  INV_X1    g0677(.A(new_n864), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n875), .A2(new_n879), .A3(KEYINPUT38), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n643), .A2(new_n380), .A3(new_n381), .A4(new_n644), .ZN(new_n881));
  INV_X1    g0681(.A(new_n873), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n868), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n383), .A2(new_n873), .A3(new_n884), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n642), .A2(new_n378), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n867), .B1(new_n886), .B2(new_n873), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n883), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT38), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n880), .A2(new_n890), .A3(KEYINPUT109), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT109), .B1(new_n880), .B2(new_n890), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT108), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n742), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n741), .A2(KEYINPUT108), .A3(new_n682), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n895), .A2(new_n743), .A3(new_n896), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n897), .A2(new_n745), .A3(new_n729), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n418), .A2(new_n421), .A3(new_n442), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n693), .A2(new_n438), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n900), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n442), .B(new_n902), .C1(new_n637), .C2(new_n438), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n901), .A2(new_n903), .A3(KEYINPUT105), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT105), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n440), .A2(new_n905), .A3(new_n442), .A4(new_n902), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n904), .A2(new_n906), .A3(new_n835), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT40), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n898), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n904), .A2(new_n835), .A3(new_n906), .ZN(new_n910));
  AOI22_X1  g0710(.A1(KEYINPUT37), .A2(new_n865), .B1(new_n872), .B2(new_n873), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n864), .B1(new_n384), .B2(new_n372), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n889), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n880), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n897), .A2(new_n745), .A3(new_n729), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n910), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  XOR2_X1   g0716(.A(KEYINPUT107), .B(KEYINPUT40), .Z(new_n917));
  AOI22_X1  g0717(.A1(new_n893), .A2(new_n909), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n471), .A2(new_n915), .ZN(new_n920));
  OAI21_X1  g0720(.A(G330), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n920), .B2(new_n919), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n880), .A2(new_n890), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT39), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n924), .B2(new_n914), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n440), .A2(new_n682), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n718), .A2(new_n835), .ZN(new_n930));
  INV_X1    g0730(.A(new_n834), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n904), .A2(new_n906), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n932), .A2(new_n914), .A3(new_n934), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n645), .A2(new_n863), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n929), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n471), .A2(new_n719), .A3(new_n725), .A4(new_n727), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n650), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n938), .B(new_n940), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n922), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n922), .A2(new_n941), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n942), .B(new_n943), .C1(new_n206), .C2(new_n754), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n241), .A2(KEYINPUT103), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n241), .A2(KEYINPUT103), .ZN(new_n946));
  OAI21_X1  g0746(.A(G77), .B1(new_n283), .B2(new_n242), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n945), .B(new_n946), .C1(new_n216), .C2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n948), .A2(G1), .A3(new_n300), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT104), .Z(new_n950));
  INV_X1    g0750(.A(G116), .ZN(new_n951));
  INV_X1    g0751(.A(new_n572), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n951), .B(new_n215), .C1(new_n952), .C2(KEYINPUT35), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(KEYINPUT35), .B2(new_n952), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT36), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n950), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(new_n955), .B2(new_n954), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n944), .A2(new_n957), .ZN(G367));
  NAND2_X1  g0758(.A1(new_n653), .A2(new_n682), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n585), .B(new_n592), .C1(new_n693), .C2(new_n574), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  OR3_X1    g0762(.A1(new_n702), .A2(KEYINPUT110), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n682), .B1(new_n655), .B2(new_n626), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n964), .A2(new_n661), .A3(new_n656), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n656), .B2(new_n964), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n967));
  OAI21_X1  g0767(.A(KEYINPUT110), .B1(new_n702), .B2(new_n962), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n963), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n708), .A2(new_n962), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n592), .B1(new_n960), .B2(new_n665), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n971), .A2(KEYINPUT42), .B1(new_n693), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(KEYINPUT42), .B2(new_n971), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n967), .B1(new_n963), .B2(new_n968), .ZN(new_n977));
  OR3_X1    g0777(.A1(new_n970), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n976), .B1(new_n970), .B2(new_n977), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n710), .B(KEYINPUT41), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n708), .B1(new_n701), .B2(new_n707), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n692), .B(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n748), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(KEYINPUT111), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT111), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n982), .A2(new_n986), .A3(new_n983), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n708), .A2(new_n703), .A3(new_n961), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT45), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n988), .A2(new_n989), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n708), .A2(new_n703), .ZN(new_n992));
  AND4_X1   g0792(.A1(KEYINPUT44), .A2(new_n992), .A3(new_n960), .A4(new_n959), .ZN(new_n993));
  AOI21_X1  g0793(.A(KEYINPUT44), .B1(new_n992), .B2(new_n962), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n702), .B1(new_n990), .B2(new_n991), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n993), .A2(new_n994), .B1(new_n990), .B2(new_n991), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n996), .A2(new_n692), .A3(new_n701), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n985), .A2(new_n987), .A3(new_n995), .A4(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n980), .B1(new_n998), .B2(new_n983), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n978), .B(new_n979), .C1(new_n999), .C2(new_n756), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n772), .A2(new_n230), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n765), .B1(new_n210), .B2(new_n452), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n757), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G283), .A2(new_n813), .B1(new_n847), .B2(G303), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT46), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n477), .B2(new_n804), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n798), .A2(new_n481), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n259), .B(new_n1007), .C1(G317), .C2(new_n807), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1004), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  NOR3_X1   g0809(.A1(new_n804), .A2(new_n1005), .A3(new_n951), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G107), .B2(new_n779), .ZN(new_n1011));
  INV_X1    g0811(.A(G311), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1011), .B1(new_n1012), .B2(new_n815), .C1(new_n787), .C2(new_n809), .ZN(new_n1013));
  INV_X1    g0813(.A(G137), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n259), .B1(new_n801), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(G143), .B2(new_n790), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n794), .B2(new_n202), .C1(new_n849), .C2(new_n795), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n804), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n1018), .A2(G58), .B1(new_n843), .B2(G77), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n242), .B2(new_n810), .C1(new_n787), .C2(new_n800), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n1009), .A2(new_n1013), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT47), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1003), .B1(new_n1022), .B2(new_n761), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n828), .B2(new_n966), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1000), .A2(new_n1024), .ZN(G387));
  NAND2_X1  g0825(.A1(new_n982), .A2(new_n756), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT112), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n234), .A2(new_n269), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n287), .A2(new_n202), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT50), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n711), .B(new_n269), .C1(new_n242), .C2(new_n265), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n771), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT113), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1028), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n1033), .B2(new_n1032), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(G107), .B2(new_n210), .C1(new_n711), .C2(new_n767), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n758), .B1(new_n1036), .B2(new_n765), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n779), .A2(new_n453), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n790), .A2(G159), .B1(new_n1018), .B2(G77), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(new_n787), .C2(new_n347), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(KEYINPUT114), .B(G150), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n254), .B(new_n1007), .C1(new_n807), .C2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n202), .B2(new_n795), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1040), .B(new_n1043), .C1(G68), .C2(new_n813), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n813), .A2(G303), .B1(G322), .B2(new_n790), .ZN(new_n1045));
  INV_X1    g0845(.A(G317), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1045), .B1(new_n1012), .B2(new_n787), .C1(new_n1046), .C2(new_n795), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT48), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G294), .A2(new_n1018), .B1(new_n779), .B2(G283), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1053), .A2(KEYINPUT49), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n254), .B1(new_n801), .B2(new_n816), .C1(new_n477), .C2(new_n798), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n1053), .B2(KEYINPUT49), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1044), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1037), .B1(new_n1057), .B2(new_n825), .C1(new_n701), .C2(new_n828), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n1027), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n710), .B1(new_n982), .B2(new_n983), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1060), .A2(KEYINPUT115), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n984), .A2(KEYINPUT115), .A3(new_n753), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(new_n983), .C2(new_n982), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1059), .A2(new_n1063), .ZN(G393));
  NAND2_X1  g0864(.A1(new_n997), .A2(new_n995), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1065), .A2(new_n755), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n962), .A2(new_n764), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n772), .A2(new_n239), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n765), .B1(new_n481), .B2(new_n210), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n757), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n254), .B1(new_n801), .B2(new_n811), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n799), .B(new_n1071), .C1(G283), .C2(new_n1018), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT117), .Z(new_n1073));
  OAI22_X1  g0873(.A1(new_n795), .A2(new_n1012), .B1(new_n1046), .B2(new_n815), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT52), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n794), .A2(new_n809), .B1(new_n477), .B2(new_n810), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(G303), .B2(new_n821), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1073), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(G159), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n795), .A2(new_n1079), .B1(new_n849), .B2(new_n815), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT51), .Z(new_n1081));
  NAND2_X1  g0881(.A1(new_n779), .A2(G77), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n347), .B2(new_n794), .C1(new_n787), .C2(new_n202), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n254), .B1(new_n807), .B2(G143), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1085), .B1(new_n242), .B2(new_n804), .C1(new_n596), .C2(new_n798), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT116), .Z(new_n1087));
  OAI21_X1  g0887(.A(new_n1078), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1070), .B1(new_n1088), .B2(new_n761), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1066), .B1(new_n1067), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1065), .A2(new_n984), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n998), .A2(new_n1091), .A3(new_n753), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1090), .A2(new_n1092), .ZN(G390));
  AOI21_X1  g0893(.A(new_n758), .B1(new_n839), .B2(new_n347), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n259), .B(new_n805), .C1(G294), .C2(new_n807), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n481), .B2(new_n794), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(G116), .B2(new_n847), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n1082), .B1(new_n242), .B2(new_n798), .C1(new_n815), .C2(new_n818), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(G107), .B2(new_n821), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(KEYINPUT54), .B(G143), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n852), .A2(new_n795), .B1(new_n794), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n254), .B1(new_n807), .B2(G125), .ZN(new_n1102));
  INV_X1    g0902(.A(G128), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1102), .B1(new_n815), .B2(new_n1103), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n810), .A2(new_n1079), .B1(new_n798), .B2(new_n202), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n1101), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1018), .A2(new_n1041), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT53), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(G137), .B2(new_n821), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1097), .A2(new_n1099), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1094), .B1(new_n1110), .B2(new_n825), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n926), .B2(new_n762), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n834), .B1(new_n718), .B2(new_n835), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n928), .B1(new_n1113), .B2(new_n933), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n926), .A2(new_n1114), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n682), .B(new_n833), .C1(new_n723), .C2(new_n717), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n934), .B1(new_n1116), .B2(new_n834), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n893), .A2(new_n1117), .A3(new_n928), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n910), .A2(G330), .A3(new_n746), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1115), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n833), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n724), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n931), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n927), .B1(new_n1123), .B2(new_n934), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1124), .A2(new_n893), .B1(new_n926), .B2(new_n1114), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n898), .A2(new_n691), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n910), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1120), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT120), .ZN(new_n1129));
  OR3_X1    g0929(.A1(new_n1128), .A2(new_n1129), .A3(new_n755), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1129), .B1(new_n1128), .B2(new_n755), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1112), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1126), .A2(new_n471), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n939), .A2(new_n1133), .A3(new_n650), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT118), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n746), .A2(G330), .A3(new_n835), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n1126), .A2(new_n910), .B1(new_n933), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n934), .B1(new_n1126), .B2(new_n835), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1122), .B(new_n931), .C1(new_n747), .C2(new_n907), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n1138), .A2(new_n1113), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n939), .A2(new_n1133), .A3(new_n650), .A4(KEYINPUT118), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1136), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  OR2_X1    g0943(.A1(new_n1128), .A2(new_n1143), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1128), .A2(new_n1143), .A3(KEYINPUT119), .ZN(new_n1145));
  AOI21_X1  g0945(.A(KEYINPUT119), .B1(new_n1128), .B2(new_n1143), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n753), .B(new_n1144), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1132), .A2(new_n1147), .ZN(G378));
  OR2_X1    g0948(.A1(new_n929), .A2(new_n937), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n325), .A2(new_n680), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n635), .B2(new_n633), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1150), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n323), .A2(new_n328), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1151), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n918), .B2(G330), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n898), .A2(new_n907), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT109), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n923), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n880), .A2(new_n890), .A3(KEYINPUT109), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1161), .A2(new_n1163), .A3(KEYINPUT40), .A4(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n914), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n915), .A2(new_n835), .A3(new_n904), .A4(new_n906), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n917), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  AND4_X1   g0968(.A1(G330), .A2(new_n1165), .A3(new_n1168), .A4(new_n1159), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1149), .B1(new_n1160), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1165), .A2(new_n1168), .A3(G330), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1159), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n918), .A2(G330), .A3(new_n1159), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1173), .A2(new_n1174), .A3(new_n938), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1170), .A2(KEYINPUT123), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1136), .A2(new_n1142), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1141), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1178), .B1(new_n1128), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT123), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1149), .B(new_n1181), .C1(new_n1160), .C2(new_n1169), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1176), .A2(new_n1180), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT57), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1184), .B1(new_n1170), .B2(new_n1175), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n710), .B1(new_n1186), .B2(new_n1180), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1176), .A2(new_n756), .A3(new_n1182), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n268), .B(new_n254), .C1(new_n801), .C2(new_n818), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n810), .A2(new_n242), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1190), .B(new_n1191), .C1(new_n813), .C2(new_n453), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n445), .B2(new_n795), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n787), .A2(new_n481), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n798), .A2(new_n283), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n815), .A2(new_n951), .B1(new_n265), .B2(new_n804), .ZN(new_n1196));
  NOR4_X1   g0996(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1201));
  AOI21_X1  g1001(.A(G50), .B1(new_n288), .B2(new_n268), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n259), .B2(G41), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n790), .A2(G125), .B1(new_n779), .B2(G150), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n804), .B2(new_n1100), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n1103), .A2(new_n795), .B1(new_n794), .B2(new_n1014), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(G132), .C2(new_n821), .ZN(new_n1208));
  XOR2_X1   g1008(.A(new_n1208), .B(KEYINPUT122), .Z(new_n1209));
  OR2_X1    g1009(.A1(new_n1209), .A2(KEYINPUT59), .ZN(new_n1210));
  AOI211_X1 g1010(.A(G33), .B(G41), .C1(new_n807), .C2(G124), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n798), .B2(new_n800), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n1209), .B2(KEYINPUT59), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1200), .B(new_n1204), .C1(new_n1210), .C2(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1214), .A2(new_n825), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n758), .B(new_n1215), .C1(new_n202), .C2(new_n839), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1172), .A2(new_n762), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1189), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1188), .A2(new_n1219), .ZN(G375));
  NAND2_X1  g1020(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n980), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1221), .A2(new_n1222), .A3(new_n1143), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n758), .B1(new_n839), .B2(new_n242), .ZN(new_n1224));
  OR2_X1    g1024(.A1(new_n787), .A2(new_n1100), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT124), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n1195), .B2(new_n254), .ZN(new_n1227));
  OAI211_X1 g1027(.A(KEYINPUT124), .B(new_n259), .C1(new_n798), .C2(new_n283), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1225), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n1014), .A2(new_n795), .B1(new_n794), .B2(new_n849), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n804), .A2(new_n1079), .B1(new_n801), .B2(new_n1103), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n815), .A2(new_n852), .B1(new_n810), .B2(new_n202), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n259), .B1(new_n807), .B2(G303), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1234), .B1(new_n265), .B2(new_n798), .C1(new_n795), .C2(new_n818), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G107), .B2(new_n813), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1038), .B1(new_n481), .B2(new_n804), .C1(new_n815), .C2(new_n809), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n476), .B2(new_n821), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1229), .A2(new_n1233), .B1(new_n1236), .B2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1224), .B1(new_n1239), .B2(new_n825), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(new_n933), .B2(new_n762), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1141), .B2(new_n756), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1223), .A2(new_n1242), .ZN(G381));
  NAND3_X1  g1043(.A1(new_n1059), .A2(new_n1063), .A3(new_n830), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(G390), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1245), .A2(new_n1246), .A3(new_n858), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n1247), .A2(G387), .A3(G381), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1248), .B(KEYINPUT125), .ZN(new_n1249));
  INV_X1    g1049(.A(G378), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1250), .A2(new_n1188), .A3(new_n1219), .ZN(new_n1251));
  OR2_X1    g1051(.A1(new_n1249), .A2(new_n1251), .ZN(G407));
  OAI211_X1 g1052(.A(G407), .B(G213), .C1(G343), .C2(new_n1251), .ZN(G409));
  NAND3_X1  g1053(.A1(new_n1000), .A2(new_n1024), .A3(G390), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(G390), .B1(new_n1000), .B2(new_n1024), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n830), .B1(new_n1059), .B2(new_n1063), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n1255), .A2(new_n1256), .B1(new_n1245), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1256), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1245), .A2(new_n1257), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(new_n1260), .A3(new_n1254), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT61), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1143), .A2(KEYINPUT60), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1264), .A2(new_n1221), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n753), .B1(new_n1264), .B2(new_n1221), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1242), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  OR2_X1    g1067(.A1(new_n1267), .A2(new_n858), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n858), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n681), .A2(G213), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(G2897), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n1268), .A2(new_n1269), .A3(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1272), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n1183), .A2(new_n980), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n755), .B1(new_n1170), .B2(new_n1175), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(new_n1217), .B2(new_n1216), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G378), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1188), .A2(G378), .A3(new_n1219), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT126), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1188), .A2(G378), .A3(KEYINPUT126), .A4(new_n1219), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1279), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1275), .B1(new_n1284), .B2(new_n1271), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1284), .A2(new_n1271), .A3(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT62), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1263), .B(new_n1285), .C1(new_n1287), .C2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1279), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n1270), .ZN(new_n1293));
  NOR3_X1   g1093(.A1(new_n1293), .A2(KEYINPUT62), .A3(new_n1286), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1262), .B1(new_n1289), .B2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT63), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(new_n1293), .B2(new_n1286), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT61), .B1(new_n1293), .B2(new_n1275), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1262), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1287), .A2(KEYINPUT63), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1297), .A2(new_n1298), .A3(new_n1299), .A4(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1295), .A2(new_n1301), .ZN(G405));
  NAND2_X1  g1102(.A1(G375), .A2(new_n1250), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1290), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1299), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1262), .A2(new_n1290), .A3(new_n1303), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1268), .A2(KEYINPUT127), .A3(new_n1269), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1308), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1305), .A2(new_n1310), .A3(new_n1306), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1309), .A2(new_n1311), .ZN(G402));
endmodule


