//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n585, new_n586, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n637,
    new_n638, new_n639, new_n642, new_n644, new_n645, new_n646, new_n648,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206, new_n1207;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n454), .A2(new_n458), .B1(new_n459), .B2(new_n455), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(new_n469), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n468), .B(new_n471), .C1(new_n472), .C2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NAND2_X1  g055(.A1(new_n476), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n465), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n477), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND2_X1  g064(.A1(KEYINPUT4), .A2(G138), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(new_n474), .B2(new_n475), .ZN(new_n491));
  NAND2_X1  g066(.A1(G102), .A2(G2104), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n477), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G126), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n474), .B2(new_n475), .ZN(new_n496));
  NAND2_X1  g071(.A1(G114), .A2(G2104), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(G2105), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  OAI211_X1 g074(.A(G138), .B(new_n477), .C1(new_n463), .C2(new_n464), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n494), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT66), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n494), .A2(new_n499), .A3(KEYINPUT66), .A4(new_n502), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G62), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n515), .A2(KEYINPUT67), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT67), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n514), .A2(new_n517), .A3(G62), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n509), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  OR2_X1    g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n511), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G50), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n520), .A2(new_n521), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(new_n514), .ZN(new_n525));
  INV_X1    g100(.A(G88), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n519), .A2(new_n527), .ZN(G166));
  AND2_X1   g103(.A1(new_n524), .A2(new_n514), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G89), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT70), .B(KEYINPUT7), .ZN(new_n531));
  AND3_X1   g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n522), .A2(G51), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n530), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT68), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n514), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n512), .A2(KEYINPUT68), .A3(new_n513), .ZN(new_n538));
  AND2_X1   g113(.A1(G63), .A2(G651), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT69), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n537), .A2(KEYINPUT69), .A3(new_n538), .A4(new_n539), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n535), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(G168));
  NAND2_X1  g121(.A1(new_n522), .A2(G52), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n525), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(G77), .A2(G543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n537), .A2(new_n538), .ZN(new_n551));
  INV_X1    g126(.A(G64), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n549), .B1(new_n553), .B2(G651), .ZN(G171));
  NAND2_X1  g129(.A1(new_n522), .A2(G43), .ZN(new_n555));
  INV_X1    g130(.A(G81), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n525), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT71), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g134(.A(new_n555), .B(KEYINPUT71), .C1(new_n525), .C2(new_n556), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n562));
  NAND2_X1  g137(.A1(G68), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G56), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n551), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G651), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n561), .A2(new_n562), .A3(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n562), .B1(new_n561), .B2(new_n566), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G860), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT73), .ZN(G153));
  NAND4_X1  g147(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g148(.A1(G1), .A2(G3), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT8), .ZN(new_n575));
  NAND4_X1  g150(.A1(G319), .A2(G483), .A3(G661), .A4(new_n575), .ZN(G188));
  NAND2_X1  g151(.A1(new_n522), .A2(G53), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT9), .ZN(new_n578));
  XNOR2_X1  g153(.A(KEYINPUT74), .B(G65), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n514), .A2(new_n579), .B1(G78), .B2(G543), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(new_n509), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n529), .A2(G91), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n578), .A2(new_n581), .A3(new_n582), .ZN(G299));
  INV_X1    g158(.A(G171), .ZN(G301));
  AND3_X1   g159(.A1(new_n535), .A2(KEYINPUT75), .A3(new_n544), .ZN(new_n585));
  AOI21_X1  g160(.A(KEYINPUT75), .B1(new_n535), .B2(new_n544), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(G286));
  INV_X1    g162(.A(G166), .ZN(G303));
  AOI21_X1  g163(.A(G74), .B1(new_n537), .B2(new_n538), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(new_n509), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n522), .A2(G49), .ZN(new_n591));
  INV_X1    g166(.A(G87), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n525), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G288));
  INV_X1    g170(.A(G61), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n596), .B1(new_n512), .B2(new_n513), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT76), .ZN(new_n598));
  INV_X1    g173(.A(G73), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n597), .A2(new_n598), .B1(new_n599), .B2(new_n511), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n514), .A2(new_n598), .A3(G61), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(G651), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n522), .A2(G48), .ZN(new_n604));
  INV_X1    g179(.A(G86), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n525), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(G305));
  NAND3_X1  g183(.A1(new_n537), .A2(G60), .A3(new_n538), .ZN(new_n609));
  NAND2_X1  g184(.A1(G72), .A2(G543), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n509), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n522), .A2(G47), .ZN(new_n612));
  XNOR2_X1  g187(.A(KEYINPUT77), .B(G85), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n525), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(G290));
  NAND2_X1  g191(.A1(G301), .A2(G868), .ZN(new_n617));
  INV_X1    g192(.A(G54), .ZN(new_n618));
  INV_X1    g193(.A(new_n522), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(KEYINPUT78), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(KEYINPUT78), .B2(new_n619), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n529), .A2(KEYINPUT10), .A3(G92), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT10), .ZN(new_n623));
  INV_X1    g198(.A(G92), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n525), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g201(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n514), .A2(G66), .ZN(new_n628));
  INV_X1    g203(.A(G79), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(new_n511), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n509), .B1(new_n630), .B2(KEYINPUT79), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(KEYINPUT79), .B2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n617), .B1(new_n634), .B2(G868), .ZN(G284));
  OAI21_X1  g210(.A(new_n617), .B1(new_n634), .B2(G868), .ZN(G321));
  INV_X1    g211(.A(G299), .ZN(new_n637));
  OAI21_X1  g212(.A(KEYINPUT80), .B1(new_n637), .B2(G868), .ZN(new_n638));
  NAND2_X1  g213(.A1(G286), .A2(G868), .ZN(new_n639));
  MUX2_X1   g214(.A(KEYINPUT80), .B(new_n638), .S(new_n639), .Z(G297));
  XOR2_X1   g215(.A(G297), .B(KEYINPUT81), .Z(G280));
  INV_X1    g216(.A(G559), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n634), .B1(new_n642), .B2(G860), .ZN(G148));
  NOR2_X1   g218(.A1(new_n633), .A2(G559), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(G868), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(G868), .B2(new_n570), .ZN(G323));
  XOR2_X1   g222(.A(KEYINPUT82), .B(KEYINPUT11), .Z(new_n648));
  XNOR2_X1  g223(.A(G323), .B(new_n648), .ZN(G282));
  NAND2_X1  g224(.A1(new_n476), .A2(new_n470), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT12), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT13), .ZN(new_n652));
  INV_X1    g227(.A(G2100), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  AOI22_X1  g230(.A1(new_n482), .A2(G123), .B1(new_n484), .B2(G135), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n477), .A2(G111), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n469), .B1(new_n657), .B2(KEYINPUT83), .ZN(new_n658));
  OAI21_X1  g233(.A(KEYINPUT83), .B1(G99), .B2(G2105), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n658), .B1(new_n657), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(G2096), .Z(new_n663));
  NAND3_X1  g238(.A1(new_n654), .A2(new_n655), .A3(new_n663), .ZN(G156));
  INV_X1    g239(.A(G14), .ZN(new_n665));
  XOR2_X1   g240(.A(KEYINPUT15), .B(G2435), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2438), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2427), .B(G2430), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT85), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n669), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(KEYINPUT14), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT86), .ZN(new_n673));
  XOR2_X1   g248(.A(G1341), .B(G1348), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2451), .B(G2454), .Z(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2443), .B(G2446), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n665), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(new_n680), .B2(new_n679), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(G401));
  XOR2_X1   g258(.A(G2084), .B(G2090), .Z(new_n684));
  XNOR2_X1  g259(.A(G2067), .B(G2678), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT87), .ZN(new_n686));
  NOR2_X1   g261(.A1(G2072), .A2(G2078), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n444), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n684), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n688), .B(KEYINPUT17), .Z(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(new_n686), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n688), .A2(new_n685), .A3(new_n684), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT18), .Z(new_n694));
  NAND3_X1  g269(.A1(new_n691), .A2(new_n686), .A3(new_n684), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n692), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(new_n653), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT88), .B(G2096), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(G227));
  XOR2_X1   g274(.A(G1971), .B(G1976), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT19), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1956), .B(G2474), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1961), .B(G1966), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT20), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n702), .A2(new_n703), .ZN(new_n707));
  NOR3_X1   g282(.A1(new_n701), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n701), .B2(new_n707), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT89), .Z(new_n711));
  XOR2_X1   g286(.A(G1981), .B(G1986), .Z(new_n712));
  XNOR2_X1  g287(.A(G1991), .B(G1996), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n711), .B(new_n716), .ZN(G229));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G20), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT23), .Z(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G299), .B2(G16), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT95), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G1956), .ZN(new_n724));
  INV_X1    g299(.A(G2090), .ZN(new_n725));
  INV_X1    g300(.A(G29), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G35), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT94), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G162), .B2(new_n726), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT29), .Z(new_n730));
  OAI22_X1  g305(.A1(new_n723), .A2(new_n724), .B1(new_n725), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n724), .B2(new_n723), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT96), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n726), .A2(G26), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT28), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n482), .A2(G128), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n484), .A2(G140), .ZN(new_n737));
  OR2_X1    g312(.A1(G104), .A2(G2105), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n738), .B(G2104), .C1(G116), .C2(new_n477), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n736), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n735), .B1(new_n741), .B2(new_n726), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT91), .ZN(new_n743));
  INV_X1    g318(.A(G2067), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n718), .A2(G4), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n634), .B2(new_n718), .ZN(new_n747));
  INV_X1    g322(.A(G1348), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(G27), .A2(G29), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G164), .B2(G29), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(new_n443), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n745), .A2(new_n749), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT30), .B(G28), .ZN(new_n754));
  OR2_X1    g329(.A1(KEYINPUT31), .A2(G11), .ZN(new_n755));
  NAND2_X1  g330(.A1(KEYINPUT31), .A2(G11), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n754), .A2(new_n726), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n662), .B2(new_n726), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT93), .Z(new_n759));
  INV_X1    g334(.A(KEYINPUT24), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(G34), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n726), .B1(new_n760), .B2(G34), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n762), .B2(KEYINPUT92), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(KEYINPUT92), .B2(new_n762), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G160), .B2(G29), .ZN(new_n765));
  INV_X1    g340(.A(G2084), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n759), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n726), .A2(G33), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n477), .A2(G103), .A3(G2104), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT25), .Z(new_n771));
  INV_X1    g346(.A(G139), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n478), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(G115), .A2(G2104), .ZN(new_n774));
  INV_X1    g349(.A(G127), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n465), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n773), .B1(G2105), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n769), .B1(new_n777), .B2(new_n726), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G2072), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n726), .A2(G32), .ZN(new_n780));
  NAND3_X1  g355(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT26), .Z(new_n782));
  INV_X1    g357(.A(G129), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n481), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n470), .A2(G105), .ZN(new_n785));
  INV_X1    g360(.A(G141), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n478), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n780), .B1(new_n788), .B2(new_n726), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT27), .B(G1996), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n789), .B(new_n790), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n718), .A2(G5), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G171), .B2(new_n718), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1961), .ZN(new_n794));
  NOR4_X1   g369(.A1(new_n768), .A2(new_n779), .A3(new_n791), .A4(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(G168), .A2(new_n718), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n718), .B2(G21), .ZN(new_n797));
  INV_X1    g372(.A(G1966), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n725), .A2(new_n730), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n795), .B(new_n799), .C1(new_n798), .C2(new_n797), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n718), .A2(G19), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n570), .B2(new_n718), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1341), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n753), .A2(new_n800), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n733), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n718), .A2(G22), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G166), .B2(new_n718), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(G1971), .Z(new_n808));
  MUX2_X1   g383(.A(G6), .B(G305), .S(G16), .Z(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT32), .B(G1981), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT90), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n809), .B(new_n811), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n718), .A2(G23), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n594), .B2(new_n718), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT33), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n815), .A2(G1976), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n815), .A2(G1976), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n808), .B(new_n812), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(KEYINPUT34), .ZN(new_n819));
  OR2_X1    g394(.A1(G95), .A2(G2105), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n820), .B(G2104), .C1(G107), .C2(new_n477), .ZN(new_n821));
  INV_X1    g396(.A(G131), .ZN(new_n822));
  INV_X1    g397(.A(G119), .ZN(new_n823));
  OAI221_X1 g398(.A(new_n821), .B1(new_n478), .B2(new_n822), .C1(new_n823), .C2(new_n481), .ZN(new_n824));
  MUX2_X1   g399(.A(G25), .B(new_n824), .S(G29), .Z(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT35), .B(G1991), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n718), .A2(G24), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n615), .B2(new_n718), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n829), .A2(G1986), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n829), .A2(G1986), .ZN(new_n831));
  OR3_X1    g406(.A1(new_n827), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(new_n818), .B2(KEYINPUT34), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n819), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(KEYINPUT36), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n834), .A2(KEYINPUT36), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n805), .B1(new_n835), .B2(new_n836), .ZN(G311));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n835), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n838), .A2(new_n804), .A3(new_n733), .ZN(G150));
  NAND3_X1  g414(.A1(new_n537), .A2(G67), .A3(new_n538), .ZN(new_n840));
  NAND2_X1  g415(.A1(G80), .A2(G543), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n509), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n522), .A2(G55), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT97), .B(G93), .Z(new_n844));
  OAI21_X1  g419(.A(new_n843), .B1(new_n525), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n568), .B2(new_n569), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n561), .A2(new_n566), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n849), .A2(new_n847), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT38), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n634), .A2(G559), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n856));
  AOI21_X1  g431(.A(G860), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n856), .B2(new_n855), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n847), .A2(G860), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT37), .Z(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(G145));
  NAND2_X1  g436(.A1(new_n503), .A2(KEYINPUT98), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT98), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n494), .A2(new_n499), .A3(new_n863), .A4(new_n502), .ZN(new_n864));
  AND2_X1   g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n741), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n777), .B(new_n788), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n824), .B(new_n651), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n482), .A2(G130), .ZN(new_n870));
  OAI21_X1  g445(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n871));
  INV_X1    g446(.A(G118), .ZN(new_n872));
  AOI22_X1  g447(.A1(new_n871), .A2(KEYINPUT99), .B1(new_n872), .B2(G2105), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(KEYINPUT99), .B2(new_n871), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n484), .A2(G142), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n870), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n869), .B(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n877), .A2(KEYINPUT100), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n868), .A2(new_n878), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n877), .A2(KEYINPUT100), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n868), .B1(new_n880), .B2(new_n878), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n662), .B(new_n479), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n488), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G37), .ZN(new_n886));
  INV_X1    g461(.A(new_n884), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n879), .A2(new_n881), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n885), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n889), .B(new_n890), .ZN(G395));
  XOR2_X1   g466(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n594), .B(KEYINPUT103), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(G305), .ZN(new_n895));
  XNOR2_X1  g470(.A(G166), .B(new_n615), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n852), .A2(new_n644), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n848), .A2(new_n645), .A3(new_n851), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n633), .A2(new_n637), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT41), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n627), .A2(G299), .A3(new_n632), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n627), .A2(KEYINPUT102), .A3(G299), .A4(new_n632), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n901), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n904), .B1(new_n908), .B2(KEYINPUT41), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n900), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n898), .A2(new_n899), .A3(new_n908), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n897), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n897), .B1(new_n911), .B2(new_n910), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n893), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n897), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n910), .A2(new_n911), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n918), .A2(new_n892), .A3(new_n912), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n915), .A2(new_n919), .A3(G868), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT105), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n915), .A2(new_n919), .A3(new_n922), .A4(G868), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n846), .A2(G868), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(new_n923), .A3(new_n924), .ZN(G295));
  NAND3_X1  g500(.A1(new_n921), .A2(new_n923), .A3(new_n924), .ZN(G331));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n927));
  OAI21_X1  g502(.A(G171), .B1(new_n585), .B2(new_n586), .ZN(new_n928));
  NAND2_X1  g503(.A1(G301), .A2(new_n545), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n849), .A2(KEYINPUT72), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n846), .B1(new_n931), .B2(new_n567), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n930), .B1(new_n932), .B2(new_n850), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n848), .A2(new_n851), .A3(new_n928), .A4(new_n929), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(new_n934), .A3(KEYINPUT106), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n852), .A2(new_n936), .A3(new_n930), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(new_n909), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n933), .A2(new_n934), .A3(new_n908), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n897), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n886), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n897), .B1(new_n938), .B2(new_n939), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n927), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n901), .A2(KEYINPUT41), .A3(new_n903), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(KEYINPUT107), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n908), .A2(new_n902), .ZN(new_n946));
  AOI22_X1  g521(.A1(new_n945), .A2(new_n946), .B1(new_n933), .B2(new_n934), .ZN(new_n947));
  INV_X1    g522(.A(new_n908), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n948), .B1(new_n935), .B2(new_n937), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n916), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n950), .A2(KEYINPUT43), .A3(new_n886), .A4(new_n940), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n943), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT44), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT43), .B1(new_n941), .B2(new_n942), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n950), .A2(new_n927), .A3(new_n886), .A4(new_n940), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n953), .A2(new_n958), .ZN(G397));
  INV_X1    g534(.A(KEYINPUT55), .ZN(new_n960));
  INV_X1    g535(.A(G8), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n960), .B1(G166), .B2(new_n961), .ZN(new_n962));
  OAI211_X1 g537(.A(KEYINPUT55), .B(G8), .C1(new_n519), .C2(new_n527), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G1384), .ZN(new_n965));
  OAI211_X1 g540(.A(KEYINPUT4), .B(G138), .C1(new_n463), .C2(new_n464), .ZN(new_n966));
  AOI21_X1  g541(.A(G2105), .B1(new_n966), .B2(new_n492), .ZN(new_n967));
  OAI21_X1  g542(.A(G126), .B1(new_n463), .B2(new_n464), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n477), .B1(new_n968), .B2(new_n497), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT66), .B1(new_n970), .B2(new_n502), .ZN(new_n971));
  INV_X1    g546(.A(new_n506), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n965), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT50), .ZN(new_n974));
  INV_X1    g549(.A(G40), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n479), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n503), .A2(KEYINPUT111), .A3(new_n965), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT111), .B1(new_n503), .B2(new_n965), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n974), .A2(new_n725), .A3(new_n976), .A4(new_n980), .ZN(new_n981));
  XOR2_X1   g556(.A(KEYINPUT108), .B(G1384), .Z(new_n982));
  NAND4_X1  g557(.A1(new_n862), .A2(KEYINPUT45), .A3(new_n864), .A4(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(G1384), .B1(new_n505), .B2(new_n506), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n976), .B(new_n983), .C1(new_n984), .C2(KEYINPUT45), .ZN(new_n985));
  XNOR2_X1  g560(.A(KEYINPUT110), .B(G1971), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n961), .B1(new_n981), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT116), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n964), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  AOI211_X1 g565(.A(KEYINPUT116), .B(new_n961), .C1(new_n981), .C2(new_n987), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT49), .ZN(new_n993));
  INV_X1    g568(.A(new_n513), .ZN(new_n994));
  NOR2_X1   g569(.A1(KEYINPUT5), .A2(G543), .ZN(new_n995));
  OAI21_X1  g570(.A(G61), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n996), .A2(KEYINPUT76), .B1(G73), .B2(G543), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n509), .B1(new_n997), .B2(new_n601), .ZN(new_n998));
  OAI21_X1  g573(.A(G1981), .B1(new_n998), .B2(new_n606), .ZN(new_n999));
  INV_X1    g574(.A(G1981), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n603), .A2(new_n607), .A3(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n999), .A2(new_n1001), .A3(KEYINPUT113), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n1003));
  NAND3_X1  g578(.A1(G305), .A2(new_n1003), .A3(G1981), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n993), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1005), .B(KEYINPUT115), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n976), .B1(new_n978), .B2(new_n979), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT112), .B(G8), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1002), .A2(new_n993), .A3(new_n1004), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1002), .A2(KEYINPUT114), .A3(new_n993), .A4(new_n1004), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1010), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1006), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n503), .A2(new_n965), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT45), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n503), .A2(KEYINPUT111), .A3(new_n965), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n965), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n1023), .A3(new_n976), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n798), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n974), .A2(new_n766), .A3(new_n976), .A4(new_n980), .ZN(new_n1026));
  AOI211_X1 g601(.A(G286), .B(new_n1008), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n594), .A2(G1976), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1007), .A2(new_n1009), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(new_n594), .B2(G1976), .ZN(new_n1031));
  OR2_X1    g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1029), .A2(KEYINPUT52), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1016), .A2(new_n1027), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT63), .B1(new_n992), .B2(new_n1035), .ZN(new_n1036));
  AOI211_X1 g611(.A(new_n961), .B(new_n964), .C1(new_n981), .C2(new_n987), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1039), .B(new_n1009), .C1(new_n586), .C2(new_n585), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT63), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1019), .A2(KEYINPUT50), .A3(new_n1021), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n977), .B(new_n965), .C1(new_n971), .C2(new_n972), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1042), .A2(new_n1043), .A3(new_n725), .A4(new_n976), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1008), .B1(new_n987), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n964), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1041), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1038), .B1(new_n1040), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1049), .B1(new_n1006), .B2(new_n1015), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1010), .ZN(new_n1052));
  AOI211_X1 g627(.A(G1976), .B(G288), .C1(new_n1006), .C2(new_n1015), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1001), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n1036), .A2(new_n1051), .A3(new_n1055), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n976), .B(new_n744), .C1(new_n978), .C2(new_n979), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n980), .B(new_n976), .C1(new_n977), .C2(new_n984), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1058), .B1(new_n1059), .B2(new_n748), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT120), .B1(new_n1060), .B2(new_n633), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1042), .A2(new_n1043), .A3(new_n976), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT117), .B(G1956), .Z(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n973), .A2(new_n1020), .ZN(new_n1065));
  XOR2_X1   g640(.A(KEYINPUT56), .B(G2072), .Z(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1065), .A2(new_n976), .A3(new_n983), .A4(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1064), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT57), .ZN(new_n1071));
  XOR2_X1   g646(.A(new_n1071), .B(KEYINPUT119), .Z(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1070), .A2(KEYINPUT57), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1073), .B1(G299), .B2(new_n1074), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n581), .A2(new_n582), .ZN(new_n1076));
  OR2_X1    g651(.A1(new_n1070), .A2(KEYINPUT57), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1076), .A2(new_n578), .A3(new_n1077), .A4(new_n1072), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT121), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1075), .A2(new_n1078), .A3(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1069), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n1084));
  NAND2_X1  g659(.A1(G160), .A2(G40), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1085), .B1(new_n1086), .B2(new_n977), .ZN(new_n1087));
  AOI21_X1  g662(.A(G1348), .B1(new_n1087), .B2(new_n974), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1084), .B(new_n634), .C1(new_n1088), .C2(new_n1058), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1061), .A2(new_n1083), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1079), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1064), .A2(new_n1068), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT60), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1094), .B1(new_n1088), .B2(new_n1058), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1059), .A2(new_n748), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1096), .A2(KEYINPUT60), .A3(new_n1057), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(new_n634), .A3(new_n1097), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT58), .B(G1341), .Z(new_n1099));
  NAND2_X1  g674(.A1(new_n1007), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1100), .B1(new_n985), .B2(G1996), .ZN(new_n1101));
  AND2_X1   g676(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n568), .A2(new_n569), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT123), .B1(KEYINPUT122), .B2(KEYINPUT59), .ZN(new_n1105));
  XOR2_X1   g680(.A(new_n1105), .B(KEYINPUT124), .Z(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1106), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1101), .A2(new_n1103), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n985), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1111), .A2(new_n1067), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1092), .B(KEYINPUT61), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1098), .A2(new_n1110), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT61), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1064), .A2(new_n1068), .A3(new_n1091), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1091), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1060), .A2(KEYINPUT60), .A3(new_n633), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1093), .B1(new_n1115), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n980), .A2(new_n976), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n984), .A2(new_n977), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1123), .A2(G2084), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1085), .B1(new_n984), .B2(KEYINPUT45), .ZN(new_n1126));
  AOI21_X1  g701(.A(G1966), .B1(new_n1126), .B2(new_n1022), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n545), .B(new_n1009), .C1(new_n1125), .C2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(G168), .A2(new_n1008), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n961), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1128), .B(KEYINPUT51), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n987), .A2(new_n1044), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1046), .B1(new_n1132), .B2(new_n1009), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1037), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1039), .A2(new_n1009), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1129), .A2(KEYINPUT51), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AND4_X1   g712(.A1(new_n1131), .A2(new_n1134), .A3(new_n1137), .A4(new_n1050), .ZN(new_n1138));
  INV_X1    g713(.A(G1961), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1059), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT53), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(new_n985), .B2(G2078), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1126), .A2(KEYINPUT53), .A3(new_n443), .A4(new_n1022), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1140), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(G171), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n865), .A2(new_n982), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n1020), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1141), .A2(new_n975), .A3(G2078), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n471), .B1(new_n478), .B2(new_n472), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT125), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n468), .B(new_n1148), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1151), .B1(new_n1150), .B2(new_n1149), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1147), .A2(new_n983), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1140), .A2(new_n1153), .A3(new_n1142), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1145), .B1(G171), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n1144), .A2(G171), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1156), .B1(new_n1154), .B2(G171), .ZN(new_n1158));
  AOI22_X1  g733(.A1(new_n1155), .A2(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1122), .A2(new_n1138), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1128), .A2(KEYINPUT51), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1130), .A2(new_n1129), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1137), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1131), .A2(KEYINPUT62), .A3(new_n1137), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1134), .A2(new_n1050), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1145), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1056), .A2(new_n1160), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT109), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1146), .A2(new_n1020), .A3(new_n976), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(G1996), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1171), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1172), .A2(KEYINPUT109), .A3(G1996), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n788), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n740), .B(new_n744), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1178), .B1(new_n1174), .B2(new_n788), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1173), .A2(new_n1179), .ZN(new_n1180));
  XOR2_X1   g755(.A(new_n824), .B(new_n826), .Z(new_n1181));
  OAI211_X1 g756(.A(new_n1177), .B(new_n1180), .C1(new_n1172), .C2(new_n1181), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n615), .B(G1986), .Z(new_n1183));
  AOI21_X1  g758(.A(new_n1182), .B1(new_n1173), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1170), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n824), .A2(new_n826), .ZN(new_n1186));
  XOR2_X1   g761(.A(new_n1186), .B(KEYINPUT126), .Z(new_n1187));
  NAND3_X1  g762(.A1(new_n1177), .A2(new_n1180), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n741), .A2(new_n744), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1172), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NOR3_X1   g765(.A1(new_n1172), .A2(G1986), .A3(G290), .ZN(new_n1191));
  XOR2_X1   g766(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1192));
  XNOR2_X1  g767(.A(new_n1191), .B(new_n1192), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1182), .A2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1172), .B1(new_n788), .B2(new_n1178), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT46), .ZN(new_n1196));
  OR3_X1    g771(.A1(new_n1175), .A2(new_n1196), .A3(new_n1176), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1196), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1195), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT47), .ZN(new_n1200));
  OR2_X1    g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1202));
  AOI211_X1 g777(.A(new_n1190), .B(new_n1194), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1185), .A2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g779(.A1(G229), .A2(G227), .A3(new_n460), .ZN(new_n1206));
  NAND3_X1  g780(.A1(new_n682), .A2(new_n889), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g781(.A(new_n1207), .B1(new_n954), .B2(new_n955), .ZN(G308));
  NAND4_X1  g782(.A1(new_n956), .A2(new_n682), .A3(new_n889), .A4(new_n1206), .ZN(G225));
endmodule


