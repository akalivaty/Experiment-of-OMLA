

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582;

  XNOR2_X1 U325 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U326 ( .A(n373), .B(n372), .ZN(n374) );
  NOR2_X1 U327 ( .A1(n525), .A2(n446), .ZN(n560) );
  XNOR2_X1 U328 ( .A(n380), .B(n293), .ZN(n381) );
  XOR2_X1 U329 ( .A(G134GAT), .B(G106GAT), .Z(n293) );
  INV_X1 U330 ( .A(KEYINPUT11), .ZN(n372) );
  INV_X1 U331 ( .A(KEYINPUT48), .ZN(n412) );
  XNOR2_X1 U332 ( .A(n412), .B(KEYINPUT64), .ZN(n413) );
  XNOR2_X1 U333 ( .A(n414), .B(n413), .ZN(n522) );
  XNOR2_X1 U334 ( .A(n382), .B(n381), .ZN(n383) );
  INV_X1 U335 ( .A(G190GAT), .ZN(n447) );
  XOR2_X1 U336 ( .A(n424), .B(n313), .Z(n525) );
  XNOR2_X1 U337 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U338 ( .A(n450), .B(n449), .ZN(G1351GAT) );
  XNOR2_X1 U339 ( .A(KEYINPUT17), .B(KEYINPUT83), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n294), .B(G183GAT), .ZN(n295) );
  XOR2_X1 U341 ( .A(n295), .B(KEYINPUT18), .Z(n297) );
  XNOR2_X1 U342 ( .A(KEYINPUT82), .B(KEYINPUT19), .ZN(n296) );
  XOR2_X1 U343 ( .A(n297), .B(n296), .Z(n424) );
  XOR2_X1 U344 ( .A(G190GAT), .B(G99GAT), .Z(n299) );
  XNOR2_X1 U345 ( .A(G43GAT), .B(G15GAT), .ZN(n298) );
  XNOR2_X1 U346 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U347 ( .A(n300), .B(G176GAT), .Z(n302) );
  XOR2_X1 U348 ( .A(G120GAT), .B(G71GAT), .Z(n389) );
  XNOR2_X1 U349 ( .A(G169GAT), .B(n389), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U351 ( .A(KEYINPUT84), .B(KEYINPUT81), .Z(n304) );
  NAND2_X1 U352 ( .A1(G227GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U353 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U354 ( .A(n306), .B(n305), .Z(n312) );
  XNOR2_X1 U355 ( .A(G127GAT), .B(KEYINPUT79), .ZN(n307) );
  XNOR2_X1 U356 ( .A(n307), .B(KEYINPUT0), .ZN(n308) );
  XOR2_X1 U357 ( .A(n308), .B(KEYINPUT80), .Z(n310) );
  XNOR2_X1 U358 ( .A(G113GAT), .B(G134GAT), .ZN(n309) );
  XNOR2_X1 U359 ( .A(n310), .B(n309), .ZN(n439) );
  XNOR2_X1 U360 ( .A(n439), .B(KEYINPUT20), .ZN(n311) );
  XNOR2_X1 U361 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U362 ( .A(G141GAT), .B(G22GAT), .Z(n336) );
  XOR2_X1 U363 ( .A(KEYINPUT90), .B(KEYINPUT22), .Z(n315) );
  XNOR2_X1 U364 ( .A(KEYINPUT23), .B(G204GAT), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U366 ( .A(n336), .B(n316), .Z(n318) );
  NAND2_X1 U367 ( .A1(G228GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U369 ( .A(n319), .B(KEYINPUT85), .Z(n322) );
  XNOR2_X1 U370 ( .A(G50GAT), .B(KEYINPUT73), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n320), .B(G162GAT), .ZN(n375) );
  XNOR2_X1 U372 ( .A(n375), .B(KEYINPUT24), .ZN(n321) );
  XNOR2_X1 U373 ( .A(n322), .B(n321), .ZN(n325) );
  XOR2_X1 U374 ( .A(G155GAT), .B(KEYINPUT2), .Z(n324) );
  XNOR2_X1 U375 ( .A(KEYINPUT3), .B(KEYINPUT89), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n324), .B(n323), .ZN(n435) );
  XOR2_X1 U377 ( .A(n325), .B(n435), .Z(n333) );
  XOR2_X1 U378 ( .A(KEYINPUT86), .B(KEYINPUT21), .Z(n327) );
  XNOR2_X1 U379 ( .A(G218GAT), .B(KEYINPUT88), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U381 ( .A(n328), .B(KEYINPUT87), .Z(n330) );
  XNOR2_X1 U382 ( .A(G197GAT), .B(G211GAT), .ZN(n329) );
  XNOR2_X1 U383 ( .A(n330), .B(n329), .ZN(n420) );
  XNOR2_X1 U384 ( .A(G106GAT), .B(G78GAT), .ZN(n331) );
  XOR2_X1 U385 ( .A(n331), .B(G148GAT), .Z(n392) );
  XOR2_X1 U386 ( .A(n420), .B(n392), .Z(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n459) );
  XOR2_X1 U388 ( .A(G15GAT), .B(G1GAT), .Z(n359) );
  XOR2_X1 U389 ( .A(G169GAT), .B(G8GAT), .Z(n421) );
  XOR2_X1 U390 ( .A(n359), .B(n421), .Z(n335) );
  NAND2_X1 U391 ( .A1(G229GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n335), .B(n334), .ZN(n337) );
  XOR2_X1 U393 ( .A(n337), .B(n336), .Z(n345) );
  XOR2_X1 U394 ( .A(G197GAT), .B(G113GAT), .Z(n339) );
  XNOR2_X1 U395 ( .A(G36GAT), .B(G50GAT), .ZN(n338) );
  XNOR2_X1 U396 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U397 ( .A(KEYINPUT68), .B(KEYINPUT29), .Z(n341) );
  XNOR2_X1 U398 ( .A(KEYINPUT69), .B(KEYINPUT30), .ZN(n340) );
  XNOR2_X1 U399 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U400 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U402 ( .A(KEYINPUT8), .B(KEYINPUT70), .Z(n347) );
  XNOR2_X1 U403 ( .A(G43GAT), .B(G29GAT), .ZN(n346) );
  XNOR2_X1 U404 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U405 ( .A(KEYINPUT7), .B(n348), .ZN(n384) );
  XNOR2_X1 U406 ( .A(n349), .B(n384), .ZN(n568) );
  INV_X1 U407 ( .A(n568), .ZN(n539) );
  XNOR2_X1 U408 ( .A(KEYINPUT45), .B(KEYINPUT113), .ZN(n387) );
  XOR2_X1 U409 ( .A(G78GAT), .B(G71GAT), .Z(n351) );
  XNOR2_X1 U410 ( .A(G183GAT), .B(G127GAT), .ZN(n350) );
  XNOR2_X1 U411 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U412 ( .A(KEYINPUT12), .B(G155GAT), .Z(n353) );
  XNOR2_X1 U413 ( .A(G22GAT), .B(G211GAT), .ZN(n352) );
  XNOR2_X1 U414 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U415 ( .A(n355), .B(n354), .Z(n361) );
  XOR2_X1 U416 ( .A(G57GAT), .B(KEYINPUT13), .Z(n388) );
  XOR2_X1 U417 ( .A(G8GAT), .B(n388), .Z(n357) );
  NAND2_X1 U418 ( .A1(G231GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U419 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U421 ( .A(n361), .B(n360), .ZN(n369) );
  XOR2_X1 U422 ( .A(KEYINPUT76), .B(KEYINPUT78), .Z(n363) );
  XNOR2_X1 U423 ( .A(G64GAT), .B(KEYINPUT75), .ZN(n362) );
  XNOR2_X1 U424 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U425 ( .A(KEYINPUT77), .B(KEYINPUT15), .Z(n365) );
  XNOR2_X1 U426 ( .A(KEYINPUT74), .B(KEYINPUT14), .ZN(n364) );
  XNOR2_X1 U427 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U428 ( .A(n367), .B(n366), .Z(n368) );
  XNOR2_X1 U429 ( .A(n369), .B(n368), .ZN(n575) );
  XOR2_X1 U430 ( .A(G36GAT), .B(G190GAT), .Z(n418) );
  XOR2_X1 U431 ( .A(KEYINPUT65), .B(n418), .Z(n371) );
  XOR2_X1 U432 ( .A(G99GAT), .B(G85GAT), .Z(n396) );
  XNOR2_X1 U433 ( .A(G218GAT), .B(n396), .ZN(n370) );
  XNOR2_X1 U434 ( .A(n371), .B(n370), .ZN(n377) );
  NAND2_X1 U435 ( .A1(G232GAT), .A2(G233GAT), .ZN(n373) );
  XOR2_X1 U436 ( .A(n377), .B(n376), .Z(n382) );
  XOR2_X1 U437 ( .A(KEYINPUT9), .B(KEYINPUT66), .Z(n379) );
  XNOR2_X1 U438 ( .A(G92GAT), .B(KEYINPUT10), .ZN(n378) );
  XNOR2_X1 U439 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U440 ( .A(n384), .B(n383), .ZN(n534) );
  XOR2_X1 U441 ( .A(KEYINPUT36), .B(KEYINPUT101), .Z(n385) );
  XNOR2_X1 U442 ( .A(n534), .B(n385), .ZN(n578) );
  AND2_X1 U443 ( .A1(n575), .A2(n578), .ZN(n386) );
  XNOR2_X1 U444 ( .A(n387), .B(n386), .ZN(n403) );
  XNOR2_X1 U445 ( .A(n389), .B(n388), .ZN(n402) );
  XOR2_X1 U446 ( .A(G64GAT), .B(G92GAT), .Z(n391) );
  XNOR2_X1 U447 ( .A(G176GAT), .B(G204GAT), .ZN(n390) );
  XNOR2_X1 U448 ( .A(n391), .B(n390), .ZN(n415) );
  XNOR2_X1 U449 ( .A(n415), .B(n392), .ZN(n400) );
  XOR2_X1 U450 ( .A(KEYINPUT32), .B(KEYINPUT71), .Z(n394) );
  XNOR2_X1 U451 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U453 ( .A(n396), .B(n395), .Z(n398) );
  NAND2_X1 U454 ( .A1(G230GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U457 ( .A(n402), .B(n401), .ZN(n571) );
  NOR2_X1 U458 ( .A1(n403), .A2(n571), .ZN(n404) );
  NAND2_X1 U459 ( .A1(n539), .A2(n404), .ZN(n411) );
  XOR2_X1 U460 ( .A(KEYINPUT112), .B(KEYINPUT47), .Z(n409) );
  XNOR2_X1 U461 ( .A(KEYINPUT41), .B(n571), .ZN(n541) );
  NOR2_X1 U462 ( .A1(n541), .A2(n539), .ZN(n405) );
  XNOR2_X1 U463 ( .A(n405), .B(KEYINPUT46), .ZN(n406) );
  NOR2_X1 U464 ( .A1(n575), .A2(n406), .ZN(n407) );
  INV_X1 U465 ( .A(n534), .ZN(n550) );
  NAND2_X1 U466 ( .A1(n407), .A2(n550), .ZN(n408) );
  XNOR2_X1 U467 ( .A(n409), .B(n408), .ZN(n410) );
  NAND2_X1 U468 ( .A1(n411), .A2(n410), .ZN(n414) );
  XOR2_X1 U469 ( .A(KEYINPUT92), .B(n415), .Z(n417) );
  NAND2_X1 U470 ( .A1(G226GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U471 ( .A(n417), .B(n416), .ZN(n419) );
  XOR2_X1 U472 ( .A(n419), .B(n418), .Z(n423) );
  XNOR2_X1 U473 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U474 ( .A(n423), .B(n422), .ZN(n425) );
  XNOR2_X1 U475 ( .A(n425), .B(n424), .ZN(n513) );
  NOR2_X1 U476 ( .A1(n522), .A2(n513), .ZN(n426) );
  XNOR2_X1 U477 ( .A(KEYINPUT54), .B(n426), .ZN(n444) );
  XOR2_X1 U478 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n428) );
  XNOR2_X1 U479 ( .A(KEYINPUT4), .B(KEYINPUT91), .ZN(n427) );
  XNOR2_X1 U480 ( .A(n428), .B(n427), .ZN(n443) );
  XOR2_X1 U481 ( .A(G85GAT), .B(G162GAT), .Z(n430) );
  XNOR2_X1 U482 ( .A(G29GAT), .B(G120GAT), .ZN(n429) );
  XNOR2_X1 U483 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U484 ( .A(G57GAT), .B(G148GAT), .Z(n432) );
  XNOR2_X1 U485 ( .A(G141GAT), .B(G1GAT), .ZN(n431) );
  XNOR2_X1 U486 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U487 ( .A(n434), .B(n433), .Z(n441) );
  XOR2_X1 U488 ( .A(n435), .B(KEYINPUT1), .Z(n437) );
  NAND2_X1 U489 ( .A1(G225GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U490 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U491 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U492 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U493 ( .A(n443), .B(n442), .Z(n509) );
  NAND2_X1 U494 ( .A1(n444), .A2(n509), .ZN(n566) );
  NOR2_X1 U495 ( .A1(n459), .A2(n566), .ZN(n445) );
  XNOR2_X1 U496 ( .A(n445), .B(KEYINPUT55), .ZN(n446) );
  NAND2_X1 U497 ( .A1(n560), .A2(n534), .ZN(n450) );
  XOR2_X1 U498 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n448) );
  NOR2_X1 U499 ( .A1(n571), .A2(n539), .ZN(n451) );
  XNOR2_X1 U500 ( .A(n451), .B(KEYINPUT72), .ZN(n485) );
  XNOR2_X1 U501 ( .A(n513), .B(KEYINPUT27), .ZN(n461) );
  NOR2_X1 U502 ( .A1(n461), .A2(n509), .ZN(n452) );
  XNOR2_X1 U503 ( .A(n452), .B(KEYINPUT93), .ZN(n521) );
  XNOR2_X1 U504 ( .A(n459), .B(KEYINPUT67), .ZN(n453) );
  XNOR2_X1 U505 ( .A(n453), .B(KEYINPUT28), .ZN(n523) );
  NAND2_X1 U506 ( .A1(n523), .A2(n525), .ZN(n454) );
  NOR2_X1 U507 ( .A1(n521), .A2(n454), .ZN(n467) );
  XNOR2_X1 U508 ( .A(KEYINPUT94), .B(KEYINPUT95), .ZN(n455) );
  XNOR2_X1 U509 ( .A(n455), .B(KEYINPUT25), .ZN(n458) );
  NOR2_X1 U510 ( .A1(n513), .A2(n525), .ZN(n456) );
  NOR2_X1 U511 ( .A1(n459), .A2(n456), .ZN(n457) );
  XNOR2_X1 U512 ( .A(n458), .B(n457), .ZN(n463) );
  NAND2_X1 U513 ( .A1(n525), .A2(n459), .ZN(n460) );
  XNOR2_X1 U514 ( .A(n460), .B(KEYINPUT26), .ZN(n567) );
  NOR2_X1 U515 ( .A1(n461), .A2(n567), .ZN(n462) );
  NOR2_X1 U516 ( .A1(n463), .A2(n462), .ZN(n465) );
  INV_X1 U517 ( .A(n509), .ZN(n464) );
  NOR2_X1 U518 ( .A1(n465), .A2(n464), .ZN(n466) );
  NOR2_X1 U519 ( .A1(n467), .A2(n466), .ZN(n482) );
  INV_X1 U520 ( .A(n575), .ZN(n547) );
  NOR2_X1 U521 ( .A1(n534), .A2(n547), .ZN(n468) );
  XOR2_X1 U522 ( .A(KEYINPUT16), .B(n468), .Z(n469) );
  NOR2_X1 U523 ( .A1(n482), .A2(n469), .ZN(n470) );
  XNOR2_X1 U524 ( .A(KEYINPUT96), .B(n470), .ZN(n496) );
  NAND2_X1 U525 ( .A1(n485), .A2(n496), .ZN(n479) );
  NOR2_X1 U526 ( .A1(n509), .A2(n479), .ZN(n472) );
  XNOR2_X1 U527 ( .A(KEYINPUT34), .B(KEYINPUT97), .ZN(n471) );
  XNOR2_X1 U528 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U529 ( .A(G1GAT), .B(n473), .ZN(G1324GAT) );
  NOR2_X1 U530 ( .A1(n513), .A2(n479), .ZN(n474) );
  XOR2_X1 U531 ( .A(KEYINPUT98), .B(n474), .Z(n475) );
  XNOR2_X1 U532 ( .A(G8GAT), .B(n475), .ZN(G1325GAT) );
  NOR2_X1 U533 ( .A1(n525), .A2(n479), .ZN(n477) );
  XNOR2_X1 U534 ( .A(KEYINPUT99), .B(KEYINPUT35), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U536 ( .A(G15GAT), .B(n478), .Z(G1326GAT) );
  NOR2_X1 U537 ( .A1(n523), .A2(n479), .ZN(n480) );
  XOR2_X1 U538 ( .A(KEYINPUT100), .B(n480), .Z(n481) );
  XNOR2_X1 U539 ( .A(G22GAT), .B(n481), .ZN(G1327GAT) );
  XNOR2_X1 U540 ( .A(KEYINPUT102), .B(KEYINPUT39), .ZN(n488) );
  NOR2_X1 U541 ( .A1(n482), .A2(n575), .ZN(n483) );
  NAND2_X1 U542 ( .A1(n483), .A2(n578), .ZN(n484) );
  XNOR2_X1 U543 ( .A(KEYINPUT37), .B(n484), .ZN(n508) );
  NAND2_X1 U544 ( .A1(n485), .A2(n508), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n486), .B(KEYINPUT38), .ZN(n494) );
  NOR2_X1 U546 ( .A1(n509), .A2(n494), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U548 ( .A(G29GAT), .B(n489), .ZN(G1328GAT) );
  NOR2_X1 U549 ( .A1(n513), .A2(n494), .ZN(n490) );
  XOR2_X1 U550 ( .A(G36GAT), .B(n490), .Z(G1329GAT) );
  NOR2_X1 U551 ( .A1(n494), .A2(n525), .ZN(n492) );
  XNOR2_X1 U552 ( .A(KEYINPUT103), .B(KEYINPUT40), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U554 ( .A(G43GAT), .B(n493), .ZN(G1330GAT) );
  NOR2_X1 U555 ( .A1(n523), .A2(n494), .ZN(n495) );
  XOR2_X1 U556 ( .A(G50GAT), .B(n495), .Z(G1331GAT) );
  XOR2_X1 U557 ( .A(n541), .B(KEYINPUT104), .Z(n557) );
  AND2_X1 U558 ( .A1(n539), .A2(n557), .ZN(n507) );
  NAND2_X1 U559 ( .A1(n507), .A2(n496), .ZN(n503) );
  NOR2_X1 U560 ( .A1(n509), .A2(n503), .ZN(n498) );
  XNOR2_X1 U561 ( .A(KEYINPUT42), .B(KEYINPUT105), .ZN(n497) );
  XNOR2_X1 U562 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U563 ( .A(G57GAT), .B(n499), .ZN(G1332GAT) );
  NOR2_X1 U564 ( .A1(n513), .A2(n503), .ZN(n500) );
  XOR2_X1 U565 ( .A(KEYINPUT106), .B(n500), .Z(n501) );
  XNOR2_X1 U566 ( .A(G64GAT), .B(n501), .ZN(G1333GAT) );
  NOR2_X1 U567 ( .A1(n525), .A2(n503), .ZN(n502) );
  XOR2_X1 U568 ( .A(G71GAT), .B(n502), .Z(G1334GAT) );
  NOR2_X1 U569 ( .A1(n523), .A2(n503), .ZN(n505) );
  XNOR2_X1 U570 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n504) );
  XNOR2_X1 U571 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U572 ( .A(G78GAT), .B(n506), .Z(G1335GAT) );
  NAND2_X1 U573 ( .A1(n508), .A2(n507), .ZN(n517) );
  NOR2_X1 U574 ( .A1(n509), .A2(n517), .ZN(n511) );
  XNOR2_X1 U575 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U577 ( .A(G85GAT), .B(n512), .ZN(G1336GAT) );
  NOR2_X1 U578 ( .A1(n513), .A2(n517), .ZN(n514) );
  XOR2_X1 U579 ( .A(G92GAT), .B(n514), .Z(G1337GAT) );
  NOR2_X1 U580 ( .A1(n525), .A2(n517), .ZN(n515) );
  XOR2_X1 U581 ( .A(KEYINPUT110), .B(n515), .Z(n516) );
  XNOR2_X1 U582 ( .A(G99GAT), .B(n516), .ZN(G1338GAT) );
  NOR2_X1 U583 ( .A1(n523), .A2(n517), .ZN(n519) );
  XNOR2_X1 U584 ( .A(KEYINPUT111), .B(KEYINPUT44), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n520), .ZN(G1339GAT) );
  NOR2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n538) );
  NAND2_X1 U588 ( .A1(n538), .A2(n523), .ZN(n524) );
  NOR2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U590 ( .A(KEYINPUT114), .B(n526), .ZN(n533) );
  NAND2_X1 U591 ( .A1(n568), .A2(n533), .ZN(n527) );
  XNOR2_X1 U592 ( .A(G113GAT), .B(n527), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n529) );
  NAND2_X1 U594 ( .A1(n557), .A2(n533), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U596 ( .A(G120GAT), .B(n530), .Z(G1341GAT) );
  NAND2_X1 U597 ( .A1(n533), .A2(n575), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n531), .B(KEYINPUT50), .ZN(n532) );
  XNOR2_X1 U599 ( .A(G127GAT), .B(n532), .ZN(G1342GAT) );
  XOR2_X1 U600 ( .A(G134GAT), .B(KEYINPUT51), .Z(n536) );
  NAND2_X1 U601 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(G1343GAT) );
  INV_X1 U603 ( .A(n567), .ZN(n537) );
  NAND2_X1 U604 ( .A1(n538), .A2(n537), .ZN(n549) );
  NOR2_X1 U605 ( .A1(n539), .A2(n549), .ZN(n540) );
  XOR2_X1 U606 ( .A(G141GAT), .B(n540), .Z(G1344GAT) );
  NOR2_X1 U607 ( .A1(n541), .A2(n549), .ZN(n546) );
  XOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT117), .Z(n543) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U611 ( .A(KEYINPUT52), .B(n544), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(G1345GAT) );
  NOR2_X1 U613 ( .A1(n547), .A2(n549), .ZN(n548) );
  XOR2_X1 U614 ( .A(G155GAT), .B(n548), .Z(G1346GAT) );
  NOR2_X1 U615 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U616 ( .A(G162GAT), .B(n551), .Z(G1347GAT) );
  XNOR2_X1 U617 ( .A(G169GAT), .B(KEYINPUT118), .ZN(n553) );
  NAND2_X1 U618 ( .A1(n568), .A2(n560), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1348GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT57), .B(KEYINPUT120), .Z(n555) );
  XNOR2_X1 U621 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U623 ( .A(KEYINPUT119), .B(n556), .Z(n559) );
  NAND2_X1 U624 ( .A1(n557), .A2(n560), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  XOR2_X1 U626 ( .A(G183GAT), .B(KEYINPUT121), .Z(n562) );
  NAND2_X1 U627 ( .A1(n560), .A2(n575), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1350GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n564) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n565) );
  XOR2_X1 U632 ( .A(KEYINPUT123), .B(n565), .Z(n570) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n579) );
  NAND2_X1 U634 ( .A1(n579), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n573) );
  NAND2_X1 U637 ( .A1(n579), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U639 ( .A(G204GAT), .B(n574), .Z(G1353GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n579), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(KEYINPUT126), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G211GAT), .B(n577), .ZN(G1354GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n581) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

