//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n447, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n577, new_n579, new_n580,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n594, new_n595, new_n596,
    new_n597, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n641, new_n642, new_n645, new_n646,
    new_n648, new_n649, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  NAND2_X1  g021(.A1(G94), .A2(G452), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT66), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(new_n463), .A3(KEYINPUT3), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n469), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n474), .A2(G137), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n468), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g053(.A1(new_n468), .A2(KEYINPUT68), .A3(new_n473), .A4(new_n475), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n471), .A2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(new_n464), .ZN(new_n483));
  INV_X1    g058(.A(G125), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n463), .A2(G2105), .ZN(new_n486));
  AOI22_X1  g061(.A1(new_n485), .A2(G2105), .B1(G101), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n480), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G160));
  NAND2_X1  g064(.A1(new_n468), .A2(new_n473), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(new_n474), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G124), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT69), .B1(G100), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NOR3_X1   g069(.A1(KEYINPUT69), .A2(G100), .A3(G2105), .ZN(new_n495));
  OAI221_X1 g070(.A(G2104), .B1(G112), .B2(new_n474), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n490), .A2(G2105), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n497), .B1(G136), .B2(new_n498), .ZN(G162));
  NAND2_X1  g074(.A1(new_n474), .A2(G138), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n473), .A2(new_n467), .A3(new_n465), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT71), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n502), .A2(new_n505), .A3(KEYINPUT4), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n507));
  INV_X1    g082(.A(new_n483), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR4_X1   g085(.A1(new_n483), .A2(KEYINPUT72), .A3(KEYINPUT4), .A4(new_n500), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n504), .A2(new_n506), .A3(new_n512), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n468), .A2(G126), .A3(G2105), .A4(new_n473), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n515));
  INV_X1    g090(.A(G114), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n515), .B1(new_n516), .B2(G2105), .ZN(new_n517));
  NOR3_X1   g092(.A1(new_n474), .A2(KEYINPUT70), .A3(G114), .ZN(new_n518));
  OAI221_X1 g093(.A(G2104), .B1(G102), .B2(G2105), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n513), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(G164));
  OR2_X1    g097(.A1(KEYINPUT73), .A2(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT73), .A2(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(KEYINPUT6), .A3(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G543), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT6), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n526), .B1(new_n527), .B2(G651), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G50), .ZN(new_n530));
  AND2_X1   g105(.A1(KEYINPUT73), .A2(G651), .ZN(new_n531));
  NOR2_X1   g106(.A1(KEYINPUT73), .A2(G651), .ZN(new_n532));
  NOR3_X1   g107(.A1(new_n531), .A2(new_n532), .A3(new_n527), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n527), .A2(G651), .ZN(new_n534));
  AND2_X1   g109(.A1(KEYINPUT5), .A2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(KEYINPUT5), .A2(G543), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G88), .ZN(new_n539));
  NAND2_X1  g114(.A1(G75), .A2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n535), .A2(new_n536), .ZN(new_n541));
  INV_X1    g116(.A(G62), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n523), .A2(new_n524), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n530), .A2(new_n539), .A3(new_n545), .ZN(G303));
  INV_X1    g121(.A(G303), .ZN(G166));
  INV_X1    g122(.A(KEYINPUT5), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(new_n526), .ZN(new_n549));
  NAND2_X1  g124(.A1(KEYINPUT5), .A2(G543), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n549), .A2(new_n550), .B1(new_n527), .B2(G651), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n551), .A2(G89), .A3(new_n525), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n525), .A2(G51), .A3(new_n528), .ZN(new_n553));
  NAND3_X1  g128(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT7), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n549), .A2(new_n550), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n556), .A2(G63), .A3(G651), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n552), .A2(new_n553), .A3(new_n555), .A4(new_n557), .ZN(G286));
  INV_X1    g133(.A(G286), .ZN(G168));
  INV_X1    g134(.A(G64), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n560), .B1(new_n549), .B2(new_n550), .ZN(new_n561));
  AND2_X1   g136(.A1(G77), .A2(G543), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n544), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n525), .A2(new_n556), .A3(G90), .A4(new_n534), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n525), .A2(G52), .A3(new_n528), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G171));
  INV_X1    g142(.A(G56), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n568), .B1(new_n549), .B2(new_n550), .ZN(new_n569));
  AND2_X1   g144(.A1(G68), .A2(G543), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n544), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  XNOR2_X1  g146(.A(KEYINPUT74), .B(G81), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n551), .A2(new_n525), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n525), .A2(G43), .A3(new_n528), .ZN(new_n574));
  AND3_X1   g149(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G860), .ZN(G153));
  NAND4_X1  g151(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n577));
  XOR2_X1   g152(.A(new_n577), .B(KEYINPUT75), .Z(G176));
  NAND2_X1  g153(.A1(G1), .A2(G3), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT8), .ZN(new_n580));
  NAND4_X1  g155(.A1(G319), .A2(G483), .A3(G661), .A4(new_n580), .ZN(G188));
  NAND3_X1  g156(.A1(new_n525), .A2(G53), .A3(new_n528), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(KEYINPUT9), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT9), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n525), .A2(new_n584), .A3(G53), .A4(new_n528), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  AND3_X1   g161(.A1(KEYINPUT76), .A2(G78), .A3(G543), .ZN(new_n587));
  AOI21_X1  g162(.A(KEYINPUT76), .B1(G78), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(G65), .B1(new_n535), .B2(new_n536), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n538), .A2(G91), .B1(new_n591), .B2(G651), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n586), .A2(new_n592), .ZN(G299));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n566), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT77), .A4(new_n565), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G301));
  OAI21_X1  g173(.A(G651), .B1(new_n556), .B2(G74), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT78), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n599), .B(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(G49), .A2(new_n529), .B1(new_n538), .B2(G87), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(G288));
  NAND2_X1  g178(.A1(new_n529), .A2(G48), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n538), .A2(G86), .ZN(new_n605));
  NAND2_X1  g180(.A1(G73), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G61), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n541), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(new_n544), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n604), .A2(new_n605), .A3(new_n609), .ZN(G305));
  INV_X1    g185(.A(KEYINPUT79), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n551), .A2(G85), .A3(new_n525), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n525), .A2(G47), .A3(new_n528), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n612), .A2(new_n611), .A3(new_n613), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(G72), .A2(G543), .ZN(new_n618));
  INV_X1    g193(.A(G60), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n541), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(new_n544), .ZN(new_n621));
  AOI21_X1  g196(.A(KEYINPUT80), .B1(new_n617), .B2(new_n621), .ZN(new_n622));
  AND3_X1   g197(.A1(new_n612), .A2(new_n611), .A3(new_n613), .ZN(new_n623));
  OAI211_X1 g198(.A(KEYINPUT80), .B(new_n621), .C1(new_n623), .C2(new_n614), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(G290));
  NAND3_X1  g202(.A1(new_n551), .A2(G92), .A3(new_n525), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(KEYINPUT10), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT10), .ZN(new_n630));
  NAND4_X1  g205(.A1(new_n551), .A2(new_n630), .A3(new_n525), .A4(G92), .ZN(new_n631));
  INV_X1    g206(.A(G66), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n632), .B1(new_n549), .B2(new_n550), .ZN(new_n633));
  AND2_X1   g208(.A1(G79), .A2(G543), .ZN(new_n634));
  OAI21_X1  g209(.A(G651), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n525), .A2(G54), .A3(new_n528), .ZN(new_n636));
  NAND4_X1  g211(.A1(new_n629), .A2(new_n631), .A3(new_n635), .A4(new_n636), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n637), .A2(G868), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n638), .B1(G868), .B2(new_n597), .ZN(G284));
  AOI21_X1  g214(.A(new_n638), .B1(G868), .B2(new_n597), .ZN(G321));
  INV_X1    g215(.A(G868), .ZN(new_n641));
  NAND2_X1  g216(.A1(G299), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(new_n641), .B2(G168), .ZN(G297));
  OAI21_X1  g218(.A(new_n642), .B1(new_n641), .B2(G168), .ZN(G280));
  INV_X1    g219(.A(new_n637), .ZN(new_n645));
  INV_X1    g220(.A(G559), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n645), .B1(new_n646), .B2(G860), .ZN(G148));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(G868), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n649), .B1(G868), .B2(new_n575), .ZN(G323));
  XNOR2_X1  g225(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g226(.A1(new_n498), .A2(G135), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n491), .A2(G123), .ZN(new_n653));
  OR2_X1    g228(.A1(G99), .A2(G2105), .ZN(new_n654));
  OAI211_X1 g229(.A(new_n654), .B(G2104), .C1(G111), .C2(new_n474), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n652), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT82), .B(G2096), .Z(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n508), .A2(new_n486), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT13), .B(G2100), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n658), .A2(new_n659), .A3(new_n664), .ZN(G156));
  XNOR2_X1  g240(.A(G2427), .B(G2438), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2430), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT15), .B(G2435), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n669), .A2(KEYINPUT14), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1341), .B(G1348), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n671), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2451), .B(G2454), .Z(new_n676));
  XNOR2_X1  g251(.A(G2443), .B(G2446), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n675), .A2(new_n678), .ZN(new_n680));
  AND3_X1   g255(.A1(new_n679), .A2(G14), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT84), .ZN(G401));
  INV_X1    g257(.A(KEYINPUT18), .ZN(new_n683));
  XOR2_X1   g258(.A(G2084), .B(G2090), .Z(new_n684));
  XNOR2_X1  g259(.A(G2067), .B(G2678), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(KEYINPUT17), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n684), .A2(new_n685), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n683), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G2100), .ZN(new_n690));
  XOR2_X1   g265(.A(G2072), .B(G2078), .Z(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(new_n686), .B2(KEYINPUT18), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G2096), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n690), .B(new_n693), .ZN(G227));
  XOR2_X1   g269(.A(G1971), .B(G1976), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT19), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1956), .B(G2474), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1961), .B(G1966), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n697), .A2(new_n698), .ZN(new_n700));
  NOR3_X1   g275(.A1(new_n696), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n696), .A2(new_n699), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT20), .Z(new_n703));
  AOI211_X1 g278(.A(new_n701), .B(new_n703), .C1(new_n696), .C2(new_n700), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1991), .B(G1996), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1981), .B(G1986), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(G229));
  NAND2_X1  g285(.A1(new_n491), .A2(G119), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n474), .A2(G107), .ZN(new_n712));
  OAI21_X1  g287(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n498), .A2(G131), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT85), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(KEYINPUT85), .B1(new_n498), .B2(G131), .ZN(new_n717));
  OAI221_X1 g292(.A(new_n711), .B1(new_n712), .B2(new_n713), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  MUX2_X1   g293(.A(G25), .B(new_n718), .S(G29), .Z(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT35), .B(G1991), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n719), .B(new_n720), .Z(new_n721));
  NOR2_X1   g296(.A1(G16), .A2(G24), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n626), .B2(G16), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(G1986), .Z(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT86), .B(KEYINPUT34), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  MUX2_X1   g301(.A(G23), .B(G288), .S(G16), .Z(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT33), .B(G1976), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n727), .B(new_n728), .Z(new_n729));
  INV_X1    g304(.A(G16), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G22), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G166), .B2(new_n730), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G1971), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n730), .A2(G6), .ZN(new_n734));
  INV_X1    g309(.A(G305), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(new_n730), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT32), .B(G1981), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT87), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n736), .B(new_n738), .Z(new_n739));
  NOR3_X1   g314(.A1(new_n729), .A2(new_n733), .A3(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n721), .B(new_n724), .C1(new_n726), .C2(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT88), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n726), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(KEYINPUT36), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT36), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n743), .A2(new_n747), .A3(new_n744), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(G29), .A2(G35), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G162), .B2(G29), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(G2090), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT97), .Z(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT27), .B(G1996), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT93), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G29), .B2(G32), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n498), .A2(G141), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT91), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n491), .A2(G129), .ZN(new_n761));
  NAND3_X1  g336(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT26), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n764), .A2(new_n765), .B1(G105), .B2(new_n486), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n761), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n760), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT92), .ZN(new_n769));
  INV_X1    g344(.A(G29), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  MUX2_X1   g346(.A(new_n758), .B(new_n757), .S(new_n771), .Z(new_n772));
  AOI21_X1  g347(.A(new_n755), .B1(new_n756), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n756), .B2(new_n772), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n508), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n775), .A2(new_n474), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT89), .Z(new_n777));
  NAND2_X1  g352(.A1(new_n498), .A2(G139), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT25), .Z(new_n780));
  NAND3_X1  g355(.A1(new_n777), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  MUX2_X1   g356(.A(G33), .B(new_n781), .S(G29), .Z(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(G2072), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n730), .A2(G4), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n645), .B2(new_n730), .ZN(new_n785));
  INV_X1    g360(.A(G1348), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n730), .A2(G20), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT23), .Z(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G299), .B2(G16), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G1956), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT90), .B(KEYINPUT24), .ZN(new_n792));
  INV_X1    g367(.A(G34), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n770), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n793), .B2(new_n792), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n488), .B2(G29), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G2084), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n783), .A2(new_n787), .A3(new_n791), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n770), .A2(G27), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G164), .B2(new_n770), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G2078), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n770), .A2(G26), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT28), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n498), .A2(G140), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n491), .A2(G128), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n474), .A2(G116), .ZN(new_n807));
  OAI21_X1  g382(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n805), .B(new_n806), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n804), .B1(new_n809), .B2(G29), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G2067), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n730), .A2(G21), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G168), .B2(new_n730), .ZN(new_n813));
  NOR2_X1   g388(.A1(G16), .A2(G19), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n575), .B2(G16), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n813), .A2(G1966), .B1(new_n815), .B2(G1341), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n811), .B(new_n816), .C1(G1341), .C2(new_n815), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT31), .B(G11), .Z(new_n818));
  NAND2_X1  g393(.A1(G171), .A2(G16), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G5), .B2(G16), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT95), .B(G1961), .Z(new_n821));
  NOR2_X1   g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(G28), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n823), .A2(KEYINPUT30), .ZN(new_n824));
  AOI21_X1  g399(.A(G29), .B1(new_n823), .B2(KEYINPUT30), .ZN(new_n825));
  AOI211_X1 g400(.A(new_n818), .B(new_n822), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n656), .A2(new_n770), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n828), .A2(KEYINPUT94), .B1(new_n820), .B2(new_n821), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n813), .A2(G1966), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n828), .A2(KEYINPUT94), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n826), .A2(new_n829), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n817), .A2(new_n832), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n802), .B(new_n833), .C1(G2090), .C2(new_n753), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n774), .A2(new_n834), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n749), .A2(new_n835), .ZN(G311));
  NAND2_X1  g411(.A1(new_n749), .A2(new_n835), .ZN(G150));
  NOR2_X1   g412(.A1(new_n637), .A2(new_n646), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT38), .ZN(new_n839));
  INV_X1    g414(.A(G67), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(new_n549), .B2(new_n550), .ZN(new_n841));
  AND2_X1   g416(.A1(G80), .A2(G543), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n544), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n525), .A2(G55), .A3(new_n528), .ZN(new_n844));
  INV_X1    g419(.A(G93), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n551), .A2(new_n525), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n843), .B(new_n844), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n839), .B(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(KEYINPUT39), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(KEYINPUT39), .ZN(new_n852));
  XOR2_X1   g427(.A(KEYINPUT98), .B(G860), .Z(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n853), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n847), .A2(new_n855), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT37), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n854), .A2(new_n857), .ZN(G145));
  XOR2_X1   g433(.A(G162), .B(new_n656), .Z(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n488), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n809), .B(new_n521), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n768), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n862), .A2(KEYINPUT92), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n781), .B1(new_n862), .B2(KEYINPUT92), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT99), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n862), .A2(new_n781), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n498), .A2(G142), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n491), .A2(G130), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n474), .A2(G118), .ZN(new_n871));
  OAI21_X1  g446(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n869), .B(new_n870), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n718), .B(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n874), .A2(new_n662), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n662), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n875), .A2(KEYINPUT100), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(KEYINPUT100), .B1(new_n875), .B2(new_n876), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n863), .A2(KEYINPUT99), .A3(new_n864), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n868), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n879), .B1(new_n868), .B2(new_n880), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n860), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n875), .A2(new_n876), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n868), .A2(new_n880), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n860), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n868), .A2(new_n880), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n885), .B(new_n886), .C1(new_n887), .C2(new_n879), .ZN(new_n888));
  INV_X1    g463(.A(G37), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n883), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n883), .A2(new_n888), .A3(new_n889), .A4(new_n891), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(G395));
  NAND2_X1  g470(.A1(G299), .A2(new_n637), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n631), .A2(new_n635), .A3(new_n636), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n897), .A2(new_n586), .A3(new_n592), .A4(new_n629), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT41), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n899), .B1(new_n896), .B2(new_n898), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n902), .B1(new_n905), .B2(new_n901), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n575), .B(new_n847), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(new_n648), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n909), .A2(KEYINPUT103), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(KEYINPUT103), .ZN(new_n911));
  AOI22_X1  g486(.A1(new_n897), .A2(new_n629), .B1(new_n586), .B2(new_n592), .ZN(new_n912));
  NOR2_X1   g487(.A1(G299), .A2(new_n637), .ZN(new_n913));
  OR3_X1    g488(.A1(new_n908), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n910), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(G288), .B(new_n735), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n621), .B1(new_n623), .B2(new_n614), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT80), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n919), .A2(G303), .A3(new_n624), .ZN(new_n920));
  AOI21_X1  g495(.A(G303), .B1(new_n919), .B2(new_n624), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n916), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(G166), .B1(new_n622), .B2(new_n625), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n919), .A2(G303), .A3(new_n624), .ZN(new_n924));
  XNOR2_X1  g499(.A(G288), .B(G305), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT104), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n927), .B1(new_n928), .B2(KEYINPUT42), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n915), .B(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(KEYINPUT42), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n641), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n932), .B1(new_n931), .B2(new_n930), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT105), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT105), .B1(new_n847), .B2(new_n641), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n935), .B1(new_n933), .B2(new_n936), .ZN(G295));
  AOI21_X1  g512(.A(new_n935), .B1(new_n933), .B2(new_n936), .ZN(G331));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n939));
  AND2_X1   g514(.A1(G286), .A2(new_n566), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n940), .B1(new_n597), .B2(G168), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n907), .ZN(new_n942));
  AOI21_X1  g517(.A(G286), .B1(new_n595), .B2(new_n596), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n849), .B1(new_n943), .B2(new_n940), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n913), .A2(new_n912), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n942), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(new_n941), .B2(new_n907), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n849), .B(KEYINPUT106), .C1(new_n943), .C2(new_n940), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n948), .A2(new_n949), .B1(new_n907), .B2(new_n941), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT41), .B1(new_n913), .B2(new_n912), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n951), .A2(new_n901), .A3(new_n900), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n903), .A2(KEYINPUT102), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n946), .B1(new_n950), .B2(new_n954), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n922), .A2(new_n926), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n939), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n948), .A2(new_n949), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n942), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n906), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n960), .A2(KEYINPUT108), .A3(new_n927), .A4(new_n946), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT43), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n958), .A2(new_n945), .A3(new_n942), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n942), .A2(new_n944), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n963), .B1(new_n905), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(G37), .B1(new_n965), .B2(new_n956), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n962), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n927), .B1(new_n955), .B2(KEYINPUT107), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n960), .A2(new_n969), .A3(new_n946), .ZN(new_n970));
  AOI21_X1  g545(.A(G37), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n957), .A2(new_n961), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT43), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n967), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n962), .A2(new_n971), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n962), .A2(new_n971), .A3(KEYINPUT109), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n946), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n984), .B1(new_n959), .B2(new_n906), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT108), .B1(new_n985), .B2(new_n927), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n955), .A2(new_n956), .A3(new_n939), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n966), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n976), .B1(new_n988), .B2(KEYINPUT43), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n978), .B1(new_n983), .B2(new_n989), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n962), .A2(new_n971), .A3(KEYINPUT109), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT109), .B1(new_n962), .B2(new_n971), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n978), .B(new_n989), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n977), .B1(new_n990), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(KEYINPUT111), .B(new_n977), .C1(new_n990), .C2(new_n994), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(G397));
  INV_X1    g574(.A(G1384), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n521), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(KEYINPUT112), .B(G40), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n480), .A2(new_n487), .A3(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1006), .A2(G1996), .A3(new_n768), .ZN(new_n1007));
  XOR2_X1   g582(.A(new_n1007), .B(KEYINPUT113), .Z(new_n1008));
  XOR2_X1   g583(.A(new_n809), .B(G2067), .Z(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(new_n769), .B2(G1996), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1008), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n718), .A2(new_n720), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n718), .A2(new_n720), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1006), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g590(.A(new_n626), .B(G1986), .Z(new_n1016));
  AOI21_X1  g591(.A(new_n1015), .B1(new_n1006), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1001), .A2(KEYINPUT50), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n480), .A2(new_n487), .A3(new_n1004), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1384), .B1(new_n513), .B2(new_n520), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1019), .A2(new_n1020), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1961), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1002), .A2(G1384), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n521), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G2078), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n1029), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1003), .A2(G160), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1028), .A2(new_n1020), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1021), .A2(KEYINPUT45), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT114), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1005), .B1(new_n521), .B2(new_n1027), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1003), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(G2078), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1026), .B(new_n1031), .C1(new_n1038), .C2(KEYINPUT53), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G171), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT124), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1039), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1018), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT125), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1046), .A2(KEYINPUT53), .A3(new_n1029), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1047), .B(new_n1026), .C1(new_n1038), .C2(KEYINPUT53), .ZN(new_n1048));
  OR3_X1    g623(.A1(new_n1048), .A2(KEYINPUT123), .A3(new_n597), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT123), .B1(new_n1048), .B2(new_n597), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n1044), .A2(new_n1045), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1021), .A2(new_n1020), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(G2067), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n1024), .B2(new_n786), .ZN(new_n1055));
  OR2_X1    g630(.A1(new_n645), .A2(KEYINPUT120), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n645), .A2(KEYINPUT120), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1055), .A2(KEYINPUT60), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT60), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1005), .B1(new_n1001), .B2(KEYINPUT50), .ZN(new_n1060));
  AOI21_X1  g635(.A(G1348), .B1(new_n1060), .B2(new_n1023), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1059), .B1(new_n1061), .B2(new_n1054), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1061), .A2(new_n1059), .A3(new_n1054), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1058), .B(new_n1062), .C1(new_n1063), .C2(new_n1056), .ZN(new_n1064));
  INV_X1    g639(.A(G1956), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1024), .A2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT56), .B(G2072), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1046), .A2(new_n1067), .ZN(new_n1068));
  XOR2_X1   g643(.A(G299), .B(KEYINPUT57), .Z(new_n1069));
  NAND3_X1  g644(.A1(new_n1066), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1069), .ZN(new_n1071));
  AOI21_X1  g646(.A(G1956), .B1(new_n1060), .B2(new_n1023), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1067), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1032), .A2(new_n1033), .A3(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1071), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1070), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT61), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1070), .A2(new_n1075), .A3(KEYINPUT61), .ZN(new_n1079));
  INV_X1    g654(.A(G1996), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1003), .A2(new_n1080), .A3(new_n1036), .ZN(new_n1081));
  XOR2_X1   g656(.A(KEYINPUT58), .B(G1341), .Z(new_n1082));
  NAND2_X1  g657(.A1(new_n1053), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n848), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT59), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1084), .B(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1064), .A2(new_n1078), .A3(new_n1079), .A4(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1055), .A2(new_n637), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1069), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1070), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1048), .A2(new_n597), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1039), .A2(new_n597), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1018), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(G303), .A2(G8), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1096), .B(KEYINPUT55), .ZN(new_n1097));
  INV_X1    g672(.A(G1971), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1034), .A2(new_n1098), .A3(new_n1037), .ZN(new_n1099));
  INV_X1    g674(.A(G2090), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1060), .A2(new_n1100), .A3(new_n1023), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G8), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1097), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1103), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1097), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n1108));
  NAND2_X1  g683(.A1(G305), .A2(G1981), .ZN(new_n1109));
  INV_X1    g684(.A(G1981), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n604), .A2(new_n605), .A3(new_n1110), .A4(new_n609), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(KEYINPUT115), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT49), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1103), .B1(new_n1021), .B2(new_n1020), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT49), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1112), .A2(KEYINPUT115), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1114), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n601), .A2(G1976), .A3(new_n602), .ZN(new_n1119));
  INV_X1    g694(.A(G1976), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT52), .B1(G288), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1115), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT52), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1124), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1108), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1125), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1127), .A2(KEYINPUT116), .A3(new_n1122), .A4(new_n1118), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1104), .A2(new_n1107), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(G2084), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1019), .A2(new_n1131), .A3(new_n1020), .A4(new_n1023), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1132), .B(G168), .C1(new_n1046), .C2(G1966), .ZN(new_n1133));
  XNOR2_X1  g708(.A(KEYINPUT122), .B(KEYINPUT51), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n1133), .A2(G8), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT51), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1137), .B1(new_n1133), .B2(G8), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1132), .B1(new_n1046), .B2(G1966), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1140), .A2(G8), .A3(G286), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT121), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1140), .A2(KEYINPUT121), .A3(G8), .A4(G286), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1139), .A2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1092), .A2(new_n1095), .A3(new_n1130), .A4(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1045), .B1(new_n1044), .B2(new_n1051), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1052), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1105), .A2(new_n1106), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1118), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1152), .A2(G1976), .A3(G288), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1111), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1115), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1093), .A2(new_n1107), .A3(new_n1104), .A4(new_n1129), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT62), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1158), .B1(new_n1139), .B2(new_n1145), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1139), .A2(new_n1145), .A3(new_n1158), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1156), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1140), .A2(G8), .A3(G168), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1163), .A2(KEYINPUT63), .A3(new_n1150), .ZN(new_n1164));
  OR3_X1    g739(.A1(new_n1105), .A2(KEYINPUT118), .A3(new_n1106), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1105), .B1(KEYINPUT118), .B2(new_n1106), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1104), .A2(new_n1129), .A3(new_n1107), .A4(new_n1163), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1168), .A2(KEYINPUT117), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT63), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1170), .B1(new_n1168), .B2(KEYINPUT117), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1167), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1162), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1017), .B1(new_n1149), .B2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1009), .A2(new_n760), .A3(new_n767), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n1006), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT126), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1176), .B(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1006), .A2(new_n1080), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(KEYINPUT46), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT47), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1181), .B(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1006), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n809), .A2(G2067), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1015), .ZN(new_n1188));
  NOR3_X1   g763(.A1(new_n1184), .A2(G1986), .A3(G290), .ZN(new_n1189));
  XNOR2_X1  g764(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1189), .B(new_n1190), .ZN(new_n1191));
  AOI211_X1 g766(.A(new_n1183), .B(new_n1187), .C1(new_n1188), .C2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1174), .A2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g768(.A1(G229), .A2(new_n461), .A3(new_n681), .A4(G227), .ZN(new_n1195));
  NAND3_X1  g769(.A1(new_n890), .A2(new_n975), .A3(new_n1195), .ZN(G225));
  INV_X1    g770(.A(G225), .ZN(G308));
endmodule


