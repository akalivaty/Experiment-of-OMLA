//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n561, new_n563, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n583, new_n584, new_n585, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1209, new_n1210;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT67), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n463));
  AND3_X1   g038(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n463), .B1(new_n460), .B2(new_n462), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g043(.A(KEYINPUT69), .B1(new_n468), .B2(G2105), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  AOI211_X1 g046(.A(new_n470), .B(new_n471), .C1(new_n466), .C2(new_n467), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT70), .B1(new_n459), .B2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n460), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n459), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n475), .A2(new_n471), .A3(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n461), .A2(G2105), .ZN(new_n479));
  AOI22_X1  g054(.A1(new_n478), .A2(G137), .B1(G101), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n484));
  INV_X1    g059(.A(G136), .ZN(new_n485));
  INV_X1    g060(.A(G124), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n475), .A2(G2105), .A3(new_n476), .ZN(new_n487));
  OAI221_X1 g062(.A(new_n484), .B1(new_n477), .B2(new_n485), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND4_X1  g064(.A1(new_n475), .A2(G126), .A3(G2105), .A4(new_n476), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G114), .C2(new_n471), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n475), .A2(G138), .A3(new_n471), .A4(new_n476), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR3_X1   g071(.A1(new_n496), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n464), .B2(new_n465), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n493), .B1(new_n495), .B2(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(KEYINPUT71), .A3(KEYINPUT5), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n501), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n508), .A2(G88), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT72), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n510), .A2(new_n516), .A3(new_n513), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G62), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n507), .B2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n515), .A2(new_n517), .B1(G651), .B2(new_n520), .ZN(G166));
  AND2_X1   g096(.A1(new_n508), .A2(new_n509), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G89), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT75), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT7), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(new_n526), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n523), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G63), .ZN(new_n530));
  INV_X1    g105(.A(G651), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n508), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT73), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n508), .A2(KEYINPUT73), .A3(new_n532), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT74), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n512), .A2(G51), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(KEYINPUT73), .B1(new_n508), .B2(new_n532), .ZN(new_n541));
  NOR4_X1   g116(.A1(new_n507), .A2(new_n534), .A3(new_n530), .A4(new_n531), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n539), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT74), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n529), .B1(new_n540), .B2(new_n544), .ZN(G168));
  NAND2_X1  g120(.A1(new_n512), .A2(G52), .ZN(new_n546));
  INV_X1    g121(.A(new_n522), .ZN(new_n547));
  XNOR2_X1  g122(.A(KEYINPUT76), .B(G90), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n531), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n549), .A2(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  NAND2_X1  g128(.A1(new_n512), .A2(G43), .ZN(new_n554));
  INV_X1    g129(.A(G81), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n547), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(new_n531), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT77), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n561), .A2(new_n565), .ZN(G188));
  NAND2_X1  g141(.A1(KEYINPUT78), .A2(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n512), .A2(G53), .A3(new_n567), .ZN(new_n568));
  XNOR2_X1  g143(.A(KEYINPUT78), .B(KEYINPUT9), .ZN(new_n569));
  INV_X1    g144(.A(G53), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n511), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT79), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  XOR2_X1   g149(.A(new_n574), .B(KEYINPUT80), .Z(new_n575));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n507), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G651), .ZN(new_n578));
  INV_X1    g153(.A(G91), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n547), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n573), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G299));
  INV_X1    g157(.A(new_n529), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n538), .B1(new_n537), .B2(new_n539), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n543), .A2(KEYINPUT74), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(G286));
  INV_X1    g161(.A(G166), .ZN(G303));
  NAND2_X1  g162(.A1(new_n522), .A2(G87), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n512), .A2(G49), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(G288));
  NAND2_X1  g166(.A1(new_n512), .A2(G48), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n505), .A2(G86), .A3(new_n506), .A4(new_n509), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n505), .A2(G61), .A3(new_n506), .ZN(new_n596));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n531), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(G305));
  AOI22_X1  g175(.A1(new_n522), .A2(G85), .B1(G47), .B2(new_n512), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n531), .B2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n522), .A2(G92), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(KEYINPUT81), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT81), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n522), .A2(new_n607), .A3(G92), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n606), .A2(KEYINPUT10), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n507), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n612), .A2(G651), .B1(G54), .B2(new_n512), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g189(.A(KEYINPUT10), .B1(new_n606), .B2(new_n608), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n604), .B1(new_n616), .B2(G868), .ZN(G284));
  XNOR2_X1  g192(.A(G284), .B(KEYINPUT82), .ZN(G321));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G868), .B2(new_n581), .ZN(G297));
  OAI21_X1  g195(.A(new_n619), .B1(G868), .B2(new_n581), .ZN(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n616), .B1(new_n622), .B2(G860), .ZN(G148));
  INV_X1    g198(.A(new_n559), .ZN(new_n624));
  INV_X1    g199(.A(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n614), .A2(new_n615), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n627), .A2(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n626), .B1(new_n628), .B2(new_n625), .ZN(G323));
  XOR2_X1   g204(.A(KEYINPUT83), .B(KEYINPUT11), .Z(new_n630));
  XNOR2_X1  g205(.A(G323), .B(new_n630), .ZN(G282));
  NOR2_X1   g206(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n459), .A2(G2104), .ZN(new_n633));
  OAI21_X1  g208(.A(KEYINPUT68), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(new_n479), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT12), .Z(new_n638));
  XOR2_X1   g213(.A(KEYINPUT84), .B(G2100), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n638), .B(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n487), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(G123), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n478), .A2(G135), .ZN(new_n644));
  INV_X1    g219(.A(KEYINPUT85), .ZN(new_n645));
  NOR3_X1   g220(.A1(new_n645), .A2(new_n471), .A3(G111), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n645), .B1(new_n471), .B2(G111), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n647), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n643), .B(new_n644), .C1(new_n646), .C2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(G2096), .Z(new_n650));
  NAND2_X1  g225(.A1(new_n641), .A2(new_n650), .ZN(G156));
  INV_X1    g226(.A(KEYINPUT14), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2430), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2435), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2427), .B(G2438), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n652), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n656), .B1(new_n655), .B2(new_n654), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT16), .B(G1341), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G1348), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n660), .B(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(G14), .B1(new_n657), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n657), .B2(new_n663), .ZN(G401));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2067), .B(G2678), .Z(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2072), .B(G2078), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT18), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n667), .A2(new_n668), .ZN(new_n673));
  AND3_X1   g248(.A1(new_n673), .A2(KEYINPUT17), .A3(new_n670), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n670), .B1(new_n673), .B2(KEYINPUT17), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n674), .A2(new_n675), .A3(new_n669), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2096), .B(G2100), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n683), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n681), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT86), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n681), .B1(new_n688), .B2(new_n686), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(new_n688), .B2(new_n686), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT20), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n685), .B(new_n687), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(new_n691), .B2(new_n690), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1991), .ZN(new_n694));
  INV_X1    g269(.A(G1996), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1981), .B(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(G229));
  XNOR2_X1  g275(.A(KEYINPUT90), .B(G1341), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n559), .A2(new_n703), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n703), .A2(G19), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n702), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OR3_X1    g281(.A1(new_n704), .A2(new_n705), .A3(new_n702), .ZN(new_n707));
  NAND2_X1  g282(.A1(G171), .A2(G16), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G5), .B2(G16), .ZN(new_n709));
  INV_X1    g284(.A(G1961), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n706), .B(new_n707), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G2084), .ZN(new_n712));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(KEYINPUT24), .B2(G34), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(KEYINPUT24), .B2(G34), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n481), .B2(G29), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n711), .B1(new_n712), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n703), .A2(G20), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT97), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT23), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G299), .B2(G16), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G1956), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n479), .A2(G103), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT25), .Z(new_n724));
  INV_X1    g299(.A(G139), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(new_n477), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n636), .A2(G127), .ZN(new_n727));
  NAND2_X1  g302(.A1(G115), .A2(G2104), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n471), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OR3_X1    g304(.A1(new_n726), .A2(new_n729), .A3(new_n713), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G29), .B2(G33), .ZN(new_n731));
  INV_X1    g306(.A(G2072), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT91), .Z(new_n734));
  NAND3_X1  g309(.A1(new_n717), .A2(new_n722), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n731), .A2(new_n732), .ZN(new_n736));
  NOR2_X1   g311(.A1(G29), .A2(G32), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n478), .A2(G141), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT92), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n642), .A2(G129), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT26), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n743), .A2(new_n744), .B1(G105), .B2(new_n479), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n739), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n737), .B1(new_n748), .B2(G29), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT27), .B(G1996), .Z(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n736), .B(new_n751), .C1(new_n710), .C2(new_n709), .ZN(new_n752));
  NAND2_X1  g327(.A1(G168), .A2(G16), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G16), .B2(G21), .ZN(new_n754));
  INV_X1    g329(.A(G1966), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT30), .B(G28), .ZN(new_n757));
  OR2_X1    g332(.A1(KEYINPUT31), .A2(G11), .ZN(new_n758));
  NAND2_X1  g333(.A1(KEYINPUT31), .A2(G11), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n757), .A2(new_n713), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n649), .B2(new_n713), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT94), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n749), .A2(new_n750), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n752), .A2(new_n756), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n735), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n703), .A2(G4), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n616), .B2(new_n703), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT89), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1348), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n713), .A2(G26), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n642), .A2(G128), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n478), .A2(G140), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n471), .A2(G116), .ZN(new_n773));
  OAI21_X1  g348(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n771), .B(new_n772), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n770), .B1(new_n775), .B2(G29), .ZN(new_n776));
  MUX2_X1   g351(.A(new_n770), .B(new_n776), .S(KEYINPUT28), .Z(new_n777));
  INV_X1    g352(.A(G2067), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n713), .A2(G35), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G162), .B2(new_n713), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT29), .Z(new_n782));
  INV_X1    g357(.A(G2090), .ZN(new_n783));
  OAI22_X1  g358(.A1(new_n782), .A2(new_n783), .B1(new_n712), .B2(new_n716), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n779), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n782), .A2(new_n783), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT96), .Z(new_n787));
  NOR2_X1   g362(.A1(new_n754), .A2(new_n755), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT93), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n713), .A2(G27), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G164), .B2(new_n713), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT95), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G2078), .ZN(new_n793));
  NOR3_X1   g368(.A1(new_n787), .A2(new_n789), .A3(new_n793), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n765), .A2(new_n769), .A3(new_n785), .A4(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT98), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n703), .A2(G23), .ZN(new_n797));
  INV_X1    g372(.A(G288), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(new_n703), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT33), .B(G1976), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT88), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n799), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n703), .A2(G22), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G166), .B2(new_n703), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n804), .A2(G1971), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(G1971), .ZN(new_n806));
  MUX2_X1   g381(.A(G6), .B(G305), .S(G16), .Z(new_n807));
  XOR2_X1   g382(.A(KEYINPUT32), .B(G1981), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n802), .A2(new_n805), .A3(new_n806), .A4(new_n809), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT34), .Z(new_n811));
  NAND2_X1  g386(.A1(new_n713), .A2(G25), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n642), .A2(G119), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n478), .A2(G131), .ZN(new_n814));
  OR2_X1    g389(.A1(G95), .A2(G2105), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n815), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n812), .B1(new_n818), .B2(new_n713), .ZN(new_n819));
  MUX2_X1   g394(.A(new_n812), .B(new_n819), .S(KEYINPUT87), .Z(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT35), .B(G1991), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  MUX2_X1   g397(.A(G24), .B(G290), .S(G16), .Z(new_n823));
  INV_X1    g398(.A(G1986), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n820), .A2(new_n821), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n811), .A2(new_n822), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT36), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n796), .A2(new_n828), .ZN(G150));
  INV_X1    g404(.A(G150), .ZN(G311));
  NAND2_X1  g405(.A1(G80), .A2(G543), .ZN(new_n831));
  INV_X1    g406(.A(G67), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n507), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(G651), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n834), .A2(KEYINPUT99), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(KEYINPUT99), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n522), .A2(G93), .B1(G55), .B2(new_n512), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(new_n559), .B2(KEYINPUT100), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(KEYINPUT100), .B2(new_n559), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT100), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n624), .A2(new_n841), .A3(new_n838), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n616), .A2(G559), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n847));
  AOI21_X1  g422(.A(G860), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n847), .B2(new_n846), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n838), .A2(G860), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT102), .ZN(new_n851));
  XNOR2_X1  g426(.A(KEYINPUT101), .B(KEYINPUT37), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n849), .A2(new_n853), .ZN(G145));
  INV_X1    g429(.A(G142), .ZN(new_n855));
  NOR3_X1   g430(.A1(new_n471), .A2(KEYINPUT104), .A3(G118), .ZN(new_n856));
  OAI21_X1  g431(.A(KEYINPUT104), .B1(new_n471), .B2(G118), .ZN(new_n857));
  OR2_X1    g432(.A1(G106), .A2(G2105), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n857), .A2(G2104), .A3(new_n858), .ZN(new_n859));
  OAI22_X1  g434(.A1(new_n477), .A2(new_n855), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n860), .B1(G130), .B2(new_n642), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n747), .B(new_n861), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n726), .A2(new_n729), .A3(KEYINPUT103), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(new_n638), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n862), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n481), .B(G162), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n495), .A2(new_n498), .ZN(new_n868));
  INV_X1    g443(.A(new_n493), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n817), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n867), .B(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n649), .B(new_n775), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(G37), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(new_n872), .B2(new_n874), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g454(.A(G290), .B(G305), .Z(new_n880));
  XNOR2_X1  g455(.A(G166), .B(new_n798), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n880), .B(new_n881), .Z(new_n882));
  INV_X1    g457(.A(KEYINPUT107), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n882), .B1(new_n883), .B2(KEYINPUT42), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT108), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n883), .A2(KEYINPUT42), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n843), .B(new_n628), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n627), .A2(new_n581), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n616), .A2(G299), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT41), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n890), .A2(KEYINPUT41), .A3(new_n891), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n889), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n895), .A2(new_n889), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n888), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n898), .A2(new_n899), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n887), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n887), .A2(new_n903), .ZN(new_n905));
  OAI21_X1  g480(.A(G868), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n838), .A2(new_n625), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(G295));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n907), .ZN(G331));
  AOI21_X1  g484(.A(G301), .B1(new_n840), .B2(new_n842), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n840), .A2(G301), .A3(new_n842), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(G168), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n912), .ZN(new_n914));
  OAI21_X1  g489(.A(G286), .B1(new_n914), .B2(new_n910), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n913), .B(new_n915), .C1(new_n896), .C2(new_n897), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n913), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n892), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n916), .A2(new_n918), .A3(new_n882), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT109), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n916), .A2(new_n918), .ZN(new_n922));
  INV_X1    g497(.A(new_n882), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n916), .A2(new_n918), .A3(KEYINPUT109), .A4(new_n882), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n921), .A2(new_n924), .A3(new_n876), .A4(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(G37), .B1(new_n919), .B2(new_n920), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n917), .B1(new_n895), .B2(new_n894), .ZN(new_n930));
  INV_X1    g505(.A(new_n918), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n923), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AND4_X1   g507(.A1(KEYINPUT43), .A2(new_n929), .A3(new_n925), .A4(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT44), .B1(new_n928), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n926), .A2(KEYINPUT43), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n929), .A2(new_n927), .A3(new_n925), .A4(new_n932), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n934), .A2(new_n939), .ZN(G397));
  INV_X1    g515(.A(KEYINPUT127), .ZN(new_n941));
  INV_X1    g516(.A(G125), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(new_n634), .B2(new_n635), .ZN(new_n943));
  INV_X1    g518(.A(new_n467), .ZN(new_n944));
  OAI21_X1  g519(.A(G2105), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n470), .ZN(new_n946));
  OAI211_X1 g521(.A(KEYINPUT69), .B(G2105), .C1(new_n943), .C2(new_n944), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n946), .A2(G40), .A3(new_n480), .A4(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT45), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n949), .B1(G164), .B2(G1384), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n747), .B(new_n695), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n775), .B(new_n778), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n817), .A2(new_n821), .ZN(new_n955));
  OR2_X1    g530(.A1(new_n817), .A2(new_n821), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n953), .A2(new_n954), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(G290), .B(new_n824), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n952), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT61), .ZN(new_n961));
  INV_X1    g536(.A(new_n580), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT57), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(new_n963), .A3(new_n572), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n964), .B1(new_n581), .B2(new_n963), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT110), .B1(G164), .B2(G1384), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT110), .ZN(new_n968));
  INV_X1    g543(.A(G1384), .ZN(new_n969));
  AOI22_X1  g544(.A1(KEYINPUT4), .A2(new_n494), .B1(new_n636), .B2(new_n497), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n968), .B(new_n969), .C1(new_n970), .C2(new_n493), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n967), .A2(KEYINPUT50), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n948), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n972), .A2(KEYINPUT112), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT112), .B1(new_n972), .B2(new_n973), .ZN(new_n975));
  NOR3_X1   g550(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT116), .B1(new_n977), .B2(G1956), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n972), .A2(new_n973), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT112), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n972), .A2(KEYINPUT112), .A3(new_n973), .ZN(new_n982));
  INV_X1    g557(.A(new_n976), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT116), .ZN(new_n985));
  INV_X1    g560(.A(G1956), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n978), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g563(.A(KEYINPUT45), .B(new_n969), .C1(new_n970), .C2(new_n493), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n480), .A2(G40), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n950), .A2(new_n473), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  XOR2_X1   g566(.A(KEYINPUT56), .B(G2072), .Z(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n966), .B1(new_n988), .B2(new_n994), .ZN(new_n995));
  AOI211_X1 g570(.A(new_n965), .B(new_n993), .C1(new_n978), .C2(new_n987), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n961), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n987), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n985), .B1(new_n984), .B2(new_n986), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n994), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n965), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n988), .A2(new_n966), .A3(new_n994), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(new_n1002), .A3(KEYINPUT61), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n991), .A2(G1996), .ZN(new_n1004));
  XNOR2_X1  g579(.A(KEYINPUT58), .B(G1341), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n967), .A2(new_n971), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1005), .B1(new_n1006), .B2(new_n973), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n559), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT118), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT118), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1010), .B(new_n559), .C1(new_n1004), .C2(new_n1007), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1009), .A2(KEYINPUT59), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT59), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1008), .A2(KEYINPUT118), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1016), .A2(new_n473), .A3(G40), .A4(new_n480), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT50), .B1(new_n967), .B2(new_n971), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT117), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT50), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n968), .B1(new_n870), .B2(new_n969), .ZN(new_n1021));
  AOI211_X1 g596(.A(KEYINPUT110), .B(G1384), .C1(new_n868), .C2(new_n869), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1020), .B1(new_n870), .B2(new_n969), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1024), .A2(new_n948), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1023), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1019), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G1348), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1006), .A2(new_n973), .A3(new_n778), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT60), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n616), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1030), .A2(KEYINPUT60), .A3(new_n627), .A4(new_n1031), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1015), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n997), .A2(new_n1003), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n627), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n995), .B1(new_n1040), .B2(new_n1002), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT124), .ZN(new_n1043));
  AOI21_X1  g618(.A(G1961), .B1(new_n1019), .B2(new_n1027), .ZN(new_n1044));
  INV_X1    g619(.A(new_n991), .ZN(new_n1045));
  INV_X1    g620(.A(G2078), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT53), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT121), .B(G2078), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n945), .A2(KEYINPUT53), .A3(new_n1048), .ZN(new_n1049));
  AND4_X1   g624(.A1(new_n989), .A2(new_n950), .A3(new_n990), .A4(new_n1049), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1044), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(G171), .B1(new_n1051), .B2(KEYINPUT123), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT123), .ZN(new_n1053));
  NOR4_X1   g628(.A1(new_n1044), .A2(new_n1053), .A3(new_n1047), .A4(new_n1050), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1043), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1047), .B1(new_n1028), .B2(new_n710), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1050), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n1053), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1051), .A2(KEYINPUT123), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1059), .A2(KEYINPUT124), .A3(new_n1060), .A4(G171), .ZN(new_n1061));
  NOR3_X1   g636(.A1(G164), .A2(new_n949), .A3(G1384), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n948), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n967), .A2(new_n949), .A3(new_n971), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(new_n1046), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT120), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1063), .A2(new_n1067), .A3(new_n1064), .A4(new_n1046), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1066), .A2(KEYINPUT53), .A3(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1056), .A2(new_n1069), .A3(G301), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n1070), .A2(KEYINPUT54), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1055), .A2(new_n1061), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1006), .A2(new_n973), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n798), .A2(G1976), .ZN(new_n1074));
  INV_X1    g649(.A(G1976), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT52), .B1(G288), .B2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1073), .A2(G8), .A3(new_n1074), .A4(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G1981), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n595), .A2(new_n1078), .A3(new_n599), .ZN(new_n1079));
  OAI21_X1  g654(.A(G1981), .B1(new_n594), .B2(new_n598), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1079), .A2(KEYINPUT49), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT49), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1083), .A2(new_n1073), .A3(G8), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1073), .A2(G8), .A3(new_n1074), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1077), .B(new_n1084), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT111), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1023), .A2(new_n1025), .A3(new_n783), .ZN(new_n1090));
  INV_X1    g665(.A(G1971), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n991), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT55), .ZN(new_n1095));
  INV_X1    g670(.A(G8), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1095), .B1(G166), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  AND4_X1   g673(.A1(new_n1089), .A2(new_n1093), .A3(G8), .A4(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1096), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1089), .B1(new_n1100), .B2(new_n1098), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1088), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1092), .B1(new_n984), .B2(G2090), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1098), .B1(new_n1103), .B2(G8), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n1106));
  AOI21_X1  g681(.A(G301), .B1(new_n1056), .B2(new_n1069), .ZN(new_n1107));
  NOR4_X1   g682(.A1(new_n1044), .A2(G171), .A3(new_n1047), .A4(new_n1050), .ZN(new_n1108));
  OAI211_X1 g683(.A(KEYINPUT122), .B(new_n1106), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n1113));
  NAND3_X1  g688(.A1(G286), .A2(new_n1113), .A3(G8), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT119), .B1(G168), .B2(new_n1096), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n967), .A2(new_n949), .A3(new_n971), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n473), .A2(G40), .A3(new_n480), .A4(new_n989), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n755), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT113), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(G1966), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT113), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1023), .A2(new_n1025), .A3(new_n712), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1121), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1116), .B1(new_n1125), .B2(G8), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1017), .A2(new_n1018), .A3(G2084), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1128), .B1(new_n1120), .B2(new_n1119), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1127), .B1(new_n1129), .B2(new_n1123), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT51), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1124), .B1(new_n1122), .B2(KEYINPUT113), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1133));
  OAI21_X1  g708(.A(G8), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n1127), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT51), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1111), .A2(new_n1112), .B1(new_n1131), .B2(new_n1137), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1072), .A2(new_n1110), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1042), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1073), .A2(G8), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1084), .A2(new_n1075), .A3(new_n798), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1141), .B1(new_n1142), .B2(new_n1079), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1143), .B1(new_n1144), .B2(new_n1088), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT115), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1088), .B(new_n1146), .C1(new_n1098), .C2(new_n1100), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1100), .A2(new_n1098), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT111), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1100), .A2(new_n1089), .A3(new_n1098), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1100), .A2(new_n1098), .ZN(new_n1152));
  OAI21_X1  g727(.A(KEYINPUT115), .B1(new_n1152), .B2(new_n1087), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1147), .A2(new_n1151), .A3(KEYINPUT63), .A4(new_n1153), .ZN(new_n1154));
  OAI211_X1 g729(.A(G8), .B(G168), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT114), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1125), .A2(KEYINPUT114), .A3(G8), .A4(G168), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1154), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(KEYINPUT63), .B1(new_n1105), .B2(new_n1159), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1145), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1125), .A2(new_n1116), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1136), .B1(new_n1135), .B2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1126), .A2(KEYINPUT51), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT62), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT62), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1131), .A2(new_n1168), .A3(new_n1137), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1087), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1103), .A2(G8), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1098), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n1170), .A2(new_n1173), .A3(new_n1107), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n1167), .A2(new_n1169), .A3(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1163), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n960), .B1(new_n1140), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n954), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n951), .B1(new_n1178), .B2(new_n747), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n952), .A2(G1996), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1179), .B1(new_n1180), .B2(KEYINPUT46), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1181), .B1(KEYINPUT46), .B2(new_n1180), .ZN(new_n1182));
  XNOR2_X1  g757(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1182), .B(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n1185));
  OAI22_X1  g760(.A1(new_n1185), .A2(new_n956), .B1(G2067), .B2(new_n775), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n952), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1188), .B1(new_n1187), .B2(new_n1186), .ZN(new_n1189));
  OR3_X1    g764(.A1(new_n952), .A2(G1986), .A3(G290), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT48), .ZN(new_n1191));
  AOI22_X1  g766(.A1(new_n957), .A2(new_n951), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1192), .B1(new_n1191), .B2(new_n1190), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1184), .A2(new_n1189), .A3(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n941), .B1(new_n1177), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1194), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1159), .A2(new_n1173), .A3(new_n1170), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT63), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1144), .A2(new_n1198), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1200), .A2(new_n1159), .A3(new_n1153), .A4(new_n1147), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1167), .A2(new_n1169), .A3(new_n1174), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1202), .A2(new_n1203), .A3(new_n1145), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1204), .B1(new_n1042), .B2(new_n1139), .ZN(new_n1205));
  OAI211_X1 g780(.A(KEYINPUT127), .B(new_n1196), .C1(new_n1205), .C2(new_n960), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1195), .A2(new_n1206), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g782(.A(G319), .ZN(new_n1209));
  NOR4_X1   g783(.A1(G229), .A2(new_n1209), .A3(G401), .A4(G227), .ZN(new_n1210));
  NAND3_X1  g784(.A1(new_n937), .A2(new_n1210), .A3(new_n878), .ZN(G225));
  INV_X1    g785(.A(G225), .ZN(G308));
endmodule


