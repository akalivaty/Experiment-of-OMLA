//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n828,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(G211gat), .ZN(new_n203));
  INV_X1    g002(.A(G218gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n202), .B1(KEYINPUT22), .B2(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G211gat), .B(G218gat), .Z(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  NOR4_X1   g007(.A1(KEYINPUT70), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT70), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NOR3_X1   g012(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n209), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT71), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT71), .ZN(new_n220));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT26), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OR2_X1    g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n214), .B1(new_n225), .B2(new_n210), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n220), .B(new_n217), .C1(new_n226), .C2(new_n209), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT27), .B(G183gat), .ZN(new_n228));
  INV_X1    g027(.A(G190gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n228), .A2(KEYINPUT28), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT27), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT69), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n231), .B1(new_n232), .B2(G183gat), .ZN(new_n233));
  INV_X1    g032(.A(G183gat), .ZN(new_n234));
  NOR3_X1   g033(.A1(new_n234), .A2(KEYINPUT69), .A3(KEYINPUT27), .ZN(new_n235));
  NOR3_X1   g034(.A1(new_n233), .A2(new_n235), .A3(G190gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n230), .B1(new_n236), .B2(KEYINPUT28), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n227), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT23), .ZN(new_n239));
  NOR3_X1   g038(.A1(new_n239), .A2(G169gat), .A3(G176gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n239), .B1(G169gat), .B2(G176gat), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n241), .B1(new_n242), .B2(new_n212), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT24), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n217), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT64), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n248), .A2(new_n249), .B1(new_n234), .B2(new_n229), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(KEYINPUT65), .ZN(new_n252));
  NAND4_X1  g051(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n247), .A2(new_n250), .A3(new_n252), .A4(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n243), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT65), .B1(new_n217), .B2(new_n244), .ZN(new_n257));
  INV_X1    g056(.A(new_n253), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n259), .A2(KEYINPUT66), .A3(new_n250), .A4(new_n252), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT25), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n248), .A2(KEYINPUT67), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT67), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n263), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n234), .A2(new_n229), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n262), .A2(new_n264), .A3(new_n245), .A4(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n212), .B1(KEYINPUT23), .B2(new_n221), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT25), .ZN(new_n270));
  NOR3_X1   g069(.A1(new_n269), .A2(new_n270), .A3(new_n240), .ZN(new_n271));
  NOR2_X1   g070(.A1(G183gat), .A2(G190gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n251), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n273), .A2(KEYINPUT68), .A3(new_n262), .A4(new_n264), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n268), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n238), .B1(new_n261), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(G226gat), .A2(G233gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT74), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  OR2_X1    g078(.A1(new_n279), .A2(KEYINPUT77), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT29), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n254), .A2(new_n255), .ZN(new_n282));
  INV_X1    g081(.A(new_n243), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(new_n260), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n275), .B1(new_n284), .B2(new_n270), .ZN(new_n285));
  AND3_X1   g084(.A1(new_n219), .A2(new_n227), .A3(new_n237), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n281), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(new_n277), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n279), .A2(KEYINPUT77), .ZN(new_n289));
  AND4_X1   g088(.A1(new_n208), .A2(new_n280), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n208), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n292));
  INV_X1    g091(.A(new_n278), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n287), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n276), .A2(G226gat), .A3(G233gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n278), .B1(new_n276), .B2(new_n281), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(new_n292), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n291), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT76), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n270), .ZN(new_n301));
  INV_X1    g100(.A(new_n275), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n277), .B1(new_n303), .B2(new_n238), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n304), .B1(new_n297), .B2(new_n292), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT29), .B1(new_n303), .B2(new_n238), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT75), .B1(new_n306), .B2(new_n278), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT76), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n308), .A2(new_n309), .A3(new_n291), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n290), .B1(new_n300), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT30), .ZN(new_n312));
  XNOR2_X1  g111(.A(G8gat), .B(G36gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(G64gat), .B(G92gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n313), .B(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n311), .A2(new_n312), .A3(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G1gat), .B(G29gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n318), .B(KEYINPUT0), .ZN(new_n319));
  XNOR2_X1  g118(.A(G57gat), .B(G85gat), .ZN(new_n320));
  XOR2_X1   g119(.A(new_n319), .B(new_n320), .Z(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT72), .ZN(new_n323));
  INV_X1    g122(.A(G113gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n324), .A2(G120gat), .ZN(new_n325));
  INV_X1    g124(.A(G120gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(G113gat), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n323), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT1), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n326), .A2(G113gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n324), .A2(G120gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT72), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n328), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(G127gat), .B(G134gat), .Z(new_n334));
  INV_X1    g133(.A(KEYINPUT73), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n331), .B1(new_n325), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n336), .B1(new_n335), .B2(new_n331), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n334), .A2(KEYINPUT1), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n333), .A2(new_n334), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(G155gat), .ZN(new_n340));
  INV_X1    g139(.A(G162gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G155gat), .A2(G162gat), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OR2_X1    g143(.A1(KEYINPUT78), .A2(KEYINPUT2), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(KEYINPUT2), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G141gat), .B(G148gat), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n344), .B(new_n345), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n348), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n345), .A2(new_n342), .A3(new_n343), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n350), .A2(new_n351), .A3(new_n346), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n339), .B(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT5), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n355), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n358), .B1(new_n353), .B2(KEYINPUT3), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT3), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n349), .A2(KEYINPUT79), .A3(new_n352), .A4(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n333), .A2(new_n334), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n337), .A2(new_n338), .ZN(new_n364));
  AOI22_X1  g163(.A1(KEYINPUT3), .A2(new_n353), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n357), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n349), .A2(new_n352), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT4), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n339), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n368), .B1(new_n339), .B2(new_n367), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT80), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n363), .A2(new_n364), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT4), .B1(new_n373), .B2(new_n353), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n374), .A2(KEYINPUT80), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n366), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT81), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT81), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n366), .B(new_n378), .C1(new_n372), .C2(new_n375), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n356), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n362), .A2(new_n365), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n374), .A2(new_n369), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NOR3_X1   g182(.A1(new_n383), .A2(KEYINPUT5), .A3(new_n357), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n322), .B1(new_n380), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT39), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n386), .B1(new_n354), .B2(new_n355), .ZN(new_n387));
  INV_X1    g186(.A(new_n383), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n387), .B1(new_n388), .B2(new_n355), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n383), .A2(new_n386), .A3(new_n357), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n389), .A2(KEYINPUT40), .A3(new_n321), .A4(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(new_n321), .A3(new_n390), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT40), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AND3_X1   g193(.A1(new_n385), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n290), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n309), .B1(new_n308), .B2(new_n291), .ZN(new_n397));
  AOI211_X1 g196(.A(KEYINPUT76), .B(new_n208), .C1(new_n305), .C2(new_n307), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n396), .B(new_n316), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT30), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n300), .A2(new_n310), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n316), .B1(new_n401), .B2(new_n396), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n317), .B(new_n395), .C1(new_n400), .C2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT84), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n315), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(KEYINPUT30), .A3(new_n399), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n408), .A2(KEYINPUT84), .A3(new_n317), .A4(new_n395), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT37), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n280), .A2(new_n288), .A3(new_n289), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n411), .B1(new_n412), .B2(new_n291), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n308), .A2(new_n208), .ZN(new_n414));
  AOI211_X1 g213(.A(KEYINPUT38), .B(new_n316), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT85), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n406), .A2(new_n416), .A3(KEYINPUT37), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT85), .B1(new_n311), .B2(new_n411), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n415), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n356), .ZN(new_n420));
  INV_X1    g219(.A(new_n379), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n374), .A2(KEYINPUT80), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n370), .A2(new_n371), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(new_n423), .A3(new_n369), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n378), .B1(new_n424), .B2(new_n366), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n420), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n384), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n321), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n385), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  OAI211_X1 g229(.A(KEYINPUT6), .B(new_n322), .C1(new_n380), .C2(new_n384), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(new_n399), .A3(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n315), .B1(new_n311), .B2(new_n411), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n416), .B1(new_n406), .B2(KEYINPUT37), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n311), .A2(KEYINPUT85), .A3(new_n411), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT38), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n419), .B(new_n433), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n360), .B1(new_n291), .B2(KEYINPUT29), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n353), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n441), .A2(KEYINPUT82), .B1(G228gat), .B2(G233gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(G78gat), .B(G106gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT31), .B(G50gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  XOR2_X1   g244(.A(new_n442), .B(new_n445), .Z(new_n446));
  AOI21_X1  g245(.A(KEYINPUT29), .B1(new_n359), .B2(new_n361), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n441), .B1(new_n447), .B2(new_n208), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(G22gat), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT83), .ZN(new_n450));
  INV_X1    g249(.A(G22gat), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n441), .B(new_n451), .C1(new_n208), .C2(new_n447), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n449), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n450), .B1(new_n449), .B2(new_n452), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n446), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n455), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n442), .B(new_n445), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n458), .A3(new_n453), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n410), .A2(new_n439), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n303), .A2(new_n373), .A3(new_n238), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n276), .A2(new_n339), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(G227gat), .A2(G233gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n467), .A2(KEYINPUT34), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(KEYINPUT34), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n463), .A2(new_n464), .A3(G227gat), .A4(G233gat), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT33), .ZN(new_n472));
  XNOR2_X1  g271(.A(G15gat), .B(G43gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(G71gat), .B(G99gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n473), .B(new_n474), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n471), .B(KEYINPUT32), .C1(new_n472), .C2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n475), .B1(new_n471), .B2(new_n472), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n471), .A2(KEYINPUT32), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n470), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n470), .B1(new_n476), .B2(new_n479), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT36), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n470), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n479), .A2(new_n476), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT36), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(new_n487), .A3(new_n480), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n430), .A2(new_n431), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n491), .B1(new_n408), .B2(new_n317), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n490), .B1(new_n492), .B2(new_n461), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n462), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n408), .A2(new_n317), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n430), .A2(new_n431), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n460), .A2(new_n481), .A3(new_n482), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n499), .B(KEYINPUT35), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  XOR2_X1   g300(.A(G15gat), .B(G22gat), .Z(new_n502));
  INV_X1    g301(.A(G1gat), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n503), .A2(KEYINPUT16), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n502), .A2(new_n503), .ZN(new_n506));
  INV_X1    g305(.A(G8gat), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n505), .A2(new_n506), .B1(KEYINPUT90), .B2(new_n507), .ZN(new_n508));
  OR2_X1    g307(.A1(new_n507), .A2(KEYINPUT90), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n508), .B(new_n509), .Z(new_n510));
  XNOR2_X1  g309(.A(G43gat), .B(G50gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(KEYINPUT87), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT15), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(G29gat), .ZN(new_n515));
  INV_X1    g314(.A(G36gat), .ZN(new_n516));
  OR3_X1    g315(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT88), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT88), .B1(new_n515), .B2(new_n516), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT14), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n519), .B1(G29gat), .B2(G36gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT14), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n517), .A2(new_n518), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n511), .A2(KEYINPUT15), .ZN(new_n523));
  OR3_X1    g322(.A1(new_n514), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n514), .A2(KEYINPUT89), .A3(new_n522), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT89), .B1(new_n514), .B2(new_n522), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT17), .ZN(new_n529));
  INV_X1    g328(.A(new_n527), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(new_n525), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(new_n532), .A3(new_n524), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n510), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G229gat), .A2(G233gat), .ZN(new_n536));
  INV_X1    g335(.A(new_n528), .ZN(new_n537));
  INV_X1    g336(.A(new_n510), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n535), .A2(new_n536), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT18), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n528), .B(new_n510), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n536), .B(KEYINPUT13), .Z(new_n544));
  AOI22_X1  g343(.A1(new_n541), .A2(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n536), .ZN(new_n546));
  NOR3_X1   g345(.A1(new_n534), .A2(new_n539), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT18), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT91), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n549), .B1(new_n541), .B2(new_n542), .ZN(new_n550));
  XNOR2_X1  g349(.A(G113gat), .B(G141gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(KEYINPUT11), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT86), .ZN(new_n553));
  XNOR2_X1  g352(.A(G169gat), .B(G197gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT12), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n545), .B(new_n548), .C1(new_n550), .C2(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT91), .B1(new_n547), .B2(KEYINPUT18), .ZN(new_n558));
  INV_X1    g357(.A(new_n556), .ZN(new_n559));
  INV_X1    g358(.A(new_n548), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n544), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n561), .B1(new_n547), .B2(KEYINPUT18), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n558), .B(new_n559), .C1(new_n560), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n557), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n501), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT92), .ZN(new_n566));
  XNOR2_X1  g365(.A(G57gat), .B(G64gat), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT93), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G71gat), .B(G78gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT21), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G127gat), .B(G155gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT20), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n577), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G183gat), .B(G211gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n538), .B1(new_n572), .B2(new_n571), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n583), .B(KEYINPUT95), .Z(new_n584));
  XOR2_X1   g383(.A(new_n582), .B(new_n584), .Z(new_n585));
  NAND2_X1  g384(.A1(G85gat), .A2(G92gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT7), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT8), .ZN(new_n588));
  AND2_X1   g387(.A1(G99gat), .A2(G106gat), .ZN(new_n589));
  OAI221_X1 g388(.A(new_n587), .B1(new_n588), .B2(new_n589), .C1(G85gat), .C2(G92gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(G99gat), .A2(G106gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n590), .B(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n594), .B1(new_n529), .B2(new_n533), .ZN(new_n595));
  AND2_X1   g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n528), .A2(new_n594), .B1(KEYINPUT41), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G190gat), .B(G218gat), .ZN(new_n599));
  OR3_X1    g398(.A1(new_n595), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n599), .B1(new_n595), .B2(new_n598), .ZN(new_n601));
  XOR2_X1   g400(.A(G134gat), .B(G162gat), .Z(new_n602));
  NOR2_X1   g401(.A1(new_n596), .A2(KEYINPUT41), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n600), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT97), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n605), .B1(new_n600), .B2(new_n601), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT96), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n608), .B(new_n609), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n590), .B(new_n592), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n571), .ZN(new_n617));
  INV_X1    g416(.A(new_n571), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n594), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT98), .B(KEYINPUT10), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n617), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n594), .A2(KEYINPUT10), .A3(new_n618), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G230gat), .A2(G233gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n617), .A2(new_n619), .ZN(new_n626));
  INV_X1    g425(.A(new_n624), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G120gat), .B(G148gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(G176gat), .B(G204gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n625), .A2(new_n628), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT99), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n625), .A2(new_n628), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n631), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n566), .A2(new_n585), .A3(new_n615), .A4(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n639), .A2(new_n497), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(new_n503), .ZN(G1324gat));
  NOR2_X1   g440(.A1(new_n639), .A2(new_n496), .ZN(new_n642));
  OAI21_X1  g441(.A(KEYINPUT42), .B1(new_n642), .B2(new_n507), .ZN(new_n643));
  XOR2_X1   g442(.A(KEYINPUT16), .B(G8gat), .Z(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  MUX2_X1   g444(.A(KEYINPUT42), .B(new_n643), .S(new_n645), .Z(G1325gat));
  OAI21_X1  g445(.A(G15gat), .B1(new_n639), .B2(new_n490), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n481), .A2(new_n482), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n649), .A2(G15gat), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n647), .B1(new_n639), .B2(new_n650), .ZN(G1326gat));
  NOR2_X1   g450(.A1(new_n639), .A2(new_n461), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT43), .B(G22gat), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(G1327gat));
  XNOR2_X1  g453(.A(new_n582), .B(new_n584), .ZN(new_n655));
  AND4_X1   g454(.A1(new_n566), .A2(new_n655), .A3(new_n614), .A4(new_n638), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n656), .A2(new_n515), .A3(new_n491), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT45), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n659), .B1(new_n492), .B2(new_n461), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n399), .A2(KEYINPUT30), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n312), .B1(new_n311), .B2(new_n316), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n661), .B1(new_n407), .B2(new_n662), .ZN(new_n663));
  OAI211_X1 g462(.A(KEYINPUT100), .B(new_n460), .C1(new_n663), .C2(new_n491), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n462), .A2(new_n665), .A3(new_n490), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n615), .B1(new_n666), .B2(new_n500), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT101), .B(KEYINPUT44), .Z(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n316), .B1(new_n406), .B2(KEYINPUT37), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n670), .B1(new_n417), .B2(new_n418), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT38), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n435), .A2(new_n436), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n432), .B1(new_n673), .B2(new_n415), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n460), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n493), .B1(new_n675), .B2(new_n410), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n499), .A2(KEYINPUT35), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT35), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n678), .B1(new_n492), .B2(new_n498), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n614), .B1(new_n676), .B2(new_n680), .ZN(new_n681));
  AOI22_X1  g480(.A1(new_n667), .A2(new_n669), .B1(new_n681), .B2(KEYINPUT44), .ZN(new_n682));
  INV_X1    g481(.A(new_n564), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n655), .A2(new_n638), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(G29gat), .B1(new_n686), .B2(new_n497), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n658), .A2(new_n687), .ZN(G1328gat));
  NAND3_X1  g487(.A1(new_n656), .A2(new_n516), .A3(new_n663), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(KEYINPUT46), .Z(new_n690));
  OAI21_X1  g489(.A(G36gat), .B1(new_n686), .B2(new_n496), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(G1329gat));
  AOI21_X1  g491(.A(G43gat), .B1(new_n656), .B2(new_n648), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n489), .A2(G43gat), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n693), .B1(new_n685), .B2(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT102), .B(KEYINPUT47), .Z(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1330gat));
  NAND2_X1  g496(.A1(new_n656), .A2(new_n460), .ZN(new_n698));
  INV_X1    g497(.A(G50gat), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n685), .A2(G50gat), .A3(new_n460), .ZN(new_n701));
  AOI211_X1 g500(.A(KEYINPUT103), .B(KEYINPUT48), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  OR2_X1    g501(.A1(KEYINPUT103), .A2(KEYINPUT48), .ZN(new_n703));
  NAND2_X1  g502(.A1(KEYINPUT103), .A2(KEYINPUT48), .ZN(new_n704));
  AND4_X1   g503(.A1(new_n703), .A2(new_n700), .A3(new_n701), .A4(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n702), .A2(new_n705), .ZN(G1331gat));
  NAND2_X1  g505(.A1(new_n666), .A2(new_n500), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n585), .A2(new_n615), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n708), .A2(new_n564), .A3(new_n638), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n491), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT104), .B(G57gat), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1332gat));
  NAND2_X1  g512(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n710), .A2(new_n663), .A3(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n716), .B(KEYINPUT105), .Z(new_n717));
  XNOR2_X1  g516(.A(new_n715), .B(new_n717), .ZN(G1333gat));
  NAND2_X1  g517(.A1(new_n710), .A2(new_n489), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n649), .A2(G71gat), .ZN(new_n720));
  AOI22_X1  g519(.A1(new_n719), .A2(G71gat), .B1(new_n710), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g521(.A1(new_n710), .A2(new_n460), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT106), .B(G78gat), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1335gat));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n655), .A2(new_n683), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT107), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n637), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n727), .B1(new_n682), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n730), .ZN(new_n732));
  AOI211_X1 g531(.A(new_n615), .B(new_n668), .C1(new_n666), .C2(new_n500), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n734), .B1(new_n501), .B2(new_n614), .ZN(new_n735));
  OAI211_X1 g534(.A(KEYINPUT108), .B(new_n732), .C1(new_n733), .C2(new_n735), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n726), .B1(new_n738), .B2(new_n497), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n737), .A2(KEYINPUT109), .A3(new_n491), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n739), .A2(G85gat), .A3(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n667), .A2(KEYINPUT51), .A3(new_n729), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n667), .A2(new_n729), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n742), .B1(new_n745), .B2(KEYINPUT110), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n746), .B1(KEYINPUT110), .B2(new_n745), .ZN(new_n747));
  OR3_X1    g546(.A1(new_n638), .A2(G85gat), .A3(new_n497), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n741), .B1(new_n747), .B2(new_n748), .ZN(G1336gat));
  INV_X1    g548(.A(KEYINPUT113), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n731), .A2(new_n663), .A3(new_n736), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n751), .A2(new_n752), .A3(G92gat), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n752), .B1(new_n751), .B2(G92gat), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT112), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n745), .A2(new_n755), .A3(new_n742), .ZN(new_n756));
  OR3_X1    g555(.A1(new_n496), .A2(G92gat), .A3(new_n638), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n743), .A2(KEYINPUT112), .A3(new_n744), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n756), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n753), .A2(new_n754), .A3(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n750), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n760), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n751), .A2(G92gat), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n765), .B2(new_n752), .ZN(new_n766));
  OAI211_X1 g565(.A(KEYINPUT113), .B(KEYINPUT52), .C1(new_n766), .C2(new_n753), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n682), .A2(new_n730), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n663), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT52), .B1(new_n769), .B2(G92gat), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(new_n747), .B2(new_n757), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n763), .A2(new_n767), .A3(new_n771), .ZN(G1337gat));
  OAI21_X1  g571(.A(G99gat), .B1(new_n738), .B2(new_n490), .ZN(new_n773));
  OR3_X1    g572(.A1(new_n649), .A2(G99gat), .A3(new_n638), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n747), .B2(new_n774), .ZN(G1338gat));
  NAND2_X1  g574(.A1(new_n768), .A2(new_n460), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT53), .B1(new_n776), .B2(G106gat), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n638), .A2(new_n461), .A3(G106gat), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n777), .B1(new_n747), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n737), .A2(new_n460), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n756), .A2(new_n759), .ZN(new_n782));
  AOI22_X1  g581(.A1(new_n781), .A2(G106gat), .B1(new_n782), .B2(new_n778), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n780), .B1(new_n783), .B2(new_n784), .ZN(G1339gat));
  AOI21_X1  g584(.A(new_n536), .B1(new_n535), .B2(new_n540), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n543), .A2(new_n544), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n555), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n545), .A2(new_n556), .A3(new_n548), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n614), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n791), .B1(new_n623), .B2(new_n624), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n621), .A2(new_n622), .A3(new_n627), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n792), .A2(KEYINPUT114), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT114), .B1(new_n792), .B2(new_n793), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI211_X1 g596(.A(KEYINPUT54), .B(new_n627), .C1(new_n621), .C2(new_n622), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT115), .B1(new_n798), .B2(new_n632), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT115), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n800), .B(new_n631), .C1(new_n625), .C2(KEYINPUT54), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT55), .B1(new_n797), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n625), .A2(KEYINPUT54), .A3(new_n793), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n802), .A2(new_n808), .A3(new_n794), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT116), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n802), .A2(KEYINPUT55), .A3(new_n808), .A4(new_n794), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n813), .A2(new_n634), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n805), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n790), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n564), .A2(new_n805), .A3(new_n812), .A4(new_n814), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n637), .A2(new_n789), .A3(new_n788), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n614), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n655), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n585), .A2(new_n683), .A3(new_n615), .A4(new_n638), .ZN(new_n821));
  AOI211_X1 g620(.A(new_n497), .B(new_n663), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n498), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(new_n683), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(new_n324), .ZN(G1340gat));
  NOR2_X1   g624(.A1(new_n823), .A2(new_n638), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(new_n326), .ZN(G1341gat));
  NOR2_X1   g626(.A1(new_n823), .A2(new_n655), .ZN(new_n828));
  XOR2_X1   g627(.A(new_n828), .B(G127gat), .Z(G1342gat));
  AOI21_X1  g628(.A(new_n615), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n822), .A2(new_n498), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n832));
  XOR2_X1   g631(.A(new_n831), .B(new_n832), .Z(G1343gat));
  INV_X1    g632(.A(G141gat), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n489), .A2(new_n461), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n822), .A2(new_n834), .A3(new_n564), .A4(new_n835), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(KEYINPUT119), .ZN(new_n837));
  INV_X1    g636(.A(new_n821), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n790), .A2(new_n815), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n564), .A2(new_n811), .A3(new_n814), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n818), .A2(KEYINPUT117), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n637), .A2(new_n789), .A3(new_n843), .A4(new_n788), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n840), .A2(new_n841), .A3(new_n842), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n615), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n813), .A2(new_n634), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(new_n803), .ZN(new_n848));
  AOI22_X1  g647(.A1(new_n848), .A2(new_n564), .B1(new_n818), .B2(KEYINPUT117), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n842), .B1(new_n849), .B2(new_n844), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n839), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n838), .B1(new_n851), .B2(new_n655), .ZN(new_n852));
  OAI21_X1  g651(.A(KEYINPUT57), .B1(new_n852), .B2(new_n461), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n663), .A2(new_n497), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n490), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n461), .B1(new_n820), .B2(new_n821), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n853), .A2(new_n564), .A3(new_n858), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n859), .A2(G141gat), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT58), .B1(new_n837), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n836), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT120), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n834), .B1(new_n859), .B2(new_n864), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n853), .A2(KEYINPUT120), .A3(new_n564), .A4(new_n858), .ZN(new_n866));
  AOI211_X1 g665(.A(KEYINPUT121), .B(new_n863), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT121), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n859), .A2(new_n864), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(G141gat), .A3(new_n866), .ZN(new_n870));
  INV_X1    g669(.A(new_n863), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n868), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n861), .B1(new_n867), .B2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI211_X1 g674(.A(KEYINPUT122), .B(new_n861), .C1(new_n867), .C2(new_n872), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(G1344gat));
  NAND2_X1  g676(.A1(new_n822), .A2(new_n835), .ZN(new_n878));
  OR3_X1    g677(.A1(new_n878), .A2(G148gat), .A3(new_n638), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n856), .A2(KEYINPUT57), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n881), .B(KEYINPUT123), .Z(new_n882));
  OR2_X1    g681(.A1(new_n852), .A2(new_n461), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT124), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n883), .A2(new_n884), .A3(new_n857), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n884), .B1(new_n883), .B2(new_n857), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n882), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n888), .A2(new_n490), .A3(new_n637), .A4(new_n854), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n880), .B1(new_n889), .B2(G148gat), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n880), .A2(G148gat), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n853), .A2(new_n858), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n891), .B1(new_n892), .B2(new_n637), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n879), .B1(new_n890), .B2(new_n893), .ZN(G1345gat));
  NOR3_X1   g693(.A1(new_n878), .A2(G155gat), .A3(new_n655), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n892), .A2(new_n585), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(G155gat), .ZN(new_n897));
  XOR2_X1   g696(.A(new_n897), .B(KEYINPUT125), .Z(G1346gat));
  AOI21_X1  g697(.A(new_n341), .B1(new_n892), .B2(new_n614), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n878), .A2(G162gat), .A3(new_n615), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n899), .A2(new_n900), .ZN(G1347gat));
  NAND2_X1  g700(.A1(new_n663), .A2(new_n497), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n902), .B1(new_n820), .B2(new_n821), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n498), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n564), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g706(.A1(new_n905), .A2(new_n637), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(G176gat), .ZN(G1349gat));
  NOR2_X1   g708(.A1(new_n904), .A2(new_n655), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n228), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n911), .B1(new_n234), .B2(new_n910), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT60), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT127), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n912), .B(new_n915), .ZN(G1350gat));
  NAND2_X1  g715(.A1(new_n905), .A2(new_n614), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(G190gat), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT61), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n919), .B1(G190gat), .B2(new_n917), .ZN(G1351gat));
  NAND2_X1  g719(.A1(new_n903), .A2(new_n835), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(G197gat), .B1(new_n922), .B2(new_n564), .ZN(new_n923));
  INV_X1    g722(.A(new_n888), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n902), .A2(new_n489), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n564), .A2(G197gat), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n923), .B1(new_n927), .B2(new_n928), .ZN(G1352gat));
  NOR3_X1   g728(.A1(new_n921), .A2(G204gat), .A3(new_n638), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT62), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n924), .A2(new_n638), .A3(new_n926), .ZN(new_n932));
  INV_X1    g731(.A(G204gat), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(G1353gat));
  NAND3_X1  g733(.A1(new_n922), .A2(new_n203), .A3(new_n585), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n888), .A2(new_n585), .A3(new_n925), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n936), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT63), .B1(new_n936), .B2(G211gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(G1354gat));
  NAND3_X1  g738(.A1(new_n922), .A2(new_n204), .A3(new_n614), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n924), .A2(new_n615), .A3(new_n926), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(new_n204), .ZN(G1355gat));
endmodule


