//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992;
  INV_X1    g000(.A(G232gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  OR2_X1    g003(.A1(new_n204), .A2(KEYINPUT41), .ZN(new_n205));
  XNOR2_X1  g004(.A(G190gat), .B(G218gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT101), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n205), .B(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n206), .A2(new_n207), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT14), .ZN(new_n212));
  OR3_X1    g011(.A1(new_n212), .A2(G29gat), .A3(G36gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n212), .B1(G29gat), .B2(G36gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XOR2_X1   g014(.A(KEYINPUT89), .B(G29gat), .Z(new_n216));
  AOI22_X1  g015(.A1(new_n215), .A2(KEYINPUT88), .B1(G36gat), .B2(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(KEYINPUT88), .B2(new_n215), .ZN(new_n218));
  NAND2_X1  g017(.A1(G43gat), .A2(G50gat), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(G43gat), .A2(G50gat), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT15), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n215), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n216), .A2(G36gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n220), .A2(KEYINPUT15), .ZN(new_n227));
  XOR2_X1   g026(.A(KEYINPUT90), .B(G50gat), .Z(new_n228));
  OAI21_X1  g027(.A(new_n227), .B1(new_n228), .B2(G43gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n225), .A2(new_n226), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT91), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT17), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT100), .B(KEYINPUT7), .ZN(new_n235));
  NAND2_X1  g034(.A1(G85gat), .A2(G92gat), .ZN(new_n236));
  OR2_X1    g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n236), .ZN(new_n238));
  NOR2_X1   g037(.A1(G85gat), .A2(G92gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(G99gat), .A2(G106gat), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n239), .B1(KEYINPUT8), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n237), .A2(new_n238), .A3(new_n241), .ZN(new_n242));
  XOR2_X1   g041(.A(G99gat), .B(G106gat), .Z(new_n243));
  OR2_X1    g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n243), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n234), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n246), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n248), .A2(new_n231), .B1(KEYINPUT41), .B2(new_n204), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n211), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G134gat), .B(G162gat), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n250), .A2(new_n252), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n210), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n255), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n257), .A2(new_n209), .A3(new_n253), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(G57gat), .B(G64gat), .Z(new_n261));
  INV_X1    g060(.A(KEYINPUT9), .ZN(new_n262));
  INV_X1    g061(.A(G71gat), .ZN(new_n263));
  INV_X1    g062(.A(G78gat), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G71gat), .B(G78gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT97), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n261), .A2(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OR2_X1    g067(.A1(new_n266), .A2(new_n267), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n270), .A2(KEYINPUT21), .ZN(new_n271));
  NAND2_X1  g070(.A1(G231gat), .A2(G233gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  XOR2_X1   g072(.A(G127gat), .B(G155gat), .Z(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(KEYINPUT20), .ZN(new_n275));
  XOR2_X1   g074(.A(new_n273), .B(new_n275), .Z(new_n276));
  XNOR2_X1  g075(.A(G15gat), .B(G22gat), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT92), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT16), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n279), .B1(new_n280), .B2(G1gat), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT93), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n277), .B(KEYINPUT92), .ZN(new_n284));
  INV_X1    g083(.A(G1gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n283), .A2(new_n287), .A3(G8gat), .ZN(new_n288));
  INV_X1    g087(.A(G8gat), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n281), .B(new_n286), .C1(new_n282), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n291), .B1(KEYINPUT21), .B2(new_n270), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n292), .B(KEYINPUT99), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n276), .B(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G183gat), .B(G211gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n294), .B(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n260), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n270), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n246), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n244), .A2(new_n270), .A3(new_n245), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(KEYINPUT102), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT102), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n246), .A2(new_n304), .A3(new_n300), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT10), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT10), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G230gat), .ZN(new_n309));
  OAI22_X1  g108(.A1(new_n306), .A2(new_n308), .B1(new_n309), .B2(new_n203), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n309), .A2(new_n203), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n303), .A2(new_n312), .A3(new_n305), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G120gat), .B(G148gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(G176gat), .B(G204gat), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n315), .B(new_n316), .Z(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NOR3_X1   g117(.A1(new_n311), .A2(new_n314), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n318), .B1(new_n311), .B2(new_n314), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n299), .A2(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n288), .A2(new_n290), .ZN(new_n325));
  INV_X1    g124(.A(new_n231), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n291), .A2(new_n231), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(KEYINPUT94), .A3(new_n328), .ZN(new_n329));
  OR3_X1    g128(.A1(new_n325), .A2(KEYINPUT94), .A3(new_n326), .ZN(new_n330));
  NAND2_X1  g129(.A1(G229gat), .A2(G233gat), .ZN(new_n331));
  XOR2_X1   g130(.A(new_n331), .B(KEYINPUT13), .Z(new_n332));
  NAND3_X1  g131(.A1(new_n329), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT95), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n329), .A2(new_n330), .A3(KEYINPUT95), .A4(new_n332), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n232), .A2(new_n233), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT17), .B1(new_n231), .B2(KEYINPUT91), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n331), .B(new_n328), .C1(new_n340), .C2(new_n291), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT18), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n234), .A2(new_n325), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT18), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n343), .A2(new_n344), .A3(new_n331), .A4(new_n328), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n337), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G113gat), .B(G141gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(G197gat), .ZN(new_n349));
  XOR2_X1   g148(.A(KEYINPUT11), .B(G169gat), .Z(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n351), .B(KEYINPUT12), .Z(new_n352));
  NAND2_X1  g151(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n335), .A2(new_n336), .B1(new_n342), .B2(new_n345), .ZN(new_n354));
  INV_X1    g153(.A(new_n352), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT71), .ZN(new_n358));
  NOR2_X1   g157(.A1(G169gat), .A2(G176gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT26), .ZN(new_n360));
  NAND2_X1  g159(.A1(G183gat), .A2(G190gat), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT26), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n362), .B1(G169gat), .B2(G176gat), .ZN(new_n363));
  AND2_X1   g162(.A1(G169gat), .A2(G176gat), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n360), .B(new_n361), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(G183gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT27), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT27), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G183gat), .ZN(new_n369));
  INV_X1    g168(.A(G190gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT28), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT27), .B(G183gat), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n374), .A2(KEYINPUT28), .A3(new_n370), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n365), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G169gat), .ZN(new_n377));
  INV_X1    g176(.A(G176gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT23), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n364), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT24), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n361), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n370), .ZN(new_n384));
  NAND3_X1  g183(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n380), .A2(G176gat), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT64), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n377), .ZN(new_n389));
  NAND2_X1  g188(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n387), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n381), .A2(new_n386), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT25), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT65), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n361), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT66), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT66), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT24), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n396), .A2(new_n397), .A3(new_n398), .A4(new_n400), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n384), .A2(new_n385), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n377), .A2(new_n378), .A3(KEYINPUT23), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT25), .ZN(new_n405));
  NAND2_X1  g204(.A1(G169gat), .A2(G176gat), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n406), .B1(new_n359), .B2(KEYINPUT23), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n403), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n376), .B1(new_n394), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(G113gat), .ZN(new_n411));
  AND2_X1   g210(.A1(new_n411), .A2(G120gat), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(G120gat), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT68), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G113gat), .B(G120gat), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT68), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT1), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n414), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(G127gat), .A2(G134gat), .ZN(new_n420));
  INV_X1    g219(.A(G134gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT67), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT67), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(G134gat), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n420), .B1(new_n425), .B2(G127gat), .ZN(new_n426));
  AND2_X1   g225(.A1(G127gat), .A2(G134gat), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n418), .B1(new_n427), .B2(new_n420), .ZN(new_n428));
  AND2_X1   g227(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n429));
  NOR2_X1   g228(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n429), .A2(new_n430), .A3(new_n411), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT70), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n428), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OR2_X1    g232(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(G113gat), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n411), .A2(G120gat), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(KEYINPUT70), .A3(new_n437), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n419), .A2(new_n426), .B1(new_n433), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n358), .B1(new_n410), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G227gat), .A2(G233gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n394), .A2(new_n409), .ZN(new_n443));
  INV_X1    g242(.A(new_n376), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n439), .A2(new_n443), .A3(new_n358), .A4(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n418), .B1(new_n415), .B2(new_n416), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n412), .A2(new_n413), .A3(KEYINPUT68), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n426), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n428), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n434), .A2(new_n432), .A3(G113gat), .A4(new_n435), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n437), .A2(KEYINPUT70), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n449), .B(new_n450), .C1(new_n431), .C2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n393), .A2(new_n392), .B1(new_n403), .B2(new_n408), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n453), .B1(new_n454), .B2(new_n376), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n441), .A2(new_n442), .A3(new_n445), .A4(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT74), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n457), .A2(KEYINPUT34), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(KEYINPUT34), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n456), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n459), .B1(new_n456), .B2(new_n458), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n442), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n455), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n463), .B1(new_n464), .B2(new_n440), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT33), .ZN(new_n466));
  XNOR2_X1  g265(.A(G15gat), .B(G43gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(G71gat), .B(G99gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n467), .B(new_n468), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n465), .B(KEYINPUT32), .C1(new_n466), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n465), .A2(KEYINPUT32), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT73), .ZN(new_n472));
  INV_X1    g271(.A(new_n469), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT73), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n465), .A2(new_n474), .A3(KEYINPUT32), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n472), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n465), .A2(KEYINPUT72), .A3(new_n466), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT72), .B1(new_n465), .B2(new_n466), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n462), .B(new_n470), .C1(new_n476), .C2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n469), .B1(new_n471), .B2(KEYINPUT73), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n482), .B(new_n475), .C1(new_n478), .C2(new_n477), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n462), .B1(new_n483), .B2(new_n470), .ZN(new_n484));
  NAND2_X1  g283(.A1(G155gat), .A2(G162gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT2), .ZN(new_n486));
  INV_X1    g285(.A(G141gat), .ZN(new_n487));
  INV_X1    g286(.A(G148gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(G141gat), .A2(G148gat), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n486), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  OR2_X1    g290(.A1(G155gat), .A2(G162gat), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT77), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n492), .A2(new_n493), .A3(new_n485), .ZN(new_n494));
  AND2_X1   g293(.A1(G155gat), .A2(G162gat), .ZN(new_n495));
  NOR2_X1   g294(.A1(G155gat), .A2(G162gat), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT77), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n491), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n495), .A2(new_n496), .ZN(new_n499));
  AND2_X1   g298(.A1(G141gat), .A2(G148gat), .ZN(new_n500));
  NOR2_X1   g299(.A1(G141gat), .A2(G148gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n499), .A2(new_n502), .A3(new_n493), .A4(new_n486), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(G211gat), .A2(G218gat), .ZN(new_n506));
  INV_X1    g305(.A(G211gat), .ZN(new_n507));
  INV_X1    g306(.A(G218gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g308(.A1(G197gat), .A2(G204gat), .ZN(new_n510));
  NOR2_X1   g309(.A1(G197gat), .A2(G204gat), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT22), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n506), .B(new_n509), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n509), .A2(new_n506), .ZN(new_n515));
  XNOR2_X1  g314(.A(G197gat), .B(G204gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n506), .A2(new_n513), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT29), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n505), .B1(new_n519), .B2(KEYINPUT3), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n514), .A2(new_n518), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT3), .B1(new_n498), .B2(new_n503), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n522), .B1(new_n523), .B2(KEYINPUT29), .ZN(new_n524));
  INV_X1    g323(.A(G228gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n525), .A2(new_n203), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n520), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT3), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT81), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n528), .B1(new_n519), .B2(new_n529), .ZN(new_n530));
  AOI211_X1 g329(.A(KEYINPUT81), .B(KEYINPUT29), .C1(new_n514), .C2(new_n518), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n505), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n524), .ZN(new_n533));
  INV_X1    g332(.A(new_n526), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT82), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT82), .ZN(new_n536));
  AOI211_X1 g335(.A(new_n536), .B(new_n526), .C1(new_n532), .C2(new_n524), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n527), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(G22gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT83), .ZN(new_n540));
  INV_X1    g339(.A(G22gat), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n541), .B(new_n527), .C1(new_n535), .C2(new_n537), .ZN(new_n542));
  XNOR2_X1  g341(.A(G78gat), .B(G106gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT80), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT31), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n545), .B(G50gat), .Z(new_n546));
  NAND4_X1  g345(.A1(new_n539), .A2(new_n540), .A3(new_n542), .A4(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n542), .A2(KEYINPUT83), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n549), .A2(new_n546), .B1(new_n539), .B2(new_n542), .ZN(new_n550));
  OAI22_X1  g349(.A1(new_n481), .A2(new_n484), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT86), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(G226gat), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n554), .A2(new_n203), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT75), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n557), .B1(new_n454), .B2(new_n376), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n443), .A2(new_n444), .A3(KEYINPUT75), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n556), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NOR3_X1   g359(.A1(new_n410), .A2(KEYINPUT29), .A3(new_n555), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n521), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n555), .A2(KEYINPUT29), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n558), .A2(new_n559), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n410), .A2(new_n555), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n564), .A2(new_n522), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G8gat), .B(G36gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(G64gat), .B(G92gat), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n567), .B(new_n568), .Z(new_n569));
  NAND3_X1  g368(.A1(new_n562), .A2(new_n566), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT30), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n562), .A2(KEYINPUT30), .A3(new_n566), .A4(new_n569), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n569), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n562), .A2(new_n566), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(KEYINPUT76), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT76), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n579), .B1(new_n562), .B2(new_n566), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n576), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n575), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G1gat), .B(G29gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT0), .ZN(new_n584));
  XNOR2_X1  g383(.A(G57gat), .B(G85gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n584), .B(new_n585), .Z(new_n586));
  NAND3_X1  g385(.A1(new_n448), .A2(new_n504), .A3(new_n452), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT4), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT4), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n448), .A2(new_n504), .A3(new_n452), .A4(new_n589), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n498), .A2(new_n503), .A3(KEYINPUT3), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n591), .A2(new_n523), .ZN(new_n592));
  AOI22_X1  g391(.A1(new_n588), .A2(new_n590), .B1(new_n592), .B2(new_n453), .ZN(new_n593));
  NAND2_X1  g392(.A1(G225gat), .A2(G233gat), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n594), .B(KEYINPUT78), .Z(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n587), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n504), .B1(new_n448), .B2(new_n452), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n595), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n593), .A2(new_n596), .B1(new_n599), .B2(KEYINPUT5), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n588), .A2(new_n590), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n592), .A2(new_n453), .ZN(new_n602));
  AND4_X1   g401(.A1(KEYINPUT5), .A2(new_n601), .A3(new_n596), .A4(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n586), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n593), .A2(new_n596), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n599), .A2(KEYINPUT5), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n586), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n593), .A2(KEYINPUT5), .A3(new_n596), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(KEYINPUT79), .B(KEYINPUT6), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n604), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n611), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n607), .A2(new_n608), .A3(new_n609), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n582), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n549), .A2(new_n546), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n539), .A2(new_n542), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(new_n547), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n621), .B(KEYINPUT86), .C1(new_n481), .C2(new_n484), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n553), .A2(new_n617), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT35), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT35), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n615), .A2(new_n575), .A3(new_n625), .A4(new_n581), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n626), .B1(new_n547), .B2(new_n620), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n483), .A2(new_n470), .ZN(new_n628));
  INV_X1    g427(.A(new_n462), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n630), .A2(KEYINPUT85), .A3(new_n480), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT85), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n632), .B1(new_n481), .B2(new_n484), .ZN(new_n633));
  AND3_X1   g432(.A1(new_n627), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n624), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n582), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n593), .A2(new_n596), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n638), .A2(KEYINPUT39), .ZN(new_n639));
  OR3_X1    g438(.A1(new_n597), .A2(new_n598), .A3(new_n595), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n638), .A2(KEYINPUT39), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n639), .A2(new_n586), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT40), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n639), .A2(KEYINPUT40), .A3(new_n586), .A4(new_n641), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n644), .A2(new_n610), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n621), .B1(new_n637), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n577), .A2(KEYINPUT37), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n648), .A2(new_n569), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT38), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n522), .B1(new_n560), .B2(new_n561), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n564), .A2(new_n521), .A3(new_n565), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n651), .A2(KEYINPUT37), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n649), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n616), .A2(new_n570), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT37), .B1(new_n578), .B2(new_n580), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n650), .B1(new_n656), .B2(new_n649), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n647), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT84), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n621), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n620), .A2(KEYINPUT84), .A3(new_n547), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n617), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n630), .A2(KEYINPUT36), .A3(new_n480), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT36), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n665), .B1(new_n481), .B2(new_n484), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  OR3_X1    g466(.A1(new_n659), .A2(new_n663), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(KEYINPUT87), .B1(new_n636), .B2(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n634), .B1(new_n623), .B2(KEYINPUT35), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n659), .A2(new_n663), .A3(new_n667), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT87), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n357), .B1(new_n669), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(KEYINPUT96), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n636), .A2(KEYINPUT87), .A3(new_n668), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n672), .B1(new_n670), .B2(new_n671), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT96), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n678), .A2(new_n679), .A3(new_n357), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n324), .B1(new_n675), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n616), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G1gat), .ZN(G1324gat));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT16), .B(G8gat), .Z(new_n685));
  NAND3_X1  g484(.A1(new_n681), .A2(new_n582), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n324), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n679), .B1(new_n678), .B2(new_n357), .ZN(new_n688));
  INV_X1    g487(.A(new_n357), .ZN(new_n689));
  AOI211_X1 g488(.A(KEYINPUT96), .B(new_n689), .C1(new_n676), .C2(new_n677), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n582), .B(new_n687), .C1(new_n688), .C2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(G8gat), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n686), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(KEYINPUT42), .ZN(new_n694));
  INV_X1    g493(.A(new_n691), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT42), .B1(new_n695), .B2(new_n685), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n684), .B1(new_n694), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT42), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n699), .B1(new_n686), .B2(new_n692), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n700), .A2(new_n696), .A3(KEYINPUT103), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n698), .A2(new_n701), .ZN(G1325gat));
  INV_X1    g501(.A(new_n681), .ZN(new_n703));
  INV_X1    g502(.A(new_n667), .ZN(new_n704));
  OAI21_X1  g503(.A(G15gat), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n631), .A2(new_n633), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n706), .A2(G15gat), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n705), .B1(new_n703), .B2(new_n707), .ZN(G1326gat));
  INV_X1    g507(.A(new_n661), .ZN(new_n709));
  INV_X1    g508(.A(new_n662), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n681), .A2(new_n712), .ZN(new_n713));
  OR2_X1    g512(.A1(new_n713), .A2(KEYINPUT104), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(KEYINPUT104), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT43), .B(G22gat), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n716), .B1(new_n714), .B2(new_n715), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(G1327gat));
  NAND2_X1  g518(.A1(new_n298), .A2(new_n323), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(new_n259), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(new_n688), .B2(new_n690), .ZN(new_n722));
  OR3_X1    g521(.A1(new_n722), .A2(new_n615), .A3(new_n216), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n724));
  OR2_X1    g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n259), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n260), .B1(new_n670), .B2(new_n671), .ZN(new_n728));
  AOI22_X1  g527(.A1(new_n678), .A2(new_n727), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n720), .A2(new_n689), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OR3_X1    g530(.A1(new_n731), .A2(KEYINPUT105), .A3(new_n615), .ZN(new_n732));
  OAI21_X1  g531(.A(KEYINPUT105), .B1(new_n731), .B2(new_n615), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n732), .A2(new_n216), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n723), .A2(new_n724), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n725), .A2(new_n734), .A3(new_n735), .ZN(G1328gat));
  NOR2_X1   g535(.A1(new_n637), .A2(G36gat), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n721), .B(new_n737), .C1(new_n688), .C2(new_n690), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(KEYINPUT106), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT46), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n738), .A2(KEYINPUT106), .ZN(new_n742));
  OR3_X1    g541(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n741), .B1(new_n740), .B2(new_n742), .ZN(new_n744));
  OAI21_X1  g543(.A(G36gat), .B1(new_n731), .B2(new_n637), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(G1329gat));
  OAI21_X1  g545(.A(G43gat), .B1(new_n731), .B2(new_n704), .ZN(new_n747));
  OR2_X1    g546(.A1(new_n706), .A2(G43gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n722), .B2(new_n748), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(new_n731), .B2(new_n621), .ZN(new_n752));
  INV_X1    g551(.A(new_n621), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n729), .A2(KEYINPUT109), .A3(new_n753), .A4(new_n730), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n752), .A2(new_n228), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT107), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n722), .A2(new_n756), .ZN(new_n757));
  OAI211_X1 g556(.A(KEYINPUT107), .B(new_n721), .C1(new_n688), .C2(new_n690), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n711), .A2(new_n228), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n755), .A2(new_n760), .A3(KEYINPUT48), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n228), .B1(new_n731), .B2(new_n711), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT48), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT108), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT108), .ZN(new_n766));
  AOI211_X1 g565(.A(new_n766), .B(KEYINPUT48), .C1(new_n760), .C2(new_n762), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n761), .B1(new_n765), .B2(new_n767), .ZN(G1331gat));
  NAND3_X1  g567(.A1(new_n299), .A2(new_n689), .A3(new_n322), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n769), .B1(new_n636), .B2(new_n668), .ZN(new_n770));
  OR2_X1    g569(.A1(new_n770), .A2(KEYINPUT110), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(KEYINPUT110), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n616), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g575(.A1(new_n773), .A2(new_n637), .ZN(new_n777));
  NOR2_X1   g576(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n778));
  AND2_X1   g577(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(new_n777), .B2(new_n778), .ZN(G1333gat));
  AOI21_X1  g580(.A(new_n263), .B1(new_n774), .B2(new_n667), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n773), .A2(G71gat), .A3(new_n706), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XOR2_X1   g583(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n785));
  XNOR2_X1  g584(.A(new_n784), .B(new_n785), .ZN(G1334gat));
  NOR2_X1   g585(.A1(new_n773), .A2(new_n711), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(new_n264), .ZN(G1335gat));
  INV_X1    g587(.A(new_n298), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(new_n357), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n791), .A2(new_n323), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n729), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(G85gat), .B1(new_n793), .B2(new_n615), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n728), .A2(new_n791), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT51), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n323), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n615), .A2(G85gat), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n794), .B1(new_n800), .B2(new_n801), .ZN(G1336gat));
  NAND2_X1  g601(.A1(new_n797), .A2(new_n798), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n323), .A2(G92gat), .A3(new_n637), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n729), .A2(new_n582), .A3(new_n792), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(G92gat), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n805), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  XOR2_X1   g608(.A(new_n804), .B(KEYINPUT112), .Z(new_n810));
  AOI22_X1  g609(.A1(new_n803), .A2(new_n810), .B1(new_n807), .B2(G92gat), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n809), .B1(new_n811), .B2(new_n806), .ZN(G1337gat));
  OAI21_X1  g611(.A(G99gat), .B1(new_n793), .B2(new_n704), .ZN(new_n813));
  OR2_X1    g612(.A1(new_n706), .A2(G99gat), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n800), .B2(new_n814), .ZN(G1338gat));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n621), .A2(G106gat), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n799), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(G106gat), .B1(new_n793), .B2(new_n621), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT53), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI211_X1 g619(.A(KEYINPUT53), .B(G106gat), .C1(new_n793), .C2(new_n711), .ZN(new_n821));
  NOR2_X1   g620(.A1(KEYINPUT113), .A2(KEYINPUT53), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n822), .B1(new_n799), .B2(new_n817), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n820), .B1(new_n821), .B2(new_n823), .ZN(G1339gat));
  NOR2_X1   g623(.A1(new_n306), .A2(new_n308), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n312), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(KEYINPUT54), .A3(new_n310), .ZN(new_n827));
  XNOR2_X1  g626(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n311), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n827), .A2(new_n829), .A3(KEYINPUT55), .A4(new_n318), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n827), .A2(new_n829), .A3(new_n318), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n319), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n347), .A2(new_n352), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n354), .A2(new_n355), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n830), .B(new_n833), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n332), .B1(new_n329), .B2(new_n330), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n343), .A2(new_n328), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n841), .A2(G229gat), .A3(G233gat), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n839), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  AOI22_X1  g642(.A1(new_n843), .A2(new_n351), .B1(new_n354), .B2(new_n355), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n322), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n260), .B1(new_n836), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n258), .A3(new_n256), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n833), .A2(new_n830), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT116), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n831), .A2(new_n832), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n852), .A2(new_n320), .A3(new_n830), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n260), .A2(new_n853), .A3(new_n844), .ZN(new_n854));
  AOI22_X1  g653(.A1(new_n853), .A2(new_n357), .B1(new_n844), .B2(new_n322), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n851), .B(new_n854), .C1(new_n855), .C2(new_n260), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n850), .A2(new_n856), .A3(new_n298), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n687), .A2(new_n689), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n582), .A2(new_n615), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n712), .A2(new_n706), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n862), .A2(new_n411), .A3(new_n689), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n615), .B1(new_n857), .B2(new_n858), .ZN(new_n864));
  AND4_X1   g663(.A1(new_n637), .A2(new_n864), .A3(new_n553), .A4(new_n622), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n357), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n863), .B1(new_n866), .B2(new_n411), .ZN(G1340gat));
  NAND4_X1  g666(.A1(new_n865), .A2(new_n434), .A3(new_n435), .A4(new_n322), .ZN(new_n868));
  OAI21_X1  g667(.A(G120gat), .B1(new_n862), .B2(new_n323), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1341gat));
  INV_X1    g669(.A(G127gat), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n865), .A2(new_n871), .A3(new_n789), .ZN(new_n872));
  OAI21_X1  g671(.A(G127gat), .B1(new_n862), .B2(new_n298), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(G1342gat));
  NAND4_X1  g673(.A1(new_n865), .A2(new_n422), .A3(new_n424), .A4(new_n260), .ZN(new_n875));
  XOR2_X1   g674(.A(new_n875), .B(KEYINPUT56), .Z(new_n876));
  OAI21_X1  g675(.A(G134gat), .B1(new_n862), .B2(new_n259), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1343gat));
  NAND2_X1  g677(.A1(new_n704), .A2(new_n753), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(new_n582), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n880), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n881), .A2(G141gat), .A3(new_n689), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n882), .A2(KEYINPUT58), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n704), .A2(new_n860), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n298), .B1(new_n846), .B2(new_n849), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n858), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n712), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n884), .B1(new_n887), .B2(KEYINPUT57), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n621), .B1(new_n857), .B2(new_n858), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT117), .B1(new_n892), .B2(new_n689), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(G141gat), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n892), .A2(KEYINPUT117), .A3(new_n689), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n883), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n892), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n487), .B1(new_n897), .B2(new_n357), .ZN(new_n898));
  OAI21_X1  g697(.A(KEYINPUT58), .B1(new_n898), .B2(new_n882), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n896), .A2(new_n899), .ZN(G1344gat));
  INV_X1    g699(.A(new_n881), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(new_n488), .A3(new_n322), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n889), .A2(KEYINPUT57), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT57), .B1(new_n886), .B2(new_n712), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n906), .A2(new_n704), .A3(new_n322), .A4(new_n860), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n903), .B1(new_n907), .B2(G148gat), .ZN(new_n908));
  AOI211_X1 g707(.A(KEYINPUT59), .B(new_n488), .C1(new_n897), .C2(new_n322), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n902), .B1(new_n908), .B2(new_n909), .ZN(G1345gat));
  OAI21_X1  g709(.A(G155gat), .B1(new_n892), .B2(new_n298), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n881), .A2(G155gat), .A3(new_n298), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  XOR2_X1   g713(.A(new_n914), .B(KEYINPUT118), .Z(G1346gat));
  OAI21_X1  g714(.A(G162gat), .B1(new_n892), .B2(new_n259), .ZN(new_n916));
  OR3_X1    g715(.A1(new_n881), .A2(G162gat), .A3(new_n259), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1347gat));
  AOI21_X1  g717(.A(new_n616), .B1(new_n857), .B2(new_n858), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n553), .A2(new_n582), .A3(new_n622), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n921), .A2(new_n357), .A3(new_n389), .A4(new_n390), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT119), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n637), .A2(new_n616), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n859), .A2(new_n861), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT120), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT120), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n859), .A2(new_n927), .A3(new_n861), .A4(new_n924), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(G169gat), .B1(new_n929), .B2(new_n689), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n923), .A2(new_n930), .ZN(G1348gat));
  OAI21_X1  g730(.A(G176gat), .B1(new_n929), .B2(new_n323), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n921), .A2(new_n378), .A3(new_n322), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1349gat));
  NAND3_X1  g733(.A1(new_n926), .A2(new_n789), .A3(new_n928), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G183gat), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n789), .A2(new_n374), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n919), .A2(new_n920), .A3(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT121), .B1(new_n940), .B2(KEYINPUT60), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n938), .B1(new_n935), .B2(G183gat), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT121), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT60), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT122), .ZN(new_n946));
  AND4_X1   g745(.A1(new_n946), .A2(new_n936), .A3(new_n944), .A4(new_n939), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n946), .B1(new_n942), .B2(new_n944), .ZN(new_n948));
  OAI22_X1  g747(.A1(new_n941), .A2(new_n945), .B1(new_n947), .B2(new_n948), .ZN(G1350gat));
  OAI21_X1  g748(.A(G190gat), .B1(new_n929), .B2(new_n259), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT123), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT123), .ZN(new_n952));
  OAI211_X1 g751(.A(new_n952), .B(G190gat), .C1(new_n929), .C2(new_n259), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n951), .A2(KEYINPUT61), .A3(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n950), .A2(KEYINPUT123), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n921), .A2(new_n370), .A3(new_n260), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n954), .A2(new_n956), .A3(new_n957), .ZN(G1351gat));
  NOR2_X1   g757(.A1(new_n879), .A2(new_n637), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT124), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n919), .A2(new_n960), .ZN(new_n961));
  OR3_X1    g760(.A1(new_n961), .A2(G197gat), .A3(new_n689), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n704), .A2(new_n924), .ZN(new_n963));
  INV_X1    g762(.A(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n906), .A2(new_n357), .A3(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(G197gat), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n965), .A2(new_n966), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n962), .B1(new_n968), .B2(new_n969), .ZN(G1352gat));
  NOR3_X1   g769(.A1(new_n961), .A2(G204gat), .A3(new_n323), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT126), .ZN(new_n972));
  OR2_X1    g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n971), .A2(new_n972), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n906), .A2(new_n322), .A3(new_n964), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n978), .A2(G204gat), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n973), .A2(new_n974), .A3(KEYINPUT62), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n977), .A2(new_n979), .A3(new_n980), .ZN(G1353gat));
  NAND3_X1  g780(.A1(new_n906), .A2(new_n789), .A3(new_n964), .ZN(new_n982));
  AND3_X1   g781(.A1(new_n982), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n983));
  AOI21_X1  g782(.A(KEYINPUT63), .B1(new_n982), .B2(G211gat), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n789), .A2(new_n507), .ZN(new_n985));
  OAI22_X1  g784(.A1(new_n983), .A2(new_n984), .B1(new_n961), .B2(new_n985), .ZN(G1354gat));
  AOI21_X1  g785(.A(KEYINPUT127), .B1(new_n906), .B2(new_n964), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n904), .A2(new_n905), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT127), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n988), .A2(new_n989), .A3(new_n963), .ZN(new_n990));
  NOR3_X1   g789(.A1(new_n987), .A2(new_n990), .A3(new_n259), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n260), .A2(new_n508), .ZN(new_n992));
  OAI22_X1  g791(.A1(new_n991), .A2(new_n508), .B1(new_n961), .B2(new_n992), .ZN(G1355gat));
endmodule


