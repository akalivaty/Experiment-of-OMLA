//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT84), .ZN(new_n189));
  INV_X1    g003(.A(G113), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G116), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n190), .B1(new_n192), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G116), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n194), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(new_n191), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT2), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(new_n190), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT66), .B1(KEYINPUT2), .B2(G113), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n204), .A2(new_n205), .B1(KEYINPUT2), .B2(G113), .ZN(new_n206));
  AOI22_X1  g020(.A1(new_n196), .A2(new_n201), .B1(new_n206), .B2(new_n200), .ZN(new_n207));
  OR2_X1    g021(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n208));
  INV_X1    g022(.A(G107), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G104), .ZN(new_n210));
  AND2_X1   g024(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n208), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G101), .ZN(new_n213));
  INV_X1    g027(.A(G104), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G107), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n214), .A2(G107), .ZN(new_n216));
  NOR2_X1   g030(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n212), .A2(new_n213), .A3(new_n215), .A4(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT80), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n209), .A2(G104), .ZN(new_n221));
  OAI21_X1  g035(.A(G101), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n219), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n220), .B1(new_n219), .B2(new_n222), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n207), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n215), .B1(new_n208), .B2(new_n210), .ZN(new_n226));
  NAND2_X1  g040(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n217), .B1(new_n216), .B2(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(G101), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(KEYINPUT4), .A3(new_n219), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n204), .A2(new_n205), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n203), .A2(new_n190), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n199), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n206), .A2(new_n200), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT4), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n236), .B(G101), .C1(new_n226), .C2(new_n228), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n230), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n225), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT6), .ZN(new_n240));
  XNOR2_X1  g054(.A(G110), .B(G122), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n225), .A2(new_n238), .A3(new_n241), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT6), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n241), .B1(new_n225), .B2(new_n238), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n189), .B(new_n243), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n246), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n248), .A2(KEYINPUT84), .A3(KEYINPUT6), .A4(new_n244), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G146), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G143), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT1), .ZN(new_n253));
  INV_X1    g067(.A(G143), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n254), .A2(G146), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n251), .A2(G143), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n253), .B(G128), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n254), .A2(G146), .ZN(new_n258));
  INV_X1    g072(.A(G128), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n252), .B(new_n258), .C1(KEYINPUT1), .C2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT85), .ZN(new_n262));
  INV_X1    g076(.A(G125), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  AND2_X1   g078(.A1(KEYINPUT0), .A2(G128), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n252), .A2(new_n258), .A3(new_n265), .ZN(new_n266));
  OR2_X1    g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  NAND2_X1  g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(G143), .B(G146), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n266), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n264), .B1(new_n263), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n262), .B1(new_n261), .B2(new_n263), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G224), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(G953), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  NOR3_X1   g093(.A1(new_n273), .A2(new_n277), .A3(new_n274), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n250), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G902), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT7), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n277), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n275), .A2(new_n286), .ZN(new_n287));
  XOR2_X1   g101(.A(new_n241), .B(KEYINPUT8), .Z(new_n288));
  NAND2_X1  g102(.A1(new_n219), .A2(new_n222), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n288), .B1(new_n207), .B2(new_n289), .ZN(new_n290));
  OR2_X1    g104(.A1(new_n196), .A2(KEYINPUT86), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n196), .A2(KEYINPUT86), .B1(KEYINPUT5), .B2(new_n200), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n291), .A2(new_n292), .B1(new_n206), .B2(new_n200), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n290), .B1(new_n293), .B2(new_n289), .ZN(new_n294));
  OAI22_X1  g108(.A1(new_n273), .A2(new_n274), .B1(new_n285), .B2(new_n277), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n287), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n244), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n284), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G210), .B1(G237), .B2(G902), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n283), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n300), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n281), .B1(new_n247), .B2(new_n249), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n302), .B1(new_n303), .B2(new_n298), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n188), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G134), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n254), .A2(G128), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n259), .A2(G143), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n307), .B1(KEYINPUT13), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT13), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n310), .B1(new_n259), .B2(G143), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n306), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT91), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n312), .B(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n308), .A2(new_n307), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n306), .ZN(new_n316));
  XNOR2_X1  g130(.A(G116), .B(G122), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n317), .A2(new_n209), .ZN(new_n318));
  INV_X1    g132(.A(new_n317), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(G107), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n314), .B(new_n316), .C1(new_n318), .C2(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n315), .B(new_n306), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n197), .A2(KEYINPUT14), .A3(G122), .ZN(new_n323));
  OAI211_X1 g137(.A(G107), .B(new_n323), .C1(new_n319), .C2(KEYINPUT14), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n322), .B(new_n324), .C1(G107), .C2(new_n319), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT9), .B(G234), .ZN(new_n326));
  INV_X1    g140(.A(G217), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n326), .A2(new_n327), .A3(G953), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n321), .A2(new_n325), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT92), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT92), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n321), .A2(new_n331), .A3(new_n325), .A4(new_n328), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n321), .A2(new_n325), .ZN(new_n333));
  INV_X1    g147(.A(new_n328), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n330), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n284), .ZN(new_n337));
  INV_X1    g151(.A(G478), .ZN(new_n338));
  NOR2_X1   g152(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n338), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n342), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n344), .B1(new_n336), .B2(new_n284), .ZN(new_n345));
  INV_X1    g159(.A(G952), .ZN(new_n346));
  AOI211_X1 g160(.A(G953), .B(new_n346), .C1(G234), .C2(G237), .ZN(new_n347));
  AND2_X1   g161(.A1(KEYINPUT67), .A2(G953), .ZN(new_n348));
  NOR2_X1   g162(.A1(KEYINPUT67), .A2(G953), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n284), .B1(G234), .B2(G237), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n353), .B(KEYINPUT94), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT21), .B(G898), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n347), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NOR3_X1   g170(.A1(new_n343), .A2(new_n345), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT90), .ZN(new_n358));
  NOR2_X1   g172(.A1(G475), .A2(G902), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n349), .ZN(new_n361));
  INV_X1    g175(.A(G237), .ZN(new_n362));
  NAND2_X1  g176(.A1(KEYINPUT67), .A2(G953), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n361), .A2(G214), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n254), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n350), .A2(G143), .A3(G214), .A4(new_n362), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(KEYINPUT18), .A3(G131), .ZN(new_n368));
  INV_X1    g182(.A(G140), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G125), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n263), .A2(G140), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G146), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n370), .A2(new_n371), .A3(new_n251), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(KEYINPUT18), .A2(G131), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n365), .A2(new_n366), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n368), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT19), .B1(new_n370), .B2(new_n371), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n370), .A2(new_n371), .A3(KEYINPUT19), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(KEYINPUT87), .A3(new_n251), .ZN(new_n383));
  INV_X1    g197(.A(new_n381), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n251), .B1(new_n384), .B2(new_n379), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT87), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n370), .A2(new_n371), .A3(KEYINPUT73), .A4(KEYINPUT16), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n370), .A2(new_n371), .A3(KEYINPUT16), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT73), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n390), .B1(new_n370), .B2(KEYINPUT16), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n388), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G146), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n383), .A2(new_n387), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G131), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n365), .A2(new_n366), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n395), .B1(new_n365), .B2(new_n366), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n378), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(G113), .B(G122), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(new_n214), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n399), .A2(KEYINPUT88), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(KEYINPUT88), .B1(new_n399), .B2(new_n402), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n251), .B(new_n388), .C1(new_n389), .C2(new_n391), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT74), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n393), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  OR3_X1    g222(.A1(new_n392), .A2(new_n407), .A3(G146), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OR2_X1    g224(.A1(new_n396), .A2(new_n397), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n410), .B1(new_n411), .B2(KEYINPUT17), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n397), .A2(KEYINPUT17), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(KEYINPUT89), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n401), .B(new_n378), .C1(new_n412), .C2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n360), .B1(new_n405), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT20), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n358), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n399), .A2(new_n402), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT88), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n399), .A2(KEYINPUT88), .A3(new_n402), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n415), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n359), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(KEYINPUT90), .A3(KEYINPUT20), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n423), .A2(new_n417), .A3(new_n359), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n418), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n378), .B1(new_n412), .B2(new_n414), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n402), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n415), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n284), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G475), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n305), .A2(new_n357), .A3(new_n427), .A4(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT10), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n261), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n435), .B1(new_n223), .B2(new_n224), .ZN(new_n436));
  OAI21_X1  g250(.A(KEYINPUT11), .B1(new_n306), .B2(G137), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT11), .ZN(new_n438));
  INV_X1    g252(.A(G137), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n439), .A3(G134), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT65), .B1(new_n439), .B2(G134), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT65), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(new_n306), .A3(G137), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n441), .A2(new_n395), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n442), .A2(new_n444), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n395), .B1(new_n447), .B2(new_n441), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n434), .B1(new_n289), .B2(new_n261), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n230), .A2(new_n272), .A3(new_n237), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n436), .A2(new_n449), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n350), .A2(G227), .ZN(new_n453));
  XOR2_X1   g267(.A(G110), .B(G140), .Z(new_n454));
  XNOR2_X1  g268(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G131), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n445), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n289), .A2(new_n261), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n219), .A2(new_n222), .B1(new_n257), .B2(new_n260), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(KEYINPUT12), .B1(new_n461), .B2(KEYINPUT81), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n464), .B(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n458), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n436), .A2(new_n450), .A3(new_n451), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n461), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n469), .A2(new_n452), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n467), .B1(new_n470), .B2(new_n456), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT82), .ZN(new_n472));
  INV_X1    g286(.A(G469), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n471), .A2(new_n472), .A3(new_n473), .A4(new_n284), .ZN(new_n474));
  OR2_X1    g288(.A1(new_n464), .A2(new_n465), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n464), .A2(new_n465), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n457), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n456), .B1(new_n469), .B2(new_n452), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n473), .B(new_n284), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT82), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n456), .B1(new_n466), .B2(new_n452), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n482), .B1(new_n458), .B2(new_n469), .ZN(new_n483));
  OAI21_X1  g297(.A(G469), .B1(new_n483), .B2(G902), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(G221), .B1(new_n326), .B2(G902), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OR2_X1    g301(.A1(new_n433), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n271), .B1(new_n460), .B2(new_n445), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n306), .A2(G137), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n439), .A2(G134), .ZN(new_n491));
  OAI21_X1  g305(.A(G131), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AND4_X1   g306(.A1(new_n445), .A2(new_n260), .A3(new_n257), .A4(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n235), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT70), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n272), .B1(new_n446), .B2(new_n448), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n233), .A2(new_n234), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n445), .A2(new_n260), .A3(new_n257), .A4(new_n492), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n494), .A2(new_n495), .A3(new_n499), .ZN(new_n500));
  OAI211_X1 g314(.A(KEYINPUT70), .B(new_n235), .C1(new_n489), .C2(new_n493), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(KEYINPUT28), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT28), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n350), .A2(G210), .A3(new_n362), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT27), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT27), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n350), .A2(new_n507), .A3(G210), .A4(new_n362), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT26), .B(G101), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n506), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n509), .B1(new_n506), .B2(new_n508), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n502), .A2(KEYINPUT29), .A3(new_n504), .A4(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n496), .A2(KEYINPUT30), .A3(new_n498), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT64), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n266), .B(new_n515), .C1(new_n269), .C2(new_n270), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n268), .B(new_n267), .C1(new_n255), .C2(new_n256), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n515), .B1(new_n518), .B2(new_n266), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n445), .A2(new_n492), .ZN(new_n521));
  INV_X1    g335(.A(new_n261), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n520), .A2(new_n461), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n235), .B(new_n514), .C1(new_n523), .C2(KEYINPUT30), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n512), .B1(new_n524), .B2(new_n499), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n271), .A2(KEYINPUT64), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n516), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n498), .B1(new_n449), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n235), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT28), .A4(new_n498), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n504), .A2(new_n529), .A3(new_n512), .A4(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT29), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n513), .B(new_n284), .C1(new_n525), .C2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT71), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n534), .A2(new_n535), .A3(G472), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n535), .B1(new_n534), .B2(G472), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n529), .A2(new_n530), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n512), .B1(new_n539), .B2(new_n504), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n499), .A2(new_n512), .A3(KEYINPUT68), .ZN(new_n541));
  AOI21_X1  g355(.A(KEYINPUT68), .B1(new_n499), .B2(new_n512), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n524), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT31), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n524), .B(KEYINPUT31), .C1(new_n541), .C2(new_n542), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n540), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(G472), .A2(G902), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT69), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT32), .ZN(new_n551));
  INV_X1    g365(.A(new_n540), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n499), .A2(new_n512), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT68), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n499), .A2(new_n512), .A3(KEYINPUT68), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT31), .B1(new_n557), .B2(new_n524), .ZN(new_n558));
  INV_X1    g372(.A(new_n546), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n552), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n551), .B1(new_n560), .B2(new_n548), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n547), .A2(KEYINPUT32), .A3(new_n549), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n550), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI211_X1 g377(.A(KEYINPUT69), .B(new_n551), .C1(new_n547), .C2(new_n549), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n538), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n327), .B1(G234), .B2(new_n284), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n350), .A2(G221), .A3(G234), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(KEYINPUT76), .ZN(new_n569));
  XOR2_X1   g383(.A(KEYINPUT22), .B(G137), .Z(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  XOR2_X1   g386(.A(G119), .B(G128), .Z(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT24), .B(G110), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(KEYINPUT72), .B1(new_n193), .B2(G128), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n576), .A2(KEYINPUT23), .B1(new_n193), .B2(G128), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(KEYINPUT23), .B2(new_n576), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n575), .B1(new_n578), .B2(G110), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n408), .A2(new_n409), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT75), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT75), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n408), .A2(new_n409), .A3(new_n582), .A4(new_n579), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n573), .A2(new_n574), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n585), .B1(new_n578), .B2(G110), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(new_n374), .A3(new_n393), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n572), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n587), .ZN(new_n589));
  AOI211_X1 g403(.A(new_n589), .B(new_n571), .C1(new_n581), .C2(new_n583), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n284), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT25), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g407(.A(KEYINPUT25), .B(new_n284), .C1(new_n588), .C2(new_n590), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n567), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n566), .A2(G902), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n588), .ZN(new_n598));
  INV_X1    g412(.A(new_n590), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT77), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(KEYINPUT77), .B1(new_n588), .B2(new_n590), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n597), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n595), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(KEYINPUT78), .B1(new_n565), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n537), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n534), .A2(new_n535), .A3(G472), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n560), .A2(new_n551), .A3(new_n548), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT32), .B1(new_n547), .B2(new_n549), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n560), .A2(new_n548), .ZN(new_n612));
  AOI22_X1  g426(.A1(new_n610), .A2(new_n611), .B1(new_n612), .B2(KEYINPUT69), .ZN(new_n613));
  INV_X1    g427(.A(new_n564), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n609), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT78), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n616), .A3(new_n604), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n488), .B1(new_n606), .B2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(new_n213), .ZN(G3));
  INV_X1    g433(.A(KEYINPUT96), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n301), .A2(KEYINPUT95), .A3(new_n304), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n187), .B1(new_n301), .B2(KEYINPUT95), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n356), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n303), .A2(new_n302), .A3(new_n298), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT95), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n188), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n301), .A2(KEYINPUT95), .A3(new_n304), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(new_n628), .A3(KEYINPUT96), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT33), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n630), .B1(new_n333), .B2(new_n334), .ZN(new_n631));
  AOI22_X1  g445(.A1(new_n336), .A2(new_n630), .B1(new_n329), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n338), .A2(G902), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT97), .B(G478), .Z(new_n634));
  AOI22_X1  g448(.A1(new_n632), .A2(new_n633), .B1(new_n337), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n427), .B2(new_n432), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n623), .A2(new_n624), .A3(new_n629), .A4(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n486), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n639), .B1(new_n481), .B2(new_n484), .ZN(new_n640));
  OAI21_X1  g454(.A(G472), .B1(new_n547), .B2(G902), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n612), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n640), .A2(new_n604), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n638), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT98), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT34), .B(G104), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  NAND3_X1  g462(.A1(new_n416), .A2(KEYINPUT99), .A3(new_n417), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT99), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n426), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n418), .A2(new_n649), .A3(new_n425), .A4(new_n651), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n652), .A2(new_n432), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n337), .B(new_n342), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n653), .A2(KEYINPUT100), .A3(new_n654), .A4(new_n624), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n627), .A2(new_n628), .A3(KEYINPUT96), .ZN(new_n656));
  AOI21_X1  g470(.A(KEYINPUT96), .B1(new_n627), .B2(new_n628), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n652), .A2(new_n432), .A3(new_n654), .A4(new_n624), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT100), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n655), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n640), .A2(new_n604), .A3(new_n643), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT35), .B(G107), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  NAND2_X1  g480(.A1(new_n584), .A2(new_n587), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n572), .A2(KEYINPUT36), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n597), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n612), .B(new_n641), .C1(new_n595), .C2(new_n670), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n433), .A2(new_n487), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT37), .B(G110), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G12));
  NOR2_X1   g488(.A1(new_n595), .A2(new_n670), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n615), .A2(new_n640), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(G900), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n354), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n679), .A2(new_n347), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n653), .A2(new_n654), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n623), .A2(new_n629), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n677), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n259), .ZN(G30));
  XOR2_X1   g499(.A(new_n680), .B(KEYINPUT39), .Z(new_n686));
  NAND2_X1  g500(.A1(new_n640), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(new_n687), .B(KEYINPUT40), .Z(new_n688));
  INV_X1    g502(.A(G472), .ZN(new_n689));
  INV_X1    g503(.A(new_n512), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n500), .A2(new_n501), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n543), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n689), .B1(new_n692), .B2(new_n284), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n563), .B2(new_n564), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n304), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(new_n625), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n697), .B(KEYINPUT38), .Z(new_n698));
  NAND2_X1  g512(.A1(new_n427), .A2(new_n432), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n654), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n700), .A2(new_n676), .A3(new_n188), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n688), .A2(new_n695), .A3(new_n698), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G143), .ZN(G45));
  NOR2_X1   g517(.A1(new_n565), .A2(new_n675), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n636), .A2(new_n681), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n704), .A2(new_n706), .A3(new_n640), .A4(new_n658), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G146), .ZN(G48));
  NAND2_X1  g522(.A1(new_n471), .A2(new_n284), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(G469), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n481), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n711), .A2(new_n639), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n615), .A2(new_n604), .A3(new_n712), .ZN(new_n713));
  OR2_X1    g527(.A1(new_n713), .A2(new_n637), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT41), .B(G113), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  NOR2_X1   g530(.A1(new_n662), .A2(new_n713), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT101), .B(G116), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G18));
  INV_X1    g533(.A(KEYINPUT103), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n623), .A2(new_n629), .A3(new_n712), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT102), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n623), .A2(new_n712), .A3(KEYINPUT102), .A4(new_n629), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n432), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT90), .B1(new_n424), .B2(KEYINPUT20), .ZN(new_n727));
  AOI211_X1 g541(.A(new_n358), .B(new_n417), .C1(new_n423), .C2(new_n359), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n726), .B1(new_n729), .B2(new_n426), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n615), .A2(new_n730), .A3(new_n357), .A4(new_n676), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n720), .B1(new_n725), .B2(new_n732), .ZN(new_n733));
  AOI211_X1 g547(.A(KEYINPUT103), .B(new_n731), .C1(new_n723), .C2(new_n724), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n193), .ZN(G21));
  NAND4_X1  g550(.A1(new_n623), .A2(new_n699), .A3(new_n654), .A4(new_n629), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n545), .A2(new_n546), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n502), .A2(new_n504), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n690), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n549), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT104), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n641), .A2(new_n742), .ZN(new_n743));
  OAI211_X1 g557(.A(KEYINPUT104), .B(G472), .C1(new_n547), .C2(G902), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n741), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n712), .A2(new_n745), .A3(new_n624), .A4(new_n604), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n737), .A2(new_n746), .ZN(new_n747));
  XOR2_X1   g561(.A(new_n747), .B(G122), .Z(G24));
  NAND4_X1  g562(.A1(new_n676), .A2(new_n636), .A3(new_n745), .A4(new_n681), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n749), .B1(new_n723), .B2(new_n724), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(new_n263), .ZN(G27));
  NAND2_X1  g565(.A1(new_n484), .A2(KEYINPUT105), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n473), .A2(KEYINPUT105), .A3(G902), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n483), .A2(new_n753), .ZN(new_n754));
  AOI22_X1  g568(.A1(new_n752), .A2(new_n754), .B1(new_n474), .B2(new_n480), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n696), .A2(new_n625), .A3(new_n188), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n755), .A2(new_n757), .A3(new_n639), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n565), .A2(new_n605), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n705), .A2(KEYINPUT42), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n610), .A2(new_n611), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n762), .A2(KEYINPUT106), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(KEYINPUT106), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n609), .A3(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n758), .A2(new_n706), .A3(new_n765), .A4(new_n604), .ZN(new_n766));
  AOI22_X1  g580(.A1(new_n760), .A2(new_n761), .B1(new_n766), .B2(KEYINPUT42), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G131), .ZN(G33));
  AND3_X1   g582(.A1(new_n653), .A2(new_n654), .A3(new_n681), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n769), .A2(new_n758), .A3(new_n759), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G134), .ZN(G36));
  OR2_X1    g585(.A1(new_n483), .A2(KEYINPUT45), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n483), .A2(KEYINPUT45), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(G469), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(G469), .A2(G902), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT46), .ZN(new_n777));
  AOI22_X1  g591(.A1(new_n776), .A2(new_n777), .B1(new_n474), .B2(new_n480), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n778), .B1(new_n777), .B2(new_n776), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n779), .A2(new_n486), .A3(new_n686), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n699), .A2(new_n635), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT43), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n782), .A2(new_n642), .A3(new_n676), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n756), .B(new_n780), .C1(new_n783), .C2(KEYINPUT44), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n783), .A2(KEYINPUT44), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(new_n439), .ZN(G39));
  NOR4_X1   g601(.A1(new_n705), .A2(new_n615), .A3(new_n604), .A4(new_n757), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n779), .A2(KEYINPUT47), .A3(new_n486), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT47), .B1(new_n779), .B2(new_n486), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G140), .ZN(G42));
  AND2_X1   g606(.A1(new_n782), .A2(new_n347), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n757), .A2(new_n639), .A3(new_n711), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n765), .A2(new_n604), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XOR2_X1   g612(.A(KEYINPUT115), .B(KEYINPUT48), .Z(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n794), .A2(new_n347), .A3(new_n604), .A4(new_n694), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AOI211_X1 g616(.A(new_n346), .B(G953), .C1(new_n802), .C2(new_n636), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n796), .A2(KEYINPUT115), .A3(KEYINPUT48), .A4(new_n797), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n793), .A2(new_n604), .A3(new_n745), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n725), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n800), .A2(new_n803), .A3(new_n804), .A4(new_n806), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n807), .B(KEYINPUT116), .Z(new_n808));
  NOR2_X1   g622(.A1(new_n698), .A2(new_n187), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n805), .A2(new_n712), .A3(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT50), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n802), .A2(new_n730), .A3(new_n635), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n676), .A2(new_n745), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n812), .B1(new_n795), .B2(new_n813), .ZN(new_n814));
  OR2_X1    g628(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n789), .A2(new_n790), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n711), .A2(new_n486), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n805), .B(new_n756), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT51), .ZN(new_n819));
  XOR2_X1   g633(.A(new_n818), .B(KEYINPUT114), .Z(new_n820));
  NOR2_X1   g634(.A1(new_n815), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n822));
  OAI221_X1 g636(.A(new_n808), .B1(new_n815), .B2(new_n819), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n677), .A2(new_n683), .ZN(new_n825));
  INV_X1    g639(.A(new_n737), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n486), .B1(new_n680), .B2(KEYINPUT110), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n827), .B1(KEYINPUT110), .B2(new_n680), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n675), .A2(new_n828), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n694), .A2(new_n829), .A3(new_n755), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n825), .A2(new_n706), .B1(new_n826), .B2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n684), .ZN(new_n832));
  INV_X1    g646(.A(new_n749), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT102), .B1(new_n658), .B2(new_n712), .ZN(new_n834));
  INV_X1    g648(.A(new_n724), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n831), .A2(new_n832), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n831), .A2(new_n836), .A3(KEYINPUT52), .A4(new_n832), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI22_X1  g655(.A1(new_n637), .A2(new_n713), .B1(new_n737), .B2(new_n746), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n717), .A2(new_n842), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n767), .B(new_n843), .C1(new_n734), .C2(new_n733), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n654), .A2(new_n680), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n653), .A2(new_n756), .A3(new_n846), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n677), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n833), .A2(new_n758), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n770), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT108), .ZN(new_n851));
  AOI211_X1 g665(.A(new_n356), .B(new_n188), .C1(new_n301), .C2(new_n304), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT107), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n730), .A2(new_n852), .A3(new_n853), .A4(new_n654), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n427), .A2(new_n654), .A3(new_n432), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n305), .A2(new_n624), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT107), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n854), .A2(new_n857), .A3(new_n644), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n644), .A2(new_n636), .A3(new_n852), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n433), .A2(new_n487), .ZN(new_n860));
  INV_X1    g674(.A(new_n671), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n858), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n851), .B1(new_n863), .B2(new_n618), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n565), .A2(KEYINPUT78), .A3(new_n605), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n616), .B1(new_n615), .B2(new_n604), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n860), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n635), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n699), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n856), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n644), .A2(new_n870), .B1(new_n860), .B2(new_n861), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n867), .A2(KEYINPUT108), .A3(new_n871), .A4(new_n858), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n850), .B1(new_n864), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n841), .A2(new_n845), .A3(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT53), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n864), .A2(new_n872), .ZN(new_n877));
  INV_X1    g691(.A(new_n850), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n877), .A2(KEYINPUT53), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(new_n844), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT109), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n836), .A2(new_n832), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT109), .B1(new_n750), .B2(new_n684), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n826), .A2(new_n830), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n884), .A2(KEYINPUT52), .A3(new_n707), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n882), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n839), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT111), .B1(new_n880), .B2(new_n887), .ZN(new_n888));
  AOI211_X1 g702(.A(new_n875), .B(new_n850), .C1(new_n864), .C2(new_n872), .ZN(new_n889));
  AND4_X1   g703(.A1(KEYINPUT111), .A2(new_n887), .A3(new_n845), .A4(new_n889), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n824), .B(new_n876), .C1(new_n888), .C2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT112), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n874), .A2(KEYINPUT53), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n887), .A2(new_n845), .A3(new_n875), .A4(new_n873), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n893), .A2(KEYINPUT54), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n887), .A2(new_n845), .A3(new_n889), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT111), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n880), .A2(KEYINPUT111), .A3(new_n887), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT112), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n900), .A2(new_n901), .A3(new_n824), .A4(new_n876), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n892), .A2(new_n895), .A3(new_n902), .ZN(new_n903));
  OAI22_X1  g717(.A1(new_n823), .A2(new_n903), .B1(G952), .B2(G953), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n711), .B(KEYINPUT49), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n730), .A2(new_n486), .A3(new_n187), .A4(new_n868), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n698), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n907), .A2(new_n604), .A3(new_n694), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n904), .A2(new_n908), .ZN(G75));
  INV_X1    g723(.A(KEYINPUT56), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n900), .A2(new_n876), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(G902), .ZN(new_n912));
  INV_X1    g726(.A(G210), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n250), .A2(new_n282), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n915), .A2(new_n303), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT55), .Z(new_n917));
  AND2_X1   g731(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n914), .A2(new_n917), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n350), .A2(G952), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(G51));
  AOI21_X1  g735(.A(new_n824), .B1(new_n900), .B2(new_n876), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n891), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n775), .B(KEYINPUT57), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n471), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n912), .A2(new_n774), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n920), .B1(new_n927), .B2(new_n928), .ZN(G54));
  INV_X1    g743(.A(KEYINPUT117), .ZN(new_n930));
  AND2_X1   g744(.A1(KEYINPUT58), .A2(G475), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n911), .A2(G902), .A3(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n423), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n920), .B1(new_n932), .B2(new_n933), .ZN(new_n935));
  AOI22_X1  g749(.A1(new_n898), .A2(new_n899), .B1(new_n875), .B2(new_n874), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(new_n284), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n937), .A2(KEYINPUT117), .A3(new_n423), .A4(new_n931), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n934), .A2(new_n935), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(KEYINPUT118), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT118), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n934), .A2(new_n935), .A3(new_n941), .A4(new_n938), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n940), .A2(new_n942), .ZN(G60));
  NAND2_X1  g757(.A1(G478), .A2(G902), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT59), .Z(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n902), .A2(new_n895), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n901), .B1(new_n936), .B2(new_n824), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n632), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n950), .A2(new_n945), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n920), .B1(new_n924), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n951), .A2(KEYINPUT119), .A3(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT119), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n632), .B1(new_n903), .B2(new_n946), .ZN(new_n956));
  INV_X1    g770(.A(new_n891), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n952), .B1(new_n957), .B2(new_n922), .ZN(new_n958));
  INV_X1    g772(.A(new_n920), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n955), .B1(new_n956), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n954), .A2(new_n961), .ZN(G63));
  INV_X1    g776(.A(KEYINPUT61), .ZN(new_n963));
  INV_X1    g777(.A(new_n669), .ZN(new_n964));
  NAND2_X1  g778(.A1(G217), .A2(G902), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT60), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n911), .A2(new_n964), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(KEYINPUT120), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n601), .B(new_n602), .C1(new_n936), .C2(new_n966), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n969), .A2(new_n959), .A3(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n968), .A2(KEYINPUT120), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n963), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n970), .A2(KEYINPUT121), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n970), .A2(KEYINPUT121), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n920), .A2(new_n963), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n974), .A2(new_n968), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n973), .A2(new_n977), .ZN(G66));
  OAI21_X1  g792(.A(G953), .B1(new_n355), .B2(new_n276), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n735), .A2(new_n717), .A3(new_n842), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n980), .A2(new_n877), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n979), .B1(new_n981), .B2(new_n351), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n247), .B(new_n249), .C1(G898), .C2(new_n350), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT122), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n982), .B(new_n984), .ZN(G69));
  AOI21_X1  g799(.A(new_n350), .B1(G227), .B2(G900), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n514), .B1(new_n523), .B2(KEYINPUT30), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(new_n382), .Z(new_n988));
  NAND3_X1  g802(.A1(new_n882), .A2(new_n883), .A3(new_n707), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT123), .Z(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n702), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(KEYINPUT62), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT62), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n990), .A2(new_n993), .A3(new_n702), .ZN(new_n994));
  INV_X1    g808(.A(new_n791), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n606), .A2(new_n617), .ZN(new_n996));
  AOI211_X1 g810(.A(new_n757), .B(new_n687), .C1(new_n869), .C2(new_n855), .ZN(new_n997));
  AOI211_X1 g811(.A(new_n995), .B(new_n786), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n992), .A2(new_n994), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n988), .B1(new_n999), .B2(new_n350), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n351), .A2(G900), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n797), .A2(new_n826), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n780), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1003), .B(KEYINPUT126), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n791), .A2(new_n767), .A3(new_n770), .ZN(new_n1005));
  NOR3_X1   g819(.A1(new_n1004), .A2(new_n786), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n990), .A2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n988), .B(new_n1001), .C1(new_n1007), .C2(new_n351), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n986), .B1(new_n1000), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n986), .B(KEYINPUT125), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT124), .ZN(new_n1012));
  OAI211_X1 g826(.A(new_n1008), .B(new_n1011), .C1(new_n1000), .C2(new_n1012), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n1000), .A2(new_n1012), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1010), .B1(new_n1013), .B2(new_n1014), .ZN(G72));
  NAND3_X1  g829(.A1(new_n524), .A2(new_n499), .A3(new_n690), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n990), .A2(new_n1006), .A3(new_n981), .ZN(new_n1017));
  NAND2_X1  g831(.A1(G472), .A2(G902), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1018), .B(KEYINPUT63), .Z(new_n1019));
  AOI21_X1  g833(.A(new_n1016), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  OR3_X1    g834(.A1(new_n1020), .A2(KEYINPUT127), .A3(new_n920), .ZN(new_n1021));
  OAI21_X1  g835(.A(KEYINPUT127), .B1(new_n1020), .B2(new_n920), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n981), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1019), .B1(new_n999), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n690), .B1(new_n524), .B2(new_n499), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(new_n525), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1028), .A2(new_n543), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n893), .A2(new_n894), .A3(new_n1019), .A4(new_n1029), .ZN(new_n1030));
  AND3_X1   g844(.A1(new_n1023), .A2(new_n1027), .A3(new_n1030), .ZN(G57));
endmodule


