//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1184, new_n1185, new_n1186, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  OAI21_X1  g0007(.A(G50), .B1(G58), .B2(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NOR3_X1   g0010(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G1), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n209), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G116), .A2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n219), .B1(G50), .B2(G226), .ZN(new_n220));
  INV_X1    g0020(.A(G58), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  INV_X1    g0022(.A(G107), .ZN(new_n223));
  INV_X1    g0023(.A(G264), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G68), .ZN(new_n226));
  INV_X1    g0026(.A(G238), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n214), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT64), .ZN(new_n230));
  INV_X1    g0030(.A(KEYINPUT65), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n230), .B1(new_n231), .B2(KEYINPUT1), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n214), .A2(G13), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n235), .B(G250), .C1(G257), .C2(G264), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n236), .A2(KEYINPUT0), .ZN(new_n237));
  OR2_X1    g0037(.A1(new_n236), .A2(KEYINPUT0), .ZN(new_n238));
  AOI211_X1 g0038(.A(new_n211), .B(new_n234), .C1(new_n237), .C2(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G250), .B(G257), .Z(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XOR2_X1   g0048(.A(G50), .B(G58), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n250), .B(new_n253), .Z(G351));
  INV_X1    g0054(.A(new_n210), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G41), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT3), .B(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n222), .A2(G1698), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n259), .B(new_n260), .C1(G226), .C2(G1698), .ZN(new_n261));
  INV_X1    g0061(.A(G97), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n258), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT69), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n212), .B1(G41), .B2(G45), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n258), .A2(KEYINPUT66), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(KEYINPUT66), .B1(new_n258), .B2(new_n267), .ZN(new_n270));
  NOR3_X1   g0070(.A1(new_n269), .A2(new_n270), .A3(new_n227), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n266), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n270), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G238), .A3(new_n268), .ZN(new_n276));
  INV_X1    g0076(.A(new_n273), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(KEYINPUT69), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n265), .B1(new_n274), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  AOI211_X1 g0082(.A(new_n280), .B(new_n265), .C1(new_n274), .C2(new_n278), .ZN(new_n283));
  OAI21_X1  g0083(.A(G169), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(KEYINPUT72), .A2(KEYINPUT14), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n274), .A2(new_n278), .ZN(new_n288));
  INV_X1    g0088(.A(new_n265), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT71), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(new_n291), .A3(KEYINPUT13), .ZN(new_n292));
  INV_X1    g0092(.A(new_n283), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT13), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT71), .B1(new_n279), .B2(new_n294), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n292), .A2(new_n293), .A3(new_n295), .A4(G179), .ZN(new_n296));
  NAND2_X1  g0096(.A1(KEYINPUT72), .A2(KEYINPUT14), .ZN(new_n297));
  OAI211_X1 g0097(.A(G169), .B(new_n285), .C1(new_n282), .C2(new_n283), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n287), .A2(new_n296), .A3(new_n297), .A4(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n210), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n301), .B1(new_n212), .B2(G20), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT68), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT12), .ZN(new_n306));
  OAI21_X1  g0106(.A(G68), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n212), .A2(G13), .A3(G20), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n308), .B(KEYINPUT68), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n226), .A2(KEYINPUT12), .ZN(new_n311));
  OAI221_X1 g0111(.A(new_n307), .B1(KEYINPUT12), .B2(new_n309), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n209), .A2(new_n256), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n209), .A2(G33), .ZN(new_n314));
  INV_X1    g0114(.A(G77), .ZN(new_n315));
  OAI22_X1  g0115(.A1(new_n313), .A2(new_n202), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n209), .A2(G68), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n301), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  XOR2_X1   g0118(.A(new_n318), .B(KEYINPUT11), .Z(new_n319));
  NOR2_X1   g0119(.A1(new_n312), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n299), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G1698), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n259), .A2(G232), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n259), .A2(G1698), .ZN(new_n325));
  OAI221_X1 g0125(.A(new_n324), .B1(new_n223), .B2(new_n259), .C1(new_n325), .C2(new_n227), .ZN(new_n326));
  INV_X1    g0126(.A(new_n258), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n273), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n269), .A2(new_n270), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G244), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G169), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XOR2_X1   g0133(.A(KEYINPUT8), .B(G58), .Z(new_n334));
  INV_X1    g0134(.A(new_n313), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n334), .A2(new_n335), .B1(G20), .B2(G77), .ZN(new_n336));
  XOR2_X1   g0136(.A(KEYINPUT15), .B(G87), .Z(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n336), .B1(new_n314), .B2(new_n338), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n301), .A2(new_n339), .B1(new_n305), .B2(G77), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(G77), .B2(new_n310), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n333), .B(new_n341), .C1(G179), .C2(new_n331), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n322), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n302), .A2(G50), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n309), .A2(new_n202), .ZN(new_n345));
  NAND2_X1  g0145(.A1(KEYINPUT67), .A2(G58), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT8), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n346), .B(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G150), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n348), .A2(new_n314), .B1(new_n349), .B2(new_n313), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n350), .B1(G20), .B2(new_n203), .ZN(new_n351));
  INV_X1    g0151(.A(new_n301), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n344), .B(new_n345), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n353), .B(KEYINPUT9), .ZN(new_n354));
  NOR2_X1   g0154(.A1(G222), .A2(G1698), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n323), .A2(G223), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n259), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n357), .B(new_n327), .C1(G77), .C2(new_n259), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n277), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n359), .B1(new_n329), .B2(G226), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G190), .ZN(new_n361));
  INV_X1    g0161(.A(G200), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n354), .B(new_n361), .C1(new_n362), .C2(new_n360), .ZN(new_n363));
  XNOR2_X1  g0163(.A(new_n363), .B(KEYINPUT10), .ZN(new_n364));
  OR2_X1    g0164(.A1(new_n360), .A2(G169), .ZN(new_n365));
  INV_X1    g0165(.A(G179), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n360), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n365), .A2(new_n353), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  OR2_X1    g0169(.A1(new_n343), .A2(new_n369), .ZN(new_n370));
  OR2_X1    g0170(.A1(new_n323), .A2(G226), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n259), .B(new_n371), .C1(G223), .C2(G1698), .ZN(new_n372));
  NAND2_X1  g0172(.A1(G33), .A2(G87), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n258), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n258), .A2(G232), .A3(new_n267), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NOR3_X1   g0176(.A1(new_n374), .A2(new_n376), .A3(new_n273), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT75), .ZN(new_n379));
  NOR4_X1   g0179(.A1(new_n374), .A2(new_n376), .A3(KEYINPUT75), .A4(new_n273), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  OAI22_X1  g0182(.A1(new_n382), .A2(G169), .B1(G179), .B2(new_n378), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n348), .A2(new_n309), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n303), .B2(new_n348), .ZN(new_n385));
  XNOR2_X1  g0185(.A(G58), .B(G68), .ZN(new_n386));
  AOI22_X1  g0186(.A1(G20), .A2(new_n386), .B1(new_n335), .B2(G159), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT3), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G33), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n392), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT73), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n259), .A2(KEYINPUT73), .ZN(new_n396));
  AOI21_X1  g0196(.A(G20), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n393), .B1(new_n397), .B2(KEYINPUT7), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n388), .B1(new_n398), .B2(G68), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n352), .B1(new_n399), .B2(KEYINPUT16), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT7), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n259), .B2(G20), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n393), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G68), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT74), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT74), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n403), .A2(new_n406), .A3(G68), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n405), .A2(new_n387), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT16), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n385), .B1(new_n400), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT18), .ZN(new_n412));
  NOR3_X1   g0212(.A1(new_n383), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n400), .A2(new_n410), .ZN(new_n414));
  INV_X1    g0214(.A(new_n385), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT75), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n377), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n418), .A2(new_n380), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n419), .A2(new_n332), .B1(new_n366), .B2(new_n377), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT18), .B1(new_n416), .B2(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n413), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n379), .A2(new_n362), .A3(new_n381), .ZN(new_n424));
  INV_X1    g0224(.A(G190), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n377), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n411), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT17), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n427), .A2(new_n411), .A3(KEYINPUT17), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n341), .B1(new_n331), .B2(G200), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n425), .B2(new_n331), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n292), .A2(new_n293), .A3(new_n295), .A4(G190), .ZN(new_n436));
  OAI21_X1  g0236(.A(G200), .B1(new_n282), .B2(new_n283), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n320), .A3(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n423), .A2(new_n433), .A3(new_n435), .A4(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n370), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n212), .A2(G33), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n310), .A2(G116), .A3(new_n352), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G283), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n443), .B(new_n209), .C1(G33), .C2(new_n262), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n444), .B(new_n301), .C1(new_n209), .C2(G116), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT20), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n445), .A2(new_n446), .ZN(new_n448));
  OAI221_X1 g0248(.A(new_n442), .B1(G116), .B2(new_n310), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT77), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n257), .A2(KEYINPUT5), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n212), .A2(G45), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n257), .A2(KEYINPUT5), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT5), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G41), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n457), .A2(KEYINPUT77), .A3(new_n212), .A4(G45), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n454), .A2(new_n455), .A3(new_n458), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n459), .A2(new_n258), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G270), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n259), .A2(G257), .A3(new_n323), .ZN(new_n462));
  INV_X1    g0262(.A(G303), .ZN(new_n463));
  OAI221_X1 g0263(.A(new_n462), .B1(new_n463), .B2(new_n259), .C1(new_n325), .C2(new_n224), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n327), .ZN(new_n465));
  OR3_X1    g0265(.A1(new_n459), .A2(new_n272), .A3(new_n327), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n461), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NOR3_X1   g0267(.A1(new_n450), .A2(new_n467), .A3(new_n366), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(G200), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n470), .B(new_n450), .C1(new_n425), .C2(new_n467), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n467), .A2(G169), .A3(new_n449), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(KEYINPUT81), .A3(KEYINPUT21), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT21), .B1(new_n472), .B2(KEYINPUT81), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n469), .B(new_n471), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n310), .A2(new_n337), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n259), .A2(new_n209), .A3(G68), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT19), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n479), .B1(new_n314), .B2(new_n262), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT79), .B(G87), .ZN(new_n481));
  OAI22_X1  g0281(.A1(new_n481), .A2(new_n206), .B1(G20), .B2(new_n263), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n478), .B(new_n480), .C1(new_n482), .C2(new_n479), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n477), .B1(new_n483), .B2(new_n301), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n352), .A2(new_n308), .A3(new_n441), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n337), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT80), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n484), .A2(KEYINPUT80), .A3(new_n487), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n389), .A2(new_n391), .A3(G238), .A4(new_n323), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT78), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT78), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n259), .A2(new_n494), .A3(G238), .A4(new_n323), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n259), .A2(G244), .A3(G1698), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G116), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n327), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n258), .A2(G250), .A3(new_n453), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n453), .A2(new_n272), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n500), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G169), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n500), .A2(G179), .A3(new_n501), .A4(new_n503), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n490), .A2(new_n491), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n476), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n259), .A2(new_n209), .A3(G87), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT22), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT22), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n259), .A2(new_n511), .A3(new_n209), .A4(G87), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n223), .A2(G20), .ZN(new_n514));
  INV_X1    g0314(.A(G116), .ZN(new_n515));
  OAI22_X1  g0315(.A1(KEYINPUT23), .A2(new_n514), .B1(new_n314), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(KEYINPUT23), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT82), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT82), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n514), .A2(new_n519), .A3(KEYINPUT23), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n516), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n513), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT24), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n513), .A2(KEYINPUT24), .A3(new_n521), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n524), .A2(new_n301), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n486), .A2(G107), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n309), .A2(KEYINPUT25), .A3(new_n223), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT83), .ZN(new_n529));
  AOI21_X1  g0329(.A(KEYINPUT25), .B1(new_n309), .B2(new_n223), .ZN(new_n530));
  XOR2_X1   g0330(.A(new_n529), .B(new_n530), .Z(new_n531));
  NAND3_X1  g0331(.A1(new_n526), .A2(new_n527), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n459), .A2(G264), .A3(new_n258), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT84), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT84), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n459), .A2(new_n535), .A3(G264), .A4(new_n258), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n389), .A2(new_n391), .A3(G250), .A4(new_n323), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n389), .A2(new_n391), .A3(G257), .A4(G1698), .ZN(new_n539));
  INV_X1    g0339(.A(G294), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n538), .B(new_n539), .C1(new_n256), .C2(new_n540), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n541), .A2(new_n327), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n537), .A2(new_n466), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT85), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n542), .B1(new_n534), .B2(new_n536), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n547), .A2(KEYINPUT85), .A3(new_n466), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n332), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n544), .A2(new_n366), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n532), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(KEYINPUT86), .ZN(new_n552));
  AND4_X1   g0352(.A1(KEYINPUT85), .A2(new_n537), .A3(new_n466), .A4(new_n543), .ZN(new_n553));
  AOI21_X1  g0353(.A(KEYINPUT85), .B1(new_n547), .B2(new_n466), .ZN(new_n554));
  OAI21_X1  g0354(.A(G169), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n550), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT86), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n558), .A3(new_n532), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n552), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n546), .A2(new_n425), .A3(new_n548), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n544), .A2(new_n362), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n532), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n460), .A2(G257), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n259), .A2(G244), .A3(new_n323), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT76), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT4), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n567), .B1(new_n565), .B2(new_n566), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n443), .B1(new_n325), .B2(new_n218), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n466), .B(new_n564), .C1(new_n571), .C2(new_n258), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n332), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n223), .A2(KEYINPUT6), .A3(G97), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n262), .A2(new_n223), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n575), .A2(new_n205), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n574), .B1(new_n576), .B2(KEYINPUT6), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n577), .A2(G20), .B1(G77), .B2(new_n335), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n403), .A2(G107), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n352), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n485), .A2(new_n262), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n308), .A2(G97), .ZN(new_n582));
  OR3_X1    g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n565), .A2(new_n566), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT4), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n327), .B1(new_n587), .B2(new_n570), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n588), .A2(new_n366), .A3(new_n466), .A4(new_n564), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n573), .A2(new_n583), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n572), .A2(G200), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n588), .A2(G190), .A3(new_n466), .A4(new_n564), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n485), .A2(new_n217), .ZN(new_n596));
  AOI211_X1 g0396(.A(new_n596), .B(new_n477), .C1(new_n483), .C2(new_n301), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n493), .A2(new_n495), .A3(new_n498), .A4(new_n497), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n502), .B1(new_n598), .B2(new_n327), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n599), .A2(G190), .A3(new_n501), .ZN(new_n600));
  INV_X1    g0400(.A(new_n501), .ZN(new_n601));
  AOI211_X1 g0401(.A(new_n601), .B(new_n502), .C1(new_n598), .C2(new_n327), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n597), .B(new_n600), .C1(new_n362), .C2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n563), .A2(new_n595), .A3(new_n604), .ZN(new_n605));
  AND4_X1   g0405(.A1(new_n440), .A2(new_n508), .A3(new_n560), .A4(new_n605), .ZN(G372));
  INV_X1    g0406(.A(new_n368), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n343), .A2(new_n433), .A3(new_n438), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n608), .A2(new_n423), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT88), .ZN(new_n610));
  OR2_X1    g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n364), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n612), .B1(new_n609), .B2(new_n610), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n607), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n440), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT87), .ZN(new_n616));
  INV_X1    g0416(.A(new_n506), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n332), .B1(new_n599), .B2(new_n501), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n506), .B(KEYINPUT87), .C1(new_n602), .C2(new_n332), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n490), .A2(new_n491), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n604), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT26), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n573), .A2(new_n583), .A3(new_n589), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n603), .A2(new_n573), .A3(new_n583), .A4(new_n589), .ZN(new_n627));
  OAI21_X1  g0427(.A(KEYINPUT26), .B1(new_n627), .B2(new_n507), .ZN(new_n628));
  INV_X1    g0428(.A(new_n620), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT87), .B1(new_n505), .B2(new_n506), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n622), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n626), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n475), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n468), .B1(new_n633), .B2(new_n473), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n634), .A2(new_n551), .B1(new_n622), .B2(new_n621), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n632), .B1(new_n635), .B2(new_n605), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n614), .B1(new_n615), .B2(new_n636), .ZN(G369));
  INV_X1    g0437(.A(new_n563), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n526), .A2(new_n527), .A3(new_n531), .ZN(new_n639));
  INV_X1    g0439(.A(G13), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(G20), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n212), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(G213), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(G343), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n560), .B(new_n638), .C1(new_n639), .C2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n557), .A2(new_n532), .A3(new_n647), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n450), .A2(new_n648), .ZN(new_n652));
  MUX2_X1   g0452(.A(new_n476), .B(new_n634), .S(new_n652), .Z(new_n653));
  INV_X1    g0453(.A(G330), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n634), .A2(new_n647), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n560), .A2(new_n638), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n557), .A2(new_n532), .A3(new_n648), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n656), .A2(new_n660), .ZN(G399));
  INV_X1    g0461(.A(new_n235), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(G41), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G1), .ZN(new_n665));
  OR3_X1    g0465(.A1(new_n481), .A2(G116), .A3(new_n206), .ZN(new_n666));
  OAI22_X1  g0466(.A1(new_n665), .A2(new_n666), .B1(new_n208), .B2(new_n664), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT28), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n560), .A2(new_n508), .A3(new_n605), .A4(new_n648), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT31), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n544), .A2(new_n467), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT30), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n617), .A2(new_n564), .A3(new_n588), .ZN(new_n673));
  OR3_X1    g0473(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n672), .B1(new_n671), .B2(new_n673), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n602), .B1(new_n547), .B2(new_n466), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n676), .A2(new_n366), .A3(new_n467), .A4(new_n572), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n674), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n647), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n670), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n675), .A2(KEYINPUT89), .A3(new_n677), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n674), .ZN(new_n682));
  AOI21_X1  g0482(.A(KEYINPUT89), .B1(new_n675), .B2(new_n677), .ZN(new_n683));
  OAI211_X1 g0483(.A(KEYINPUT31), .B(new_n647), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n654), .B1(new_n680), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n558), .B1(new_n557), .B2(new_n532), .ZN(new_n686));
  AOI211_X1 g0486(.A(KEYINPUT86), .B(new_n639), .C1(new_n555), .C2(new_n556), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n634), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT93), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n560), .A2(KEYINPUT93), .A3(new_n634), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(new_n605), .A3(new_n691), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n631), .A2(new_n625), .A3(KEYINPUT26), .A4(new_n603), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT91), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n623), .A2(KEYINPUT91), .A3(KEYINPUT26), .A4(new_n625), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n624), .B1(new_n627), .B2(new_n507), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT92), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT92), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n699), .B(new_n624), .C1(new_n627), .C2(new_n507), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n695), .A2(new_n696), .A3(new_n698), .A4(new_n700), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n701), .A2(new_n631), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n647), .B1(new_n692), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT29), .ZN(new_n704));
  INV_X1    g0504(.A(new_n632), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n635), .A2(new_n605), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n647), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT90), .B1(new_n707), .B2(KEYINPUT29), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT90), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n709), .B(new_n710), .C1(new_n636), .C2(new_n647), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n685), .B1(new_n704), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n668), .B1(new_n713), .B2(G1), .ZN(G364));
  INV_X1    g0514(.A(new_n655), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n665), .B1(G45), .B2(new_n641), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n653), .A2(new_n654), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n715), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NOR3_X1   g0519(.A1(G13), .A2(G20), .A3(G33), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT98), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n653), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n210), .B1(G20), .B2(new_n332), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n209), .A2(G190), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G179), .A2(G200), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(G159), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT32), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n209), .A2(new_n366), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G190), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n362), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n728), .B1(new_n732), .B2(new_n202), .ZN(new_n733));
  INV_X1    g0533(.A(new_n729), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n734), .A2(new_n362), .A3(G190), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n726), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G159), .ZN(new_n738));
  OAI22_X1  g0538(.A1(new_n736), .A2(new_n226), .B1(KEYINPUT32), .B2(new_n738), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n734), .A2(G190), .A3(G200), .ZN(new_n740));
  AOI211_X1 g0540(.A(new_n733), .B(new_n739), .C1(G77), .C2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n362), .A2(G179), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n724), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G107), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n742), .A2(G20), .A3(G190), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n481), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n209), .B1(new_n725), .B2(G190), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n749), .A2(KEYINPUT97), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(KEYINPUT97), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n748), .B1(new_n752), .B2(new_n262), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n730), .A2(G200), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n753), .B1(G58), .B2(new_n754), .ZN(new_n755));
  AND4_X1   g0555(.A1(new_n259), .A2(new_n741), .A3(new_n745), .A4(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G283), .ZN(new_n757));
  INV_X1    g0557(.A(new_n740), .ZN(new_n758));
  INV_X1    g0558(.A(G311), .ZN(new_n759));
  OAI221_X1 g0559(.A(new_n392), .B1(new_n743), .B2(new_n757), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n747), .A2(G303), .B1(new_n737), .B2(G329), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n754), .A2(G322), .ZN(new_n762));
  XOR2_X1   g0562(.A(KEYINPUT33), .B(G317), .Z(new_n763));
  OAI211_X1 g0563(.A(new_n761), .B(new_n762), .C1(new_n736), .C2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G326), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n732), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n752), .A2(new_n540), .ZN(new_n767));
  NOR4_X1   g0567(.A1(new_n760), .A2(new_n764), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n723), .B1(new_n756), .B2(new_n768), .ZN(new_n769));
  XOR2_X1   g0569(.A(G355), .B(KEYINPUT94), .Z(new_n770));
  NOR2_X1   g0570(.A1(new_n662), .A2(new_n392), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n770), .A2(new_n771), .B1(new_n515), .B2(new_n662), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n395), .A2(new_n396), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n662), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(G45), .B2(new_n208), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n776), .B(KEYINPUT96), .Z(new_n777));
  NAND2_X1  g0577(.A1(new_n250), .A2(G45), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT95), .Z(new_n779));
  OAI21_X1  g0579(.A(new_n772), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n723), .A2(new_n720), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n722), .A2(new_n769), .A3(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n719), .B1(new_n717), .B2(new_n783), .ZN(G396));
  NAND2_X1  g0584(.A1(new_n341), .A2(new_n647), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n435), .A2(new_n785), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n786), .A2(new_n342), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n342), .A2(new_n647), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n707), .B(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(new_n685), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n717), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G13), .A2(G33), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(new_n787), .B2(new_n788), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G159), .A2(new_n740), .B1(new_n754), .B2(G143), .ZN(new_n795));
  INV_X1    g0595(.A(G137), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n795), .B1(new_n796), .B2(new_n732), .C1(new_n349), .C2(new_n736), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT34), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n774), .B1(new_n221), .B2(new_n752), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n797), .A2(new_n798), .B1(G68), .B2(new_n744), .ZN(new_n800));
  INV_X1    g0600(.A(G132), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n801), .B2(new_n726), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n799), .B(new_n802), .C1(G50), .C2(new_n747), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n731), .A2(G303), .B1(new_n744), .B2(G87), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n804), .B1(new_n736), .B2(new_n757), .C1(new_n262), .C2(new_n752), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT99), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n392), .B1(new_n746), .B2(new_n223), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n806), .A2(new_n807), .B1(new_n740), .B2(G116), .ZN(new_n808));
  INV_X1    g0608(.A(new_n754), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n808), .B1(new_n806), .B2(new_n807), .C1(new_n540), .C2(new_n809), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n805), .B(new_n810), .C1(G311), .C2(new_n737), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n723), .B1(new_n803), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n723), .A2(new_n793), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n315), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n794), .A2(new_n716), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n792), .A2(new_n815), .ZN(G384));
  INV_X1    g0616(.A(new_n679), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n817), .A2(KEYINPUT31), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n680), .A2(new_n819), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n440), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT40), .ZN(new_n822));
  INV_X1    g0622(.A(new_n645), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n400), .B1(KEYINPUT16), .B2(new_n399), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n415), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n823), .B(new_n825), .C1(new_n422), .C2(new_n432), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n383), .A2(new_n645), .B1(new_n415), .B2(new_n824), .ZN(new_n827));
  INV_X1    g0627(.A(new_n428), .ZN(new_n828));
  OAI21_X1  g0628(.A(KEYINPUT37), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n416), .A2(new_n420), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n416), .A2(new_n823), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT37), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n830), .A2(new_n831), .A3(new_n832), .A4(new_n428), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  AND3_X1   g0634(.A1(new_n826), .A2(KEYINPUT38), .A3(new_n834), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n416), .B(new_n823), .C1(new_n422), .C2(new_n432), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n830), .A2(new_n831), .A3(new_n428), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(KEYINPUT37), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n833), .ZN(new_n839));
  AOI21_X1  g0639(.A(KEYINPUT38), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n835), .A2(new_n840), .ZN(new_n841));
  AND3_X1   g0641(.A1(new_n299), .A2(new_n321), .A3(new_n648), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n321), .A2(new_n647), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n299), .A2(new_n321), .B1(new_n438), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n817), .B1(new_n669), .B2(KEYINPUT31), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n789), .B(new_n845), .C1(new_n846), .C2(new_n818), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT102), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n841), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(KEYINPUT40), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n820), .A2(new_n789), .A3(new_n845), .A4(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n822), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT38), .B1(new_n826), .B2(new_n834), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n835), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n821), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(G330), .B1(new_n852), .B2(new_n856), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n821), .A2(G330), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n857), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n788), .B1(new_n707), .B2(new_n789), .ZN(new_n863));
  INV_X1    g0663(.A(new_n845), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n854), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n423), .B2(new_n823), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT39), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n841), .A2(KEYINPUT101), .A3(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT101), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n854), .B2(KEYINPUT39), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n835), .A2(new_n840), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n872), .A2(KEYINPUT39), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n869), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n867), .B1(new_n874), .B2(new_n842), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n862), .B(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n704), .A2(new_n712), .A3(new_n440), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n614), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n876), .B(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n212), .B2(new_n641), .ZN(new_n880));
  OAI211_X1 g0680(.A(G20), .B(new_n255), .C1(new_n577), .C2(KEYINPUT35), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n515), .B(new_n881), .C1(KEYINPUT35), .C2(new_n577), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n882), .B(KEYINPUT36), .Z(new_n883));
  INV_X1    g0683(.A(KEYINPUT100), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n226), .B2(G50), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n202), .A2(KEYINPUT100), .A3(G68), .ZN(new_n886));
  OAI21_X1  g0686(.A(G77), .B1(new_n221), .B2(new_n226), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n885), .B(new_n886), .C1(new_n887), .C2(new_n208), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n888), .A2(G1), .A3(new_n640), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n880), .A2(new_n883), .A3(new_n889), .ZN(G367));
  NOR2_X1   g0690(.A1(new_n752), .A2(new_n226), .ZN(new_n891));
  OAI22_X1  g0691(.A1(new_n746), .A2(new_n221), .B1(new_n726), .B2(new_n796), .ZN(new_n892));
  INV_X1    g0692(.A(G143), .ZN(new_n893));
  OAI221_X1 g0693(.A(new_n259), .B1(new_n892), .B2(KEYINPUT108), .C1(new_n893), .C2(new_n732), .ZN(new_n894));
  AOI211_X1 g0694(.A(new_n891), .B(new_n894), .C1(KEYINPUT108), .C2(new_n892), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n743), .A2(new_n315), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n740), .B2(G50), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  OAI221_X1 g0698(.A(new_n898), .B1(new_n349), .B2(new_n809), .C1(new_n727), .C2(new_n736), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n743), .A2(new_n262), .ZN(new_n900));
  INV_X1    g0700(.A(new_n752), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n746), .A2(new_n515), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n901), .A2(G107), .B1(KEYINPUT46), .B2(new_n902), .ZN(new_n903));
  OAI221_X1 g0703(.A(new_n903), .B1(KEYINPUT46), .B2(new_n902), .C1(new_n759), .C2(new_n732), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n758), .A2(new_n757), .ZN(new_n905));
  XOR2_X1   g0705(.A(KEYINPUT107), .B(G317), .Z(new_n906));
  NOR2_X1   g0706(.A1(new_n906), .A2(new_n726), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n736), .A2(new_n540), .ZN(new_n908));
  NOR4_X1   g0708(.A1(new_n904), .A2(new_n905), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n909), .B(new_n773), .C1(new_n463), .C2(new_n809), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n899), .B1(new_n900), .B2(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT47), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n723), .ZN(new_n913));
  INV_X1    g0713(.A(new_n775), .ZN(new_n914));
  OAI221_X1 g0714(.A(new_n781), .B1(new_n235), .B2(new_n338), .C1(new_n914), .C2(new_n246), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n913), .A2(new_n716), .A3(new_n915), .ZN(new_n916));
  OR3_X1    g0716(.A1(new_n631), .A2(new_n597), .A3(new_n648), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n623), .B1(new_n597), .B2(new_n648), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n916), .B1(new_n721), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n590), .B(new_n594), .C1(new_n592), .C2(new_n648), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n625), .A2(new_n647), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n660), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT44), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n660), .A2(new_n925), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT45), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n928), .B(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(new_n656), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n658), .B1(new_n651), .B2(new_n657), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n655), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n715), .B(new_n658), .C1(new_n651), .C2(new_n657), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AND3_X1   g0736(.A1(new_n713), .A2(KEYINPUT104), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT104), .B1(new_n713), .B2(new_n936), .ZN(new_n938));
  OAI21_X1  g0738(.A(KEYINPUT105), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n713), .A2(new_n936), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT104), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT105), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n713), .A2(KEYINPUT104), .A3(new_n936), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n932), .A2(new_n939), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n713), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n663), .B(KEYINPUT41), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT106), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT106), .ZN(new_n950));
  INV_X1    g0750(.A(new_n948), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n950), .B(new_n951), .C1(new_n946), .C2(new_n713), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n212), .B1(new_n641), .B2(G45), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NOR3_X1   g0754(.A1(new_n949), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n658), .B1(new_n923), .B2(new_n924), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT42), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n590), .B1(new_n560), .B2(new_n923), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n648), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n919), .B(KEYINPUT43), .Z(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT103), .ZN(new_n963));
  NOR3_X1   g0763(.A1(new_n960), .A2(KEYINPUT43), .A3(new_n919), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n656), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n925), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n965), .B(new_n967), .Z(new_n968));
  OAI21_X1  g0768(.A(new_n922), .B1(new_n955), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(KEYINPUT109), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT109), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n971), .B(new_n922), .C1(new_n955), .C2(new_n968), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(G387));
  NAND2_X1  g0773(.A1(new_n942), .A2(new_n944), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n974), .B(new_n663), .C1(new_n713), .C2(new_n936), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n936), .A2(new_n954), .ZN(new_n976));
  AOI22_X1  g0776(.A1(G303), .A2(new_n740), .B1(new_n731), .B2(G322), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n977), .B1(new_n759), .B2(new_n736), .C1(new_n809), .C2(new_n906), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT48), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n979), .B1(new_n757), .B2(new_n752), .C1(new_n540), .C2(new_n746), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT49), .Z(new_n981));
  OAI221_X1 g0781(.A(new_n773), .B1(new_n515), .B2(new_n743), .C1(new_n765), .C2(new_n726), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT111), .Z(new_n983));
  NOR2_X1   g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n736), .A2(new_n348), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n900), .B(new_n985), .C1(G150), .C2(new_n737), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n226), .B2(new_n758), .C1(new_n727), .C2(new_n732), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n752), .A2(new_n338), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n809), .A2(new_n202), .B1(new_n315), .B2(new_n746), .ZN(new_n989));
  NOR4_X1   g0789(.A1(new_n987), .A2(new_n773), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n723), .B1(new_n984), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n334), .A2(new_n202), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT110), .Z(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT50), .ZN(new_n994));
  INV_X1    g0794(.A(G45), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n226), .B2(new_n315), .ZN(new_n996));
  NOR3_X1   g0796(.A1(new_n994), .A2(new_n666), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n771), .A2(new_n666), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n775), .B1(new_n243), .B2(new_n995), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n235), .A2(G107), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n781), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n649), .A2(new_n650), .A3(new_n721), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n991), .A2(new_n716), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n975), .A2(new_n976), .A3(new_n1004), .ZN(G393));
  XNOR2_X1  g0805(.A(new_n931), .B(new_n966), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1006), .A2(KEYINPUT112), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(KEYINPUT112), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1007), .A2(new_n954), .A3(new_n1008), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(G150), .A2(new_n731), .B1(new_n754), .B2(G159), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT51), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G68), .B2(new_n747), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n735), .A2(G50), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n773), .B1(new_n901), .B2(G77), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n743), .A2(new_n217), .B1(new_n726), .B2(new_n893), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n334), .B2(new_n740), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .A4(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G311), .A2(new_n754), .B1(new_n731), .B2(G317), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT113), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT52), .Z(new_n1020));
  AOI22_X1  g0820(.A1(new_n747), .A2(G283), .B1(new_n737), .B2(G322), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n745), .B1(new_n752), .B2(new_n515), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n259), .B(new_n1022), .C1(G303), .C2(new_n735), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1020), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n758), .A2(new_n540), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1017), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n723), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n781), .B1(new_n262), .B2(new_n235), .C1(new_n914), .C2(new_n253), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n923), .A2(new_n924), .A3(new_n720), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1027), .A2(new_n716), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1009), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1006), .A2(new_n974), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n946), .A2(new_n663), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1031), .A2(new_n1033), .ZN(G390));
  NAND3_X1  g0834(.A1(new_n820), .A2(G330), .A3(new_n789), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n864), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n685), .A2(new_n789), .A3(new_n845), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n787), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n788), .B1(new_n703), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1036), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT115), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1036), .A2(KEYINPUT115), .A3(new_n1037), .A4(new_n1039), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n845), .B1(new_n685), .B2(new_n789), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n847), .A2(new_n654), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1042), .B(new_n1043), .C1(new_n863), .C2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n878), .A2(new_n861), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(KEYINPUT116), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n842), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n872), .B(new_n1051), .C1(new_n1039), .C2(new_n844), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(KEYINPUT114), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n844), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n647), .B(new_n787), .C1(new_n692), .C2(new_n702), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1054), .B1(new_n1055), .B2(new_n788), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT114), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1056), .A2(new_n1057), .A3(new_n872), .A4(new_n1051), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1051), .B1(new_n863), .B2(new_n864), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n869), .B(new_n1059), .C1(new_n871), .C2(new_n873), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1053), .A2(new_n1037), .A3(new_n1058), .A4(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1053), .A2(new_n1060), .A3(new_n1058), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n1045), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1050), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1061), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1065), .A2(new_n1049), .A3(KEYINPUT116), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n663), .A3(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1063), .A2(new_n954), .A3(new_n1061), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT117), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1063), .A2(KEYINPUT117), .A3(new_n954), .A4(new_n1061), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n793), .B(new_n869), .C1(new_n871), .C2(new_n873), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n813), .A2(new_n348), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n743), .A2(new_n226), .B1(new_n726), .B2(new_n540), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n901), .A2(G77), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n259), .B1(new_n747), .B2(G87), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n740), .A2(G97), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n731), .A2(G283), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n1075), .B(new_n1080), .C1(G107), .C2(new_n735), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n754), .A2(G116), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n754), .A2(G132), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n747), .A2(G150), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n1084), .A2(KEYINPUT53), .B1(new_n731), .B2(G128), .ZN(new_n1085));
  INV_X1    g0885(.A(G125), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1085), .B1(new_n202), .B2(new_n743), .C1(new_n1086), .C2(new_n726), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT54), .B(G143), .Z(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n259), .B1(new_n758), .B2(new_n1089), .C1(new_n752), .C2(new_n727), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n736), .A2(new_n796), .B1(new_n1084), .B2(KEYINPUT53), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1087), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1081), .A2(new_n1082), .B1(new_n1083), .B2(new_n1092), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT118), .Z(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n723), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1073), .A2(new_n716), .A3(new_n1074), .A4(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(KEYINPUT119), .B1(new_n1072), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT119), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1096), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1098), .B(new_n1099), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1067), .B1(new_n1097), .B2(new_n1100), .ZN(G378));
  INV_X1    g0901(.A(KEYINPUT55), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n369), .B(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1103), .A2(new_n353), .A3(new_n823), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n369), .B(KEYINPUT55), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n353), .A2(new_n823), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  XOR2_X1   g0907(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1108));
  AND3_X1   g0908(.A1(new_n1104), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1108), .B1(new_n1104), .B2(new_n1107), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n858), .A2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1111), .B(G330), .C1(new_n852), .C2(new_n856), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n875), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1113), .A2(new_n875), .A3(new_n1114), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n954), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1112), .A2(new_n793), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n758), .A2(new_n338), .B1(new_n221), .B2(new_n743), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(G97), .B2(new_n735), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n731), .A2(G116), .B1(new_n747), .B2(G77), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NOR4_X1   g0925(.A1(new_n1125), .A2(G41), .A3(new_n774), .A4(new_n891), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1126), .B1(new_n223), .B2(new_n809), .C1(new_n757), .C2(new_n726), .ZN(new_n1127));
  XOR2_X1   g0927(.A(new_n1127), .B(KEYINPUT58), .Z(new_n1128));
  OAI22_X1  g0928(.A1(new_n736), .A2(new_n801), .B1(new_n732), .B2(new_n1086), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(G137), .B2(new_n740), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n901), .A2(G150), .B1(G128), .B2(new_n754), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1130), .B(new_n1131), .C1(new_n746), .C2(new_n1089), .ZN(new_n1132));
  XOR2_X1   g0932(.A(new_n1132), .B(KEYINPUT59), .Z(new_n1133));
  NOR2_X1   g0933(.A1(G33), .A2(G41), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT120), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G124), .B2(new_n737), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1133), .B(new_n1136), .C1(new_n727), .C2(new_n743), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n202), .B(new_n1135), .C1(new_n774), .C2(G41), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n723), .B1(new_n1128), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n813), .A2(new_n202), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1121), .A2(new_n716), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1120), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1063), .A2(new_n1047), .A3(new_n1061), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1117), .A2(new_n1118), .B1(new_n1144), .B2(new_n1048), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n663), .B1(new_n1145), .B2(KEYINPUT57), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT57), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(new_n1144), .B2(new_n1048), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT122), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1117), .A2(new_n1149), .A3(new_n1118), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1115), .A2(KEYINPUT122), .A3(new_n1116), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1148), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1143), .B1(new_n1146), .B2(new_n1152), .ZN(G375));
  AOI211_X1 g0953(.A(new_n896), .B(new_n988), .C1(G283), .C2(new_n754), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n731), .A2(G294), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n746), .A2(new_n262), .B1(new_n726), .B2(new_n463), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT123), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n758), .A2(new_n223), .B1(new_n736), .B2(new_n515), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1158), .A2(new_n259), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1154), .A2(new_n1155), .A3(new_n1157), .A4(new_n1159), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n752), .A2(new_n202), .B1(new_n758), .B2(new_n349), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT124), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n735), .A2(new_n1088), .B1(new_n731), .B2(G132), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(G58), .A2(new_n744), .B1(new_n737), .B2(G128), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n773), .B1(G159), .B2(new_n747), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .A4(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n809), .A2(new_n796), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1160), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1168), .A2(new_n723), .B1(new_n226), .B2(new_n813), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n716), .ZN(new_n1170));
  XOR2_X1   g0970(.A(new_n1170), .B(KEYINPUT125), .Z(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(new_n864), .B2(new_n793), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n1047), .B2(new_n954), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1049), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n948), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1173), .B1(new_n1174), .B2(new_n1175), .ZN(G381));
  INV_X1    g0976(.A(G390), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(G381), .A2(G384), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n970), .A2(new_n972), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(G378), .A2(G375), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(G393), .A2(G396), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1179), .A2(new_n1182), .ZN(G407));
  NAND2_X1  g0983(.A1(new_n1180), .A2(new_n646), .ZN(new_n1184));
  OAI211_X1 g0984(.A(G213), .B(new_n1184), .C1(new_n1179), .C2(new_n1182), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT126), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1185), .B(new_n1186), .ZN(G409));
  NAND2_X1  g0987(.A1(G378), .A2(G375), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1150), .A2(new_n954), .A3(new_n1151), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1144), .A2(new_n1048), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1119), .A2(new_n1190), .A3(new_n948), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n1189), .A2(new_n1142), .A3(new_n1191), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1192), .B(new_n1067), .C1(new_n1097), .C2(new_n1100), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT60), .ZN(new_n1194));
  OR3_X1    g0994(.A1(new_n1047), .A2(new_n1194), .A3(new_n1048), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1194), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1195), .A2(new_n663), .A3(new_n1049), .A4(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n1173), .ZN(new_n1198));
  INV_X1    g0998(.A(G384), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1197), .A2(G384), .A3(new_n1173), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n646), .A2(G213), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1188), .A2(new_n1193), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(KEYINPUT62), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1188), .A2(new_n1193), .A3(new_n1203), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n646), .A2(G213), .A3(G2897), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1200), .A2(new_n1201), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1207), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1206), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT61), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G378), .A2(G375), .B1(G213), .B2(new_n646), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT62), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1213), .A2(new_n1214), .A3(new_n1202), .A4(new_n1193), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1205), .A2(new_n1211), .A3(new_n1212), .A4(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n969), .A2(G390), .ZN(new_n1217));
  XOR2_X1   g1017(.A(G393), .B(G396), .Z(new_n1218));
  OAI211_X1 g1018(.A(new_n1177), .B(new_n922), .C1(new_n955), .C2(new_n968), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n970), .A2(new_n972), .A3(new_n1177), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n1217), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1218), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1220), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1216), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT63), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1204), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT127), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1204), .A2(KEYINPUT127), .A3(new_n1226), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1213), .A2(KEYINPUT63), .A3(new_n1202), .A4(new_n1193), .ZN(new_n1232));
  AOI21_X1  g1032(.A(KEYINPUT61), .B1(new_n1206), .B2(new_n1210), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1218), .B1(new_n1221), .B2(new_n1217), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1232), .B(new_n1233), .C1(new_n1234), .C2(new_n1220), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1225), .B1(new_n1231), .B2(new_n1235), .ZN(G405));
  OR2_X1    g1036(.A1(G378), .A2(G375), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1202), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1237), .A2(new_n1238), .A3(new_n1188), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1238), .B1(new_n1237), .B2(new_n1188), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1224), .A2(new_n1241), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n1234), .A2(new_n1220), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(G402));
endmodule


