//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n584, new_n585, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n627, new_n629, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT66), .Z(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n455), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n455), .A2(G2106), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n458), .A2(KEYINPUT67), .A3(G567), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n463));
  INV_X1    g038(.A(G567), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n463), .B1(new_n457), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n461), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(G319));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n473), .B(KEYINPUT68), .ZN(new_n474));
  OAI21_X1  g049(.A(G2105), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(G137), .B(new_n476), .C1(new_n468), .C2(new_n469), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n476), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  AND3_X1   g054(.A1(new_n477), .A2(new_n479), .A3(KEYINPUT69), .ZN(new_n480));
  AOI21_X1  g055(.A(KEYINPUT69), .B1(new_n477), .B2(new_n479), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n475), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT70), .ZN(G160));
  NOR2_X1   g058(.A1(new_n470), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n470), .A2(new_n476), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n476), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  XNOR2_X1  g066(.A(KEYINPUT3), .B(G2104), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n492), .A2(G126), .A3(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(G114), .B2(new_n476), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n492), .A2(KEYINPUT4), .A3(G138), .A4(new_n476), .ZN(new_n499));
  OAI211_X1 g074(.A(G138), .B(new_n476), .C1(new_n468), .C2(new_n469), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n497), .A2(new_n498), .A3(new_n499), .A4(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n502), .A2(new_n499), .A3(new_n493), .A4(new_n496), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT71), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT72), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT72), .A2(G651), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT6), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n508), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n518), .B1(new_n511), .B2(new_n513), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G88), .ZN(new_n520));
  NAND2_X1  g095(.A1(G75), .A2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G62), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n509), .A2(new_n510), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n515), .A2(new_n520), .A3(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  NAND2_X1  g103(.A1(new_n519), .A2(G89), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT6), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n531));
  INV_X1    g106(.A(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(KEYINPUT72), .A2(G651), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n530), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g110(.A(G51), .B(G543), .C1(new_n535), .C2(new_n512), .ZN(new_n536));
  OR2_X1    g111(.A1(KEYINPUT5), .A2(G543), .ZN(new_n537));
  NAND2_X1  g112(.A1(KEYINPUT5), .A2(G543), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n532), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(KEYINPUT7), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT7), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n542), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n539), .A2(G63), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n529), .A2(new_n536), .A3(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(G168));
  NAND2_X1  g121(.A1(new_n519), .A2(G90), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n514), .A2(G52), .ZN(new_n548));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G64), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n518), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(new_n525), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n547), .A2(new_n548), .A3(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  NAND2_X1  g129(.A1(new_n537), .A2(new_n538), .ZN(new_n555));
  OAI211_X1 g130(.A(G81), .B(new_n555), .C1(new_n535), .C2(new_n512), .ZN(new_n556));
  OAI211_X1 g131(.A(G43), .B(G543), .C1(new_n535), .C2(new_n512), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(new_n537), .B2(new_n538), .ZN(new_n559));
  INV_X1    g134(.A(G68), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(new_n508), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n525), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n556), .A2(new_n557), .A3(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT73), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT73), .A4(new_n562), .ZN(new_n566));
  AND2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  OAI211_X1 g147(.A(G53), .B(G543), .C1(new_n535), .C2(new_n512), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT74), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT9), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n555), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n573), .A2(new_n575), .B1(new_n532), .B2(new_n576), .ZN(new_n577));
  XOR2_X1   g152(.A(KEYINPUT74), .B(KEYINPUT9), .Z(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(new_n514), .B2(G53), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g155(.A(G91), .B(new_n555), .C1(new_n535), .C2(new_n512), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT75), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(G299));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n545), .B(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G286));
  NAND2_X1  g161(.A1(new_n519), .A2(G87), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n514), .A2(G49), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT77), .ZN(new_n589));
  OAI211_X1 g164(.A(new_n589), .B(G651), .C1(new_n555), .C2(G74), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n555), .B2(G74), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(KEYINPUT77), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n587), .A2(new_n588), .A3(new_n590), .A4(new_n592), .ZN(G288));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G61), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n518), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n514), .A2(G48), .B1(new_n596), .B2(new_n525), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n519), .A2(G86), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g175(.A(KEYINPUT78), .B1(new_n519), .B2(G86), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n597), .B1(new_n600), .B2(new_n601), .ZN(G305));
  AOI22_X1  g177(.A1(new_n555), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(new_n524), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT79), .ZN(new_n605));
  AOI22_X1  g180(.A1(G47), .A2(new_n514), .B1(new_n519), .B2(G85), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(G290));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  OR3_X1    g183(.A1(G171), .A2(KEYINPUT80), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(KEYINPUT80), .B1(G171), .B2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n514), .A2(G54), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n518), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G651), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  OAI211_X1 g191(.A(G92), .B(new_n555), .C1(new_n535), .C2(new_n512), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT10), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n519), .A2(KEYINPUT10), .A3(G92), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n616), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n609), .B(new_n610), .C1(G868), .C2(new_n621), .ZN(G284));
  OAI211_X1 g197(.A(new_n609), .B(new_n610), .C1(G868), .C2(new_n621), .ZN(G321));
  NOR2_X1   g198(.A1(G299), .A2(G868), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(G868), .B2(new_n585), .ZN(G297));
  AOI21_X1  g200(.A(new_n624), .B1(G868), .B2(new_n585), .ZN(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n621), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND2_X1  g203(.A1(new_n565), .A2(new_n566), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(new_n608), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n621), .A2(new_n627), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n630), .B1(new_n632), .B2(new_n608), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n492), .A2(new_n478), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2100), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n486), .A2(G123), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT83), .Z(new_n641));
  NAND2_X1  g216(.A1(new_n484), .A2(G135), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT82), .ZN(new_n643));
  OAI21_X1  g218(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n644));
  INV_X1    g219(.A(KEYINPUT84), .ZN(new_n645));
  INV_X1    g220(.A(G111), .ZN(new_n646));
  AOI22_X1  g221(.A1(new_n644), .A2(new_n645), .B1(new_n646), .B2(G2105), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n645), .B2(new_n644), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n641), .A2(new_n643), .A3(new_n648), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n649), .A2(G2096), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(G2096), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n639), .A2(new_n650), .A3(new_n651), .ZN(G156));
  XNOR2_X1  g227(.A(G2427), .B(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2430), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(KEYINPUT14), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1341), .B(G1348), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2451), .B(G2454), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT16), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT85), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n662), .A2(new_n665), .ZN(new_n667));
  AND3_X1   g242(.A1(new_n666), .A2(G14), .A3(new_n667), .ZN(G401));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT86), .ZN(new_n671));
  NOR2_X1   g246(.A1(G2072), .A2(G2078), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n442), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n669), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(KEYINPUT17), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n674), .B1(new_n671), .B2(new_n675), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n669), .B(new_n670), .C1(new_n442), .C2(new_n672), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT18), .Z(new_n678));
  NAND3_X1  g253(.A1(new_n675), .A2(new_n671), .A3(new_n669), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n676), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G2096), .B(G2100), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G227));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  AND2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n686), .A2(new_n687), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n685), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT89), .ZN(new_n694));
  OR3_X1    g269(.A1(new_n685), .A2(new_n688), .A3(new_n692), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n691), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(G229));
  AOI22_X1  g277(.A1(new_n484), .A2(G141), .B1(G105), .B2(new_n478), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n486), .A2(G129), .ZN(new_n704));
  NAND3_X1  g279(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT26), .Z(new_n706));
  NAND3_X1  g281(.A1(new_n703), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT98), .Z(new_n708));
  MUX2_X1   g283(.A(G32), .B(new_n708), .S(G29), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT27), .ZN(new_n710));
  INV_X1    g285(.A(G1996), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G35), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G162), .B2(new_n714), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G2090), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT101), .Z(new_n719));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G20), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT23), .ZN(new_n722));
  INV_X1    g297(.A(G299), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(new_n720), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT102), .B(G1956), .Z(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n712), .A2(new_n713), .A3(new_n719), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT30), .B(G28), .ZN(new_n728));
  OR2_X1    g303(.A1(KEYINPUT31), .A2(G11), .ZN(new_n729));
  NAND2_X1  g304(.A1(KEYINPUT31), .A2(G11), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n728), .A2(new_n714), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n649), .B2(new_n714), .ZN(new_n732));
  AND2_X1   g307(.A1(new_n732), .A2(KEYINPUT99), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n717), .A2(G2090), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT25), .Z(new_n736));
  NAND2_X1  g311(.A1(new_n484), .A2(G139), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n492), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n736), .B(new_n737), .C1(new_n476), .C2(new_n738), .ZN(new_n739));
  MUX2_X1   g314(.A(G33), .B(new_n739), .S(G29), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G2072), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n720), .A2(G21), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G168), .B2(new_n720), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n743), .A2(G1966), .ZN(new_n744));
  NOR4_X1   g319(.A1(new_n733), .A2(new_n734), .A3(new_n741), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n714), .A2(G27), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G164), .B2(new_n714), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT100), .ZN(new_n748));
  INV_X1    g323(.A(G2078), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(new_n749), .ZN(new_n751));
  OAI22_X1  g326(.A1(new_n732), .A2(KEYINPUT99), .B1(G1966), .B2(new_n743), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n720), .A2(G5), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G171), .B2(new_n720), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1961), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n745), .A2(new_n750), .A3(new_n751), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(G160), .A2(G29), .ZN(new_n758));
  INV_X1    g333(.A(G34), .ZN(new_n759));
  AOI21_X1  g334(.A(G29), .B1(new_n759), .B2(KEYINPUT24), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(KEYINPUT24), .B2(new_n759), .ZN(new_n761));
  AOI21_X1  g336(.A(G2084), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n758), .A2(G2084), .A3(new_n761), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n725), .B2(new_n724), .ZN(new_n764));
  NOR4_X1   g339(.A1(new_n727), .A2(new_n757), .A3(new_n762), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n714), .A2(G26), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT28), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n484), .A2(G140), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n486), .A2(G128), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n476), .A2(G116), .ZN(new_n770));
  OAI21_X1  g345(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n768), .B(new_n769), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n772), .A2(KEYINPUT95), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(KEYINPUT95), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n767), .B1(new_n775), .B2(G29), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT96), .ZN(new_n777));
  INV_X1    g352(.A(G2067), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n720), .A2(G4), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n621), .B2(new_n720), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT94), .B(G1348), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n720), .A2(G19), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n567), .B2(new_n720), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(G1341), .Z(new_n786));
  NAND3_X1  g361(.A1(new_n779), .A2(new_n783), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT97), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n765), .A2(new_n788), .ZN(new_n789));
  MUX2_X1   g364(.A(G6), .B(G305), .S(G16), .Z(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT32), .B(G1981), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G16), .A2(G23), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT92), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G288), .B2(new_n720), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT33), .B(G1976), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n720), .A2(G22), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G303), .B2(G16), .ZN(new_n799));
  INV_X1    g374(.A(G1971), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n797), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n792), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT93), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT34), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n714), .A2(G25), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n484), .A2(G131), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n486), .A2(G119), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n476), .A2(G107), .ZN(new_n812));
  OAI21_X1  g387(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n810), .B(new_n811), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n814), .A2(KEYINPUT90), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(KEYINPUT90), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n809), .B1(new_n818), .B2(new_n714), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT35), .B(G1991), .Z(new_n820));
  XOR2_X1   g395(.A(new_n819), .B(new_n820), .Z(new_n821));
  INV_X1    g396(.A(KEYINPUT91), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  MUX2_X1   g399(.A(G24), .B(G290), .S(G16), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1986), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n807), .A2(new_n808), .A3(new_n823), .A4(new_n827), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n828), .A2(KEYINPUT36), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(KEYINPUT36), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n789), .B1(new_n829), .B2(new_n830), .ZN(G311));
  AND2_X1   g406(.A1(new_n828), .A2(KEYINPUT36), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n828), .A2(KEYINPUT36), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n788), .B(new_n765), .C1(new_n832), .C2(new_n833), .ZN(G150));
  OAI211_X1 g409(.A(G55), .B(G543), .C1(new_n535), .C2(new_n512), .ZN(new_n835));
  OAI211_X1 g410(.A(G93), .B(new_n555), .C1(new_n535), .C2(new_n512), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT104), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n835), .A2(new_n836), .A3(KEYINPUT104), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT103), .ZN(new_n841));
  AND2_X1   g416(.A1(G80), .A2(G543), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(new_n555), .B2(G67), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n841), .B1(new_n843), .B2(new_n524), .ZN(new_n844));
  INV_X1    g419(.A(G67), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n518), .A2(new_n845), .ZN(new_n846));
  OAI211_X1 g421(.A(KEYINPUT103), .B(new_n525), .C1(new_n846), .C2(new_n842), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n839), .A2(new_n840), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G860), .ZN(new_n850));
  XOR2_X1   g425(.A(KEYINPUT107), .B(KEYINPUT37), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n621), .A2(G559), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT106), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT38), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT105), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n849), .A2(new_n856), .A3(new_n565), .A4(new_n566), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n839), .A2(new_n848), .A3(new_n563), .A4(new_n840), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n856), .B1(new_n567), .B2(new_n849), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n855), .B(new_n861), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n862), .A2(KEYINPUT39), .ZN(new_n863));
  INV_X1    g438(.A(G860), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n862), .B2(KEYINPUT39), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n852), .B1(new_n863), .B2(new_n865), .ZN(G145));
  XNOR2_X1  g441(.A(new_n708), .B(new_n775), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n484), .A2(G142), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n486), .A2(G130), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n476), .A2(G118), .ZN(new_n870));
  OAI21_X1  g445(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n868), .B(new_n869), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n867), .B(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n817), .B(new_n637), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n739), .B(new_n504), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n873), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(G160), .B(G162), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n649), .ZN(new_n879));
  AOI21_X1  g454(.A(G37), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n880), .B1(new_n879), .B2(new_n877), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g457(.A1(new_n861), .A2(new_n631), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n632), .B1(new_n859), .B2(new_n860), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT41), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n619), .A2(new_n620), .ZN(new_n886));
  AOI22_X1  g461(.A1(new_n514), .A2(G54), .B1(new_n614), .B2(G651), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n576), .A2(new_n532), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n514), .A2(new_n574), .A3(KEYINPUT9), .A4(G53), .ZN(new_n890));
  INV_X1    g465(.A(new_n573), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n889), .B(new_n890), .C1(new_n891), .C2(new_n578), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT75), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n581), .B(new_n893), .ZN(new_n894));
  NOR3_X1   g469(.A1(new_n888), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  AOI22_X1  g470(.A1(new_n580), .A2(new_n582), .B1(new_n886), .B2(new_n887), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n885), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(G299), .A2(new_n888), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n621), .A2(new_n582), .A3(new_n580), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(KEYINPUT41), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n883), .A2(new_n884), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n895), .A2(new_n896), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n904), .B1(new_n883), .B2(new_n884), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT42), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n905), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(new_n908), .A3(new_n902), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(G290), .B(G305), .ZN(new_n911));
  XNOR2_X1  g486(.A(G166), .B(G288), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n911), .B(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n906), .A2(new_n909), .A3(new_n913), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(G868), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n839), .A2(new_n840), .A3(new_n848), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n919), .A2(G868), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(new_n921), .ZN(G295));
  INV_X1    g497(.A(KEYINPUT108), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n923), .B1(new_n918), .B2(new_n921), .ZN(new_n924));
  AOI211_X1 g499(.A(KEYINPUT108), .B(new_n920), .C1(new_n917), .C2(G868), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(G331));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n927));
  NAND2_X1  g502(.A1(G301), .A2(new_n545), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n929), .B1(new_n585), .B2(G171), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n930), .B1(new_n859), .B2(new_n860), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n536), .A2(new_n544), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT76), .B1(new_n932), .B2(new_n529), .ZN(new_n933));
  AND4_X1   g508(.A1(KEYINPUT76), .A2(new_n529), .A3(new_n536), .A4(new_n544), .ZN(new_n934));
  OAI21_X1  g509(.A(G171), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n928), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT105), .B1(new_n919), .B2(new_n629), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n936), .A2(new_n937), .A3(new_n858), .A4(new_n857), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n931), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n901), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n931), .A2(new_n938), .A3(new_n904), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n927), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n927), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n913), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G37), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n931), .A2(new_n938), .A3(new_n904), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n901), .B1(new_n938), .B2(new_n931), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT109), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n951), .A2(new_n914), .A3(new_n944), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT43), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT111), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n941), .A2(new_n942), .ZN(new_n956));
  AOI21_X1  g531(.A(G37), .B1(new_n956), .B2(new_n913), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n952), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n955), .B1(new_n952), .B2(new_n957), .ZN(new_n960));
  OAI221_X1 g535(.A(KEYINPUT44), .B1(new_n948), .B2(new_n954), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n946), .A2(new_n947), .A3(new_n952), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n952), .A2(new_n953), .A3(new_n957), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n962), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI211_X1 g543(.A(KEYINPUT110), .B(KEYINPUT44), .C1(new_n964), .C2(new_n965), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n961), .B1(new_n968), .B2(new_n969), .ZN(G397));
  INV_X1    g545(.A(KEYINPUT118), .ZN(new_n971));
  INV_X1    g546(.A(G1384), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n506), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n971), .B1(new_n973), .B2(KEYINPUT50), .ZN(new_n974));
  AOI21_X1  g549(.A(G1384), .B1(new_n503), .B2(new_n505), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n975), .A2(KEYINPUT118), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT113), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n504), .A2(new_n979), .A3(new_n972), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n979), .B1(new_n504), .B2(new_n972), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT50), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n475), .B(G40), .C1(new_n480), .C2(new_n481), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n983), .A2(KEYINPUT117), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT117), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n504), .A2(new_n972), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(KEYINPUT113), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n976), .B1(new_n989), .B2(new_n980), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n987), .B1(new_n990), .B2(new_n984), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n978), .A2(new_n986), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G1956), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n972), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n996), .A2(new_n984), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(KEYINPUT45), .B2(new_n975), .ZN(new_n998));
  XNOR2_X1  g573(.A(KEYINPUT56), .B(G2072), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n994), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT57), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n723), .A2(KEYINPUT121), .A3(new_n1004), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n1004), .A2(KEYINPUT121), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(KEYINPUT121), .ZN(new_n1007));
  NAND3_X1  g582(.A1(G299), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1003), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1001), .B1(new_n992), .B2(new_n993), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1009), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1010), .A2(KEYINPUT61), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT61), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1016));
  AOI211_X1 g591(.A(new_n1009), .B(new_n1001), .C1(new_n992), .C2(new_n993), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n629), .B1(KEYINPUT123), .B2(KEYINPUT59), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n997), .B(new_n711), .C1(KEYINPUT45), .C2(new_n975), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT122), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n985), .A2(new_n989), .A3(new_n980), .ZN(new_n1022));
  XOR2_X1   g597(.A(KEYINPUT58), .B(G1341), .Z(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1020), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1021), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1019), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n989), .A2(new_n976), .A3(new_n980), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n985), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n975), .A2(new_n976), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n782), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OR2_X1    g608(.A1(new_n1022), .A2(G2067), .ZN(new_n1034));
  OR2_X1    g609(.A1(new_n621), .A2(KEYINPUT60), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n621), .A2(KEYINPUT60), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n1037), .B(KEYINPUT124), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1038), .A2(new_n1033), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI221_X1 g617(.A(new_n1019), .B1(KEYINPUT123), .B2(KEYINPUT59), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1029), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1014), .A2(new_n1018), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n888), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1016), .B1(new_n1013), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(G303), .A2(G8), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1049), .B(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G2090), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n978), .A2(new_n986), .A3(new_n1052), .A4(new_n991), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n998), .A2(new_n800), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1051), .B1(new_n1055), .B2(G8), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n973), .A2(KEYINPUT50), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1057), .A2(new_n1052), .A3(new_n985), .A4(new_n1030), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n1054), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1059), .A2(G8), .A3(new_n1051), .ZN(new_n1060));
  INV_X1    g635(.A(G1976), .ZN(new_n1061));
  OR2_X1    g636(.A1(G288), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT52), .B1(G288), .B2(new_n1061), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1022), .A2(new_n1062), .A3(G8), .A4(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n1064), .B(KEYINPUT115), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1022), .A2(G8), .A3(new_n1062), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT52), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1022), .A2(G8), .ZN(new_n1068));
  INV_X1    g643(.A(G1981), .ZN(new_n1069));
  AOI211_X1 g644(.A(KEYINPUT116), .B(new_n1069), .C1(new_n597), .C2(new_n598), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1069), .B(new_n597), .C1(new_n600), .C2(new_n601), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n514), .A2(G48), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n596), .A2(new_n525), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1073), .A2(new_n598), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1072), .B1(new_n1075), .B2(G1981), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1070), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT49), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1068), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1079), .B1(new_n1078), .B2(new_n1077), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1060), .A2(new_n1065), .A3(new_n1067), .A4(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1056), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n975), .A2(KEYINPUT45), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT45), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n981), .B2(new_n982), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1083), .A2(new_n1085), .A3(new_n985), .ZN(new_n1086));
  INV_X1    g661(.A(G1966), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G2084), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1057), .A2(new_n1089), .A3(new_n985), .A4(new_n1030), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(G168), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(G8), .ZN(new_n1092));
  AOI21_X1  g667(.A(G168), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT51), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT51), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1091), .A2(new_n1095), .A3(G8), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n997), .B(new_n749), .C1(KEYINPUT45), .C2(new_n975), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(G1961), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1100), .A2(G2078), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1083), .A2(new_n1085), .A3(new_n985), .A4(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(G301), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n984), .B(KEYINPUT125), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n988), .A2(new_n1084), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1108), .A2(new_n995), .A3(new_n1105), .A4(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1101), .A2(new_n1103), .A3(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(G171), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1098), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1082), .A2(new_n1097), .A3(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1104), .A2(G301), .A3(new_n1106), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1098), .B1(new_n1111), .B2(G171), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1115), .A2(new_n1116), .A3(KEYINPUT126), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT126), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1114), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1048), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1060), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT63), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1124), .A2(G8), .A3(new_n585), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1122), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1080), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1051), .B1(new_n1059), .B2(G8), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1127), .A2(new_n1128), .A3(KEYINPUT119), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1068), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1071), .A2(new_n1076), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1070), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1132), .A2(new_n1133), .A3(new_n1078), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1067), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT115), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1064), .B(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1059), .A2(G8), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1051), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1130), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1126), .B1(new_n1129), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g722(.A(KEYINPUT120), .B(new_n1126), .C1(new_n1129), .C2(new_n1144), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n1056), .A2(new_n1081), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1123), .B1(new_n1149), .B2(new_n1125), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1071), .ZN(new_n1152));
  NOR2_X1   g727(.A1(G288), .A2(G1976), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1152), .B1(new_n1080), .B2(new_n1153), .ZN(new_n1154));
  OAI22_X1  g729(.A1(new_n1154), .A2(new_n1068), .B1(new_n1127), .B2(new_n1060), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT62), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1094), .A2(new_n1156), .A3(new_n1096), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1157), .A2(new_n1082), .A3(new_n1107), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1097), .A2(KEYINPUT62), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1155), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1121), .A2(new_n1151), .A3(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n817), .B(new_n820), .ZN(new_n1162));
  XOR2_X1   g737(.A(new_n1162), .B(KEYINPUT112), .Z(new_n1163));
  XNOR2_X1  g738(.A(new_n708), .B(new_n711), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n775), .A2(G2067), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n773), .A2(new_n778), .A3(new_n774), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1163), .A2(new_n1168), .ZN(new_n1169));
  XOR2_X1   g744(.A(G290), .B(G1986), .Z(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1109), .A2(new_n984), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1161), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1172), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1169), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT48), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n1175), .A2(G1986), .A3(G290), .ZN(new_n1178));
  XOR2_X1   g753(.A(new_n1178), .B(KEYINPUT127), .Z(new_n1179));
  AOI21_X1  g754(.A(new_n1176), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1180), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1167), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1172), .B1(new_n1182), .B2(new_n708), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1172), .A2(KEYINPUT46), .A3(new_n711), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT46), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1185), .B1(new_n1175), .B2(G1996), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1183), .A2(new_n1184), .A3(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n1187), .B(KEYINPUT47), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n818), .A2(new_n820), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1166), .B1(new_n1168), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1190), .A2(new_n1172), .ZN(new_n1191));
  AND3_X1   g766(.A1(new_n1181), .A2(new_n1188), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1174), .A2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g768(.A1(G229), .A2(G401), .A3(new_n466), .A4(G227), .ZN(new_n1195));
  NAND3_X1  g769(.A1(new_n966), .A2(new_n881), .A3(new_n1195), .ZN(G225));
  INV_X1    g770(.A(G225), .ZN(G308));
endmodule


