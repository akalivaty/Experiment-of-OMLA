//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1263, new_n1264, new_n1265, new_n1267,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1328, new_n1329,
    new_n1330, new_n1331;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  AOI22_X1  g0003(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n204));
  AOI22_X1  g0004(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g0009(.A(new_n203), .B1(new_n206), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT1), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT64), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n212), .B1(new_n203), .B2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G13), .ZN(new_n214));
  NAND4_X1  g0014(.A1(new_n214), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT0), .Z(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(G50), .B1(G58), .B2(G68), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  AOI211_X1 g0023(.A(new_n211), .B(new_n218), .C1(new_n221), .C2(new_n223), .ZN(G361));
  XOR2_X1   g0024(.A(G238), .B(G244), .Z(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT65), .B(G232), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT66), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n229), .B(new_n233), .ZN(G358));
  XNOR2_X1  g0034(.A(G50), .B(G68), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT67), .ZN(new_n236));
  XOR2_X1   g0036(.A(G58), .B(G77), .Z(new_n237));
  XOR2_X1   g0037(.A(new_n236), .B(new_n237), .Z(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G351));
  XNOR2_X1  g0042(.A(KEYINPUT8), .B(G58), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n220), .A2(G33), .ZN(new_n244));
  INV_X1    g0044(.A(G150), .ZN(new_n245));
  NOR2_X1   g0045(.A1(G20), .A2(G33), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  OAI22_X1  g0047(.A1(new_n243), .A2(new_n244), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  NOR2_X1   g0048(.A1(G58), .A2(G68), .ZN(new_n249));
  INV_X1    g0049(.A(G50), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n220), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OR2_X1    g0051(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n219), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT70), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT70), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n253), .A2(new_n256), .A3(new_n219), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n252), .A2(new_n258), .B1(new_n250), .B2(new_n261), .ZN(new_n262));
  AND3_X1   g0062(.A1(new_n255), .A2(new_n260), .A3(new_n257), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n259), .A2(G20), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(G50), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n266), .B(KEYINPUT9), .ZN(new_n267));
  INV_X1    g0067(.A(new_n219), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G223), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT69), .ZN(new_n273));
  AND2_X1   g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n273), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT3), .ZN(new_n279));
  INV_X1    g0079(.A(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(KEYINPUT69), .A3(G1698), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n272), .B1(new_n278), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n277), .ZN(new_n286));
  INV_X1    g0086(.A(G222), .ZN(new_n287));
  INV_X1    g0087(.A(G77), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n286), .A2(new_n287), .B1(new_n288), .B2(new_n283), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n271), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n269), .A2(KEYINPUT68), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT68), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(G33), .A3(G41), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n291), .A2(new_n293), .A3(new_n268), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n294), .A2(G274), .ZN(new_n295));
  INV_X1    g0095(.A(G41), .ZN(new_n296));
  INV_X1    g0096(.A(G45), .ZN(new_n297));
  AOI21_X1  g0097(.A(G1), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n219), .B1(KEYINPUT68), .B2(new_n269), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n298), .B1(new_n299), .B2(new_n293), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n295), .A2(new_n298), .B1(G226), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n290), .A2(G190), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n290), .A2(new_n301), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G200), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n267), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT10), .ZN(new_n306));
  INV_X1    g0106(.A(new_n266), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n307), .B1(new_n303), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(G179), .B2(new_n303), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n243), .B1(new_n259), .B2(G20), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n263), .A2(new_n312), .B1(new_n261), .B2(new_n243), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT7), .B1(new_n276), .B2(new_n220), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n281), .A2(KEYINPUT7), .A3(new_n220), .A4(new_n282), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(G68), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G58), .ZN(new_n318));
  INV_X1    g0118(.A(G68), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(G20), .B1(new_n320), .B2(new_n249), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n246), .A2(G159), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(KEYINPUT16), .B1(new_n317), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n281), .A2(new_n220), .A3(new_n282), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT7), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n319), .B1(new_n328), .B2(new_n315), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n321), .A2(KEYINPUT16), .A3(new_n322), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n254), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT76), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n325), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n254), .ZN(new_n334));
  INV_X1    g0134(.A(new_n330), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n334), .B1(new_n317), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT16), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n329), .B2(new_n323), .ZN(new_n338));
  AOI21_X1  g0138(.A(KEYINPUT76), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n313), .B1(new_n333), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT18), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n272), .A2(new_n277), .ZN(new_n342));
  INV_X1    g0142(.A(G226), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G1698), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n342), .B(new_n344), .C1(new_n274), .C2(new_n275), .ZN(new_n345));
  AND3_X1   g0145(.A1(KEYINPUT77), .A2(G33), .A3(G87), .ZN(new_n346));
  AOI21_X1  g0146(.A(KEYINPUT77), .B1(G33), .B2(G87), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n271), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n294), .A2(G274), .A3(new_n298), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT78), .ZN(new_n353));
  INV_X1    g0153(.A(G179), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n300), .A2(G232), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n352), .A2(new_n353), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n350), .A2(new_n355), .A3(new_n351), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT78), .B1(new_n357), .B2(G179), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n308), .ZN(new_n359));
  AND3_X1   g0159(.A1(new_n356), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n340), .A2(new_n341), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G200), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(G190), .B2(new_n357), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n313), .B(new_n364), .C1(new_n333), .C2(new_n339), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT17), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n313), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n332), .B1(new_n325), .B2(new_n331), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n336), .A2(KEYINPUT76), .A3(new_n338), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n356), .A2(new_n358), .A3(new_n359), .ZN(new_n372));
  OAI21_X1  g0172(.A(KEYINPUT18), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(KEYINPUT17), .A3(new_n364), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n361), .A2(new_n367), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  XOR2_X1   g0175(.A(KEYINPUT15), .B(G87), .Z(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n377), .A2(new_n244), .ZN(new_n378));
  OAI22_X1  g0178(.A1(new_n243), .A2(new_n247), .B1(new_n220), .B2(new_n288), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n254), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n261), .A2(new_n254), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n264), .A2(G77), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n381), .A2(new_n383), .B1(new_n288), .B2(new_n261), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g0185(.A(new_n385), .B(KEYINPUT71), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n300), .A2(G244), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n351), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n276), .A2(G107), .ZN(new_n390));
  INV_X1    g0190(.A(G232), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n390), .B1(new_n286), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n278), .A2(new_n284), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n392), .B1(G238), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n389), .B1(new_n394), .B2(new_n270), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G200), .ZN(new_n396));
  INV_X1    g0196(.A(G190), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n386), .B(new_n396), .C1(new_n397), .C2(new_n395), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n395), .A2(new_n308), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n354), .B(new_n389), .C1(new_n394), .C2(new_n270), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(new_n400), .A3(new_n385), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n311), .A2(new_n375), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n259), .A2(G13), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n319), .A2(G20), .ZN(new_n405));
  AOI211_X1 g0205(.A(new_n404), .B(new_n405), .C1(KEYINPUT74), .C2(KEYINPUT12), .ZN(new_n406));
  NOR2_X1   g0206(.A1(KEYINPUT74), .A2(KEYINPUT12), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n406), .B(new_n407), .ZN(new_n408));
  OAI221_X1 g0208(.A(new_n405), .B1(new_n244), .B2(new_n288), .C1(new_n247), .C2(new_n250), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n409), .A2(new_n258), .A3(KEYINPUT11), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n381), .A2(G68), .A3(new_n264), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n408), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT11), .B1(new_n409), .B2(new_n258), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT75), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT72), .ZN(new_n416));
  INV_X1    g0216(.A(new_n298), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n294), .A2(G238), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(G97), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n280), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(G226), .A2(G1698), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n421), .B1(new_n391), .B2(G1698), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n420), .B1(new_n422), .B2(new_n283), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n351), .B(new_n418), .C1(new_n423), .C2(new_n270), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n416), .B1(new_n424), .B2(KEYINPUT13), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n391), .A2(G1698), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(G226), .B2(G1698), .ZN(new_n427));
  OAI22_X1  g0227(.A1(new_n427), .A2(new_n276), .B1(new_n280), .B2(new_n419), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n428), .A2(new_n271), .B1(new_n300), .B2(G238), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT13), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n429), .A2(KEYINPUT72), .A3(new_n430), .A4(new_n351), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n424), .A2(KEYINPUT13), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n425), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT14), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(new_n434), .A3(G169), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT73), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n424), .B2(KEYINPUT13), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n429), .A2(KEYINPUT73), .A3(new_n430), .A4(new_n351), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n437), .A2(new_n438), .A3(G179), .A4(new_n432), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n434), .B1(new_n433), .B2(G169), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n415), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n441), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n443), .A2(KEYINPUT75), .A3(new_n439), .A4(new_n435), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n414), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n433), .A2(G200), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n437), .A2(new_n438), .A3(G190), .A4(new_n432), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n446), .A2(new_n414), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n403), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(G107), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n261), .A2(new_n452), .B1(KEYINPUT89), .B2(KEYINPUT25), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT89), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT25), .ZN(new_n455));
  NOR4_X1   g0255(.A1(new_n260), .A2(new_n454), .A3(new_n455), .A4(G107), .ZN(new_n456));
  NOR2_X1   g0256(.A1(KEYINPUT89), .A2(KEYINPUT25), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n453), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(G87), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(KEYINPUT88), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n460), .B(new_n220), .C1(new_n275), .C2(new_n274), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT22), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n283), .A2(KEYINPUT22), .A3(new_n220), .A4(new_n460), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G116), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(G20), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT23), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n220), .B2(G107), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n452), .A2(KEYINPUT23), .A3(G20), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n463), .A2(new_n464), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT24), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n334), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT24), .A4(new_n470), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n458), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n259), .A2(G33), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n263), .A2(KEYINPUT80), .A3(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n255), .A2(new_n260), .A3(new_n476), .A4(new_n257), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT80), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G107), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n475), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n259), .B(G45), .C1(new_n296), .C2(KEYINPUT5), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  OR2_X1    g0285(.A1(KEYINPUT81), .A2(KEYINPUT5), .ZN(new_n486));
  NAND2_X1  g0286(.A1(KEYINPUT81), .A2(KEYINPUT5), .ZN(new_n487));
  AOI21_X1  g0287(.A(G41), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT82), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AND2_X1   g0290(.A1(KEYINPUT81), .A2(KEYINPUT5), .ZN(new_n491));
  NOR2_X1   g0291(.A1(KEYINPUT81), .A2(KEYINPUT5), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n489), .B(new_n296), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(G264), .B(new_n294), .C1(new_n490), .C2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n283), .A2(G257), .A3(G1698), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n283), .A2(G250), .A3(new_n277), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G294), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n271), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n296), .B1(new_n491), .B2(new_n492), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n484), .B1(new_n501), .B2(KEYINPUT82), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n295), .A2(new_n493), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n495), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n308), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n502), .A2(new_n493), .B1(new_n293), .B2(new_n299), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n506), .A2(G264), .B1(new_n271), .B2(new_n499), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n507), .A2(new_n354), .A3(new_n503), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n483), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(G190), .A3(new_n503), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n504), .A2(G200), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n510), .A2(new_n511), .A3(new_n475), .A4(new_n482), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n478), .A2(new_n479), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n478), .A2(new_n479), .ZN(new_n514));
  OAI21_X1  g0314(.A(G97), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n246), .A2(G77), .ZN(new_n516));
  XNOR2_X1  g0316(.A(new_n516), .B(KEYINPUT79), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT6), .ZN(new_n518));
  NOR3_X1   g0318(.A1(new_n518), .A2(new_n419), .A3(G107), .ZN(new_n519));
  XNOR2_X1  g0319(.A(G97), .B(G107), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n519), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n517), .B1(new_n220), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n452), .B1(new_n328), .B2(new_n315), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n254), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n261), .A2(new_n419), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n515), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(G257), .B(new_n294), .C1(new_n490), .C2(new_n494), .ZN(new_n527));
  OAI211_X1 g0327(.A(G244), .B(new_n277), .C1(new_n274), .C2(new_n275), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT4), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G283), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G250), .A2(G1698), .ZN(new_n533));
  NAND2_X1  g0333(.A1(KEYINPUT4), .A2(G244), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(G1698), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n532), .B1(new_n283), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n530), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n271), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n527), .A2(new_n538), .A3(new_n503), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n308), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n490), .A2(new_n494), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n541), .A2(new_n295), .B1(new_n271), .B2(new_n537), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n542), .A2(new_n354), .A3(new_n527), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n526), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(G107), .B1(new_n314), .B2(new_n316), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n545), .B(new_n517), .C1(new_n220), .C2(new_n521), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n546), .A2(new_n254), .B1(new_n419), .B2(new_n261), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n539), .A2(G200), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n527), .A2(new_n538), .A3(G190), .A4(new_n503), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n515), .A4(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n509), .A2(new_n512), .A3(new_n544), .A4(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(G244), .B(G1698), .C1(new_n274), .C2(new_n275), .ZN(new_n552));
  OAI211_X1 g0352(.A(G238), .B(new_n277), .C1(new_n274), .C2(new_n275), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(new_n553), .A3(new_n465), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n297), .A2(G1), .A3(G274), .ZN(new_n555));
  AOI21_X1  g0355(.A(G250), .B1(new_n259), .B2(G45), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n554), .A2(new_n271), .B1(new_n294), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(new_n362), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(G190), .B2(new_n558), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n283), .A2(new_n220), .A3(G68), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n244), .A2(new_n419), .ZN(new_n562));
  NOR3_X1   g0362(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n563));
  XNOR2_X1  g0363(.A(new_n563), .B(KEYINPUT83), .ZN(new_n564));
  AOI21_X1  g0364(.A(G20), .B1(new_n420), .B2(KEYINPUT19), .ZN(new_n565));
  OAI221_X1 g0365(.A(new_n561), .B1(KEYINPUT19), .B2(new_n562), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n566), .A2(new_n254), .B1(new_n261), .B2(new_n377), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n481), .A2(KEYINPUT84), .A3(G87), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT84), .B1(new_n481), .B2(G87), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n560), .B(new_n567), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n481), .A2(new_n376), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n558), .A2(new_n308), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n558), .A2(G179), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n572), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n551), .A2(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n531), .B(new_n220), .C1(G33), .C2(new_n419), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n220), .A2(G116), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n581), .A3(new_n254), .ZN(new_n582));
  XNOR2_X1  g0382(.A(new_n582), .B(KEYINPUT20), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n381), .A2(G116), .A3(new_n476), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n581), .B2(new_n404), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(G270), .B(new_n294), .C1(new_n490), .C2(new_n494), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n588), .A2(new_n503), .ZN(new_n589));
  OAI211_X1 g0389(.A(G264), .B(G1698), .C1(new_n274), .C2(new_n275), .ZN(new_n590));
  OAI211_X1 g0390(.A(G257), .B(new_n277), .C1(new_n274), .C2(new_n275), .ZN(new_n591));
  XNOR2_X1  g0391(.A(KEYINPUT85), .B(G303), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n590), .B(new_n591), .C1(new_n283), .C2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n354), .B1(new_n593), .B2(new_n271), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n587), .A2(new_n589), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(G169), .B1(new_n583), .B2(new_n585), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n593), .A2(new_n271), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n588), .A2(new_n503), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT86), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n588), .A2(KEYINPUT86), .A3(new_n503), .A4(new_n597), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n596), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n595), .B1(new_n602), .B2(KEYINPUT21), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n600), .A2(new_n601), .ZN(new_n604));
  INV_X1    g0404(.A(new_n596), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(KEYINPUT21), .A3(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT87), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n602), .A2(KEYINPUT87), .A3(KEYINPUT21), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n603), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n587), .B1(new_n604), .B2(G200), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n397), .B2(new_n604), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n578), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n451), .A2(new_n613), .ZN(G372));
  AND2_X1   g0414(.A1(new_n367), .A2(new_n374), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT91), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n401), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n399), .A2(KEYINPUT91), .A3(new_n400), .A4(new_n385), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n617), .A2(new_n448), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n615), .B1(new_n445), .B2(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n361), .A2(new_n373), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n306), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n623), .A2(new_n310), .ZN(new_n624));
  INV_X1    g0424(.A(new_n595), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n604), .A2(new_n605), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT21), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n609), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT87), .B1(new_n602), .B2(KEYINPUT21), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n628), .B(new_n509), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n550), .A2(new_n544), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n632), .A2(new_n570), .A3(new_n512), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT90), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n575), .B2(new_n573), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n574), .B(KEYINPUT90), .C1(new_n308), .C2(new_n558), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n572), .ZN(new_n639));
  INV_X1    g0439(.A(new_n544), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(new_n570), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n640), .A2(new_n570), .A3(new_n576), .A4(KEYINPUT26), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n634), .A2(new_n639), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n624), .B1(new_n451), .B2(new_n647), .ZN(G369));
  XNOR2_X1  g0448(.A(KEYINPUT92), .B(G330), .ZN(new_n649));
  INV_X1    g0449(.A(new_n610), .ZN(new_n650));
  OR3_X1    g0450(.A1(new_n404), .A2(KEYINPUT27), .A3(G20), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT27), .B1(new_n404), .B2(G20), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(G213), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(G343), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n650), .A2(new_n587), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n655), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n610), .B(new_n612), .C1(new_n586), .C2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n649), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n509), .A2(new_n655), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n483), .A2(new_n655), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n512), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n660), .B1(new_n509), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n660), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n610), .A2(new_n655), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n663), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n664), .A2(new_n665), .A3(new_n667), .ZN(G399));
  INV_X1    g0468(.A(G116), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n564), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n216), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G41), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n670), .A2(new_n672), .A3(new_n259), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n673), .B1(new_n223), .B2(new_n672), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT28), .Z(new_n675));
  INV_X1    g0475(.A(KEYINPUT96), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n507), .A2(new_n542), .A3(new_n527), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n588), .A2(new_n594), .A3(new_n558), .A4(new_n503), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT93), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT30), .ZN(new_n680));
  AND4_X1   g0480(.A1(new_n588), .A2(new_n594), .A3(new_n558), .A4(new_n503), .ZN(new_n681));
  INV_X1    g0481(.A(new_n539), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT93), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n681), .A2(new_n682), .A3(new_n683), .A4(new_n507), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n679), .A2(new_n680), .A3(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n558), .A2(G179), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n504), .A2(new_n539), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n604), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n495), .A2(new_n500), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n678), .A2(new_n539), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(KEYINPUT95), .B1(new_n691), .B2(KEYINPUT30), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT95), .ZN(new_n693));
  NOR4_X1   g0493(.A1(new_n677), .A2(new_n693), .A3(new_n678), .A4(new_n680), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n676), .B1(new_n689), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT31), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n681), .A2(new_n682), .A3(new_n507), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n693), .B1(new_n698), .B2(new_n680), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n691), .A2(KEYINPUT95), .A3(KEYINPUT30), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n701), .A2(KEYINPUT96), .A3(new_n685), .A4(new_n688), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n696), .A2(new_n697), .A3(new_n702), .ZN(new_n703));
  AOI22_X1  g0503(.A1(new_n703), .A2(new_n655), .B1(KEYINPUT31), .B2(new_n613), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n657), .A2(new_n697), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT94), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n695), .B1(new_n689), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n685), .A2(KEYINPUT94), .A3(new_n688), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n706), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n704), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n649), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n639), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n631), .B2(new_n633), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n642), .B1(new_n577), .B2(new_n544), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(new_n642), .B2(new_n641), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(KEYINPUT29), .A3(new_n657), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n647), .A2(new_n655), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n719), .B1(new_n720), .B2(KEYINPUT29), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n713), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n675), .B1(new_n722), .B2(G1), .ZN(G364));
  NAND2_X1  g0523(.A1(new_n656), .A2(new_n658), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n712), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT97), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n214), .A2(G20), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n259), .B1(new_n727), .B2(G45), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n672), .A2(new_n729), .ZN(new_n730));
  OR3_X1    g0530(.A1(new_n726), .A2(new_n659), .A3(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n730), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n219), .B1(G20), .B2(new_n308), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n220), .A2(G179), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G190), .A2(G200), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G159), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n736), .A2(KEYINPUT32), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n734), .A2(G190), .A3(G200), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n734), .A2(new_n397), .A3(G200), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI22_X1  g0542(.A1(new_n740), .A2(G87), .B1(new_n742), .B2(G107), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n220), .A2(new_n354), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G200), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G190), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n397), .A2(G179), .A3(G200), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n220), .ZN(new_n749));
  OAI221_X1 g0549(.A(new_n743), .B1(new_n319), .B2(new_n747), .C1(new_n419), .C2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(KEYINPUT32), .B1(new_n736), .B2(new_n737), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n745), .A2(new_n397), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n751), .B1(new_n753), .B2(new_n250), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n744), .A2(new_n735), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n744), .A2(G190), .A3(new_n362), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n283), .B1(new_n755), .B2(new_n288), .C1(new_n318), .C2(new_n756), .ZN(new_n757));
  OR4_X1    g0557(.A1(new_n738), .A2(new_n750), .A3(new_n754), .A4(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G322), .ZN(new_n759));
  INV_X1    g0559(.A(G311), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n756), .A2(new_n759), .B1(new_n755), .B2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n736), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n283), .B(new_n761), .C1(G329), .C2(new_n762), .ZN(new_n763));
  XOR2_X1   g0563(.A(new_n739), .B(KEYINPUT98), .Z(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G303), .ZN(new_n765));
  INV_X1    g0565(.A(new_n749), .ZN(new_n766));
  AOI22_X1  g0566(.A1(G294), .A2(new_n766), .B1(new_n752), .B2(G326), .ZN(new_n767));
  XNOR2_X1  g0567(.A(KEYINPUT33), .B(G317), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n746), .A2(new_n768), .B1(new_n742), .B2(G283), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n763), .A2(new_n765), .A3(new_n767), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n758), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n733), .B1(new_n772), .B2(KEYINPUT99), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(KEYINPUT99), .B2(new_n772), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n733), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n216), .A2(G355), .A3(new_n283), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n238), .A2(new_n297), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n216), .B(new_n276), .C1(G45), .C2(new_n222), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n779), .B1(G116), .B2(new_n216), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n732), .B(new_n774), .C1(new_n778), .C2(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(KEYINPUT100), .Z(new_n784));
  INV_X1    g0584(.A(new_n777), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n724), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n731), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT101), .ZN(G396));
  NAND4_X1  g0588(.A1(new_n617), .A2(new_n385), .A3(new_n618), .A4(new_n655), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n385), .A2(new_n655), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n398), .A2(new_n401), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(new_n647), .B2(new_n655), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n402), .A2(new_n655), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n796), .B1(new_n715), .B2(new_n645), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n730), .B1(new_n713), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n713), .B2(new_n799), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n733), .A2(new_n775), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n730), .B1(G77), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n756), .ZN(new_n804));
  INV_X1    g0604(.A(new_n755), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n804), .A2(G143), .B1(new_n805), .B2(G159), .ZN(new_n806));
  INV_X1    g0606(.A(G137), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n806), .B1(new_n753), .B2(new_n807), .C1(new_n245), .C2(new_n747), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT102), .Z(new_n809));
  OR2_X1    g0609(.A1(new_n809), .A2(KEYINPUT34), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(KEYINPUT34), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n276), .B1(new_n762), .B2(G132), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n812), .B1(new_n318), .B2(new_n749), .C1(new_n319), .C2(new_n741), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(G50), .B2(new_n764), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n810), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G294), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n756), .A2(new_n816), .B1(new_n736), .B2(new_n760), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n283), .B(new_n817), .C1(G116), .C2(new_n805), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n764), .A2(G107), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G97), .A2(new_n766), .B1(new_n752), .B2(G303), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n741), .A2(new_n459), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(G283), .B2(new_n746), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n818), .A2(new_n819), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n815), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n803), .B1(new_n824), .B2(new_n733), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n792), .B2(new_n776), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n801), .A2(new_n826), .ZN(G384));
  INV_X1    g0627(.A(new_n521), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n828), .A2(KEYINPUT35), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(KEYINPUT35), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n829), .A2(G116), .A3(new_n221), .A4(new_n830), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(KEYINPUT36), .Z(new_n832));
  OAI211_X1 g0632(.A(new_n223), .B(G77), .C1(new_n318), .C2(new_n319), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n250), .A2(G68), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n259), .B(G13), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n401), .A2(new_n655), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT103), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(new_n646), .B2(new_n795), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n414), .A2(new_n657), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n442), .A2(new_n444), .ZN(new_n843));
  INV_X1    g0643(.A(new_n414), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n842), .B1(new_n845), .B2(new_n448), .ZN(new_n846));
  NOR3_X1   g0646(.A1(new_n445), .A2(new_n449), .A3(new_n841), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n840), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT38), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n365), .B1(new_n371), .B2(new_n372), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n371), .A2(new_n653), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n851), .A2(KEYINPUT37), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n337), .A2(KEYINPUT104), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n329), .B2(new_n323), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n317), .A2(new_n324), .A3(new_n854), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n856), .A2(new_n857), .A3(new_n258), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n313), .ZN(new_n859));
  AND4_X1   g0659(.A1(new_n354), .A2(new_n350), .A3(new_n351), .A4(new_n355), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n860), .A2(new_n353), .B1(new_n308), .B2(new_n357), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n859), .A2(new_n861), .A3(new_n358), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n365), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT106), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n365), .A2(new_n862), .A3(KEYINPUT106), .ZN(new_n866));
  INV_X1    g0666(.A(new_n653), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT105), .B1(new_n859), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT105), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n869), .B(new_n653), .C1(new_n858), .C2(new_n313), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n865), .A2(new_n866), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n853), .B1(new_n872), .B2(KEYINPUT37), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n871), .B1(new_n621), .B2(new_n615), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n850), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n258), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n317), .A2(new_n324), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n876), .B1(new_n877), .B2(new_n855), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n368), .B1(new_n878), .B2(new_n857), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n869), .B1(new_n879), .B2(new_n653), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n859), .A2(KEYINPUT105), .A3(new_n867), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n375), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT37), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT106), .B1(new_n365), .B2(new_n862), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n885), .A2(new_n882), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n884), .B1(new_n886), .B2(new_n866), .ZN(new_n887));
  OAI211_X1 g0687(.A(KEYINPUT38), .B(new_n883), .C1(new_n887), .C2(new_n853), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n875), .A2(KEYINPUT107), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT107), .B1(new_n875), .B2(new_n888), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n849), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT37), .B1(new_n851), .B2(new_n852), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n340), .A2(new_n360), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n340), .A2(new_n867), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n893), .A2(new_n894), .A3(new_n884), .A4(new_n365), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n375), .A2(new_n852), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n850), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n888), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT39), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n875), .A2(new_n888), .A3(KEYINPUT39), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n902), .A2(new_n445), .A3(new_n657), .A4(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n621), .A2(new_n867), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n891), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT108), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT107), .ZN(new_n910));
  INV_X1    g0710(.A(new_n866), .ZN(new_n911));
  NOR3_X1   g0711(.A1(new_n911), .A2(new_n885), .A3(new_n882), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n895), .B1(new_n912), .B2(new_n884), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT38), .B1(new_n913), .B2(new_n883), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n873), .A2(new_n850), .A3(new_n874), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n910), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n875), .A2(new_n888), .A3(KEYINPUT107), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n905), .B1(new_n918), .B2(new_n849), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(KEYINPUT108), .A3(new_n904), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n909), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n624), .B1(new_n721), .B2(new_n451), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n921), .B(new_n922), .Z(new_n923));
  OAI21_X1  g0723(.A(new_n792), .B1(new_n846), .B2(new_n847), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n696), .A2(new_n702), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n705), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT109), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n925), .A2(KEYINPUT109), .A3(new_n705), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n704), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n924), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT40), .B1(new_n918), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n900), .A2(KEYINPUT40), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n933), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n704), .B1(new_n928), .B2(new_n929), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n937), .A2(new_n451), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n936), .A2(new_n938), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n939), .A2(new_n712), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n923), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n259), .B2(new_n727), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n923), .A2(new_n941), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n836), .B1(new_n943), .B2(new_n944), .ZN(G367));
  AND3_X1   g0745(.A1(new_n233), .A2(new_n216), .A3(new_n276), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n778), .B1(new_n216), .B2(new_n377), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n730), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NOR3_X1   g0748(.A1(new_n739), .A2(KEYINPUT46), .A3(new_n669), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n764), .A2(G116), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n949), .B1(new_n950), .B2(KEYINPUT46), .ZN(new_n951));
  AOI22_X1  g0751(.A1(G107), .A2(new_n766), .B1(new_n752), .B2(G311), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n283), .B1(new_n762), .B2(G317), .ZN(new_n953));
  INV_X1    g0753(.A(new_n592), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n804), .A2(new_n954), .B1(new_n805), .B2(G283), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n746), .A2(G294), .B1(new_n742), .B2(G97), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n952), .A2(new_n953), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n755), .A2(new_n250), .B1(new_n736), .B2(new_n807), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(G150), .B2(new_n804), .ZN(new_n959));
  AOI22_X1  g0759(.A1(G143), .A2(new_n752), .B1(new_n746), .B2(G159), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n766), .A2(G68), .B1(new_n740), .B2(G58), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n283), .B1(new_n741), .B2(new_n288), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT114), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n951), .A2(new_n957), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT47), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n948), .B1(new_n966), .B2(new_n733), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n655), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n969), .A2(new_n639), .A3(new_n570), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n639), .B2(new_n969), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n967), .B1(new_n971), .B2(new_n785), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT115), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n666), .B(new_n663), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(new_n659), .ZN(new_n976));
  AND3_X1   g0776(.A1(new_n713), .A2(new_n976), .A3(new_n721), .ZN(new_n977));
  INV_X1    g0777(.A(new_n526), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n632), .B1(new_n978), .B2(new_n657), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n640), .A2(new_n655), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n667), .A2(new_n665), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(KEYINPUT110), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT110), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n667), .A2(new_n984), .A3(new_n665), .A4(new_n981), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT45), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n981), .B1(new_n667), .B2(new_n665), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n989), .A2(KEYINPUT44), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(KEYINPUT44), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n664), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(KEYINPUT111), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n983), .A2(KEYINPUT45), .A3(new_n985), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n988), .A2(new_n992), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n977), .A2(new_n996), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n986), .A2(new_n987), .B1(new_n990), .B2(new_n991), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n994), .B1(new_n998), .B2(new_n995), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n722), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n672), .B(KEYINPUT41), .Z(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  AND3_X1   g0802(.A1(new_n1000), .A2(KEYINPUT112), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(KEYINPUT112), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n728), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n666), .A2(new_n663), .A3(new_n981), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1006), .A2(KEYINPUT42), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n544), .B1(new_n979), .B2(new_n509), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n1006), .A2(KEYINPUT42), .B1(new_n657), .B2(new_n1008), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n1007), .A2(new_n1009), .B1(KEYINPUT43), .B2(new_n971), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n993), .A2(new_n981), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  AND3_X1   g0814(.A1(new_n1005), .A2(KEYINPUT113), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(KEYINPUT113), .B1(new_n1005), .B2(new_n1014), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n974), .B1(new_n1015), .B2(new_n1016), .ZN(G387));
  NAND2_X1  g0817(.A1(new_n976), .A2(new_n729), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n663), .A2(new_n785), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n755), .A2(new_n319), .B1(new_n736), .B2(new_n245), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n276), .B(new_n1020), .C1(G50), .C2(new_n804), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n740), .A2(G77), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n243), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n376), .A2(new_n766), .B1(new_n746), .B2(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n752), .A2(G159), .B1(new_n742), .B2(G97), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n283), .B1(new_n762), .B2(G326), .ZN(new_n1027));
  INV_X1    g0827(.A(G283), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n749), .A2(new_n1028), .B1(new_n739), .B2(new_n816), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n804), .A2(G317), .B1(new_n805), .B2(new_n954), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n753), .B2(new_n759), .C1(new_n760), .C2(new_n747), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT48), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1029), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n1032), .B2(new_n1031), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT49), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1027), .B1(new_n669), .B2(new_n741), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1026), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1038), .A2(KEYINPUT116), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(KEYINPUT116), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1039), .A2(new_n733), .A3(new_n1040), .ZN(new_n1041));
  OR3_X1    g0841(.A1(new_n243), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1042));
  OAI21_X1  g0842(.A(KEYINPUT50), .B1(new_n243), .B2(G50), .ZN(new_n1043));
  AOI21_X1  g0843(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n670), .B1(new_n1045), .B2(new_n276), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n283), .A2(new_n297), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1046), .B1(new_n229), .B2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1048), .A2(new_n671), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n778), .B1(new_n452), .B2(new_n216), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1041), .B(new_n730), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n977), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n672), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n722), .A2(new_n976), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1018), .B1(new_n1019), .B2(new_n1051), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT117), .ZN(G393));
  INV_X1    g0856(.A(new_n672), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n997), .A2(new_n999), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n998), .A2(new_n664), .A3(new_n995), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT118), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n988), .A2(new_n992), .A3(new_n995), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n993), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1061), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1057), .B(new_n1058), .C1(new_n1065), .C2(new_n1052), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n241), .A2(new_n216), .A3(new_n276), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1067), .B(new_n778), .C1(new_n419), .C2(new_n216), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n730), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n766), .A2(G77), .B1(new_n805), .B2(new_n1023), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n250), .B2(new_n747), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT119), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n753), .A2(new_n245), .B1(new_n737), .B2(new_n756), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT51), .ZN(new_n1074));
  INV_X1    g0874(.A(G143), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n283), .B1(new_n736), .B2(new_n1075), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n821), .B(new_n1076), .C1(G68), .C2(new_n740), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1072), .A2(new_n1074), .A3(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G317), .A2(new_n752), .B1(new_n804), .B2(G311), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT52), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n747), .A2(new_n592), .B1(new_n452), .B2(new_n741), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n276), .B1(new_n736), .B2(new_n759), .C1(new_n816), .C2(new_n755), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n749), .A2(new_n669), .B1(new_n739), .B2(new_n1028), .ZN(new_n1083));
  OR3_X1    g0883(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1078), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1069), .B1(new_n1085), .B2(new_n733), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n981), .B2(new_n785), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n1065), .B2(new_n728), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1066), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(G390));
  NAND3_X1  g0890(.A1(new_n718), .A2(new_n657), .A3(new_n792), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n838), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n712), .B(new_n792), .C1(new_n704), .C2(new_n710), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n845), .A2(new_n448), .A3(new_n842), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n841), .B1(new_n445), .B2(new_n449), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1092), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(KEYINPUT109), .B1(new_n925), .B2(new_n705), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n927), .B(new_n706), .C1(new_n696), .C2(new_n702), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g0901(.A(G330), .B(new_n792), .C1(new_n1101), .C2(new_n704), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1095), .A2(KEYINPUT120), .A3(new_n1096), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT120), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n846), .B2(new_n847), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1102), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1098), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1093), .A2(new_n848), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n793), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1109));
  OAI211_X1 g0909(.A(G330), .B(new_n1109), .C1(new_n1101), .C2(new_n704), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n840), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1107), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n451), .ZN(new_n1115));
  INV_X1    g0915(.A(G330), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n937), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n922), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1110), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1097), .B1(new_n797), .B2(new_n839), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n445), .A2(new_n657), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n902), .A2(new_n903), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT38), .B1(new_n896), .B2(new_n897), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1122), .B1(new_n915), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1105), .A2(new_n1103), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1125), .B1(new_n1126), .B2(new_n1092), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1120), .B1(new_n1123), .B2(new_n1127), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n846), .A2(new_n847), .A3(new_n1104), .ZN(new_n1129));
  AOI21_X1  g0929(.A(KEYINPUT120), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n655), .B(new_n793), .C1(new_n715), .C2(new_n717), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n1129), .A2(new_n1130), .B1(new_n1131), .B2(new_n839), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1125), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n872), .A2(KEYINPUT37), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n874), .B1(new_n1135), .B2(new_n895), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1124), .B1(new_n1136), .B2(KEYINPUT38), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n903), .B1(new_n1137), .B2(KEYINPUT39), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n711), .A2(new_n712), .A3(new_n792), .A4(new_n1097), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1134), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1128), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1057), .B1(new_n1119), .B2(new_n1143), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1106), .A2(new_n1098), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1117), .A2(new_n1115), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1146), .B(new_n624), .C1(new_n451), .C2(new_n721), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1148), .A2(new_n1142), .A3(new_n1128), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1144), .A2(new_n1149), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n756), .A2(new_n669), .B1(new_n755), .B2(new_n419), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n283), .B(new_n1151), .C1(G294), .C2(new_n762), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n764), .A2(G87), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n766), .A2(G77), .B1(new_n742), .B2(G68), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(G107), .A2(new_n746), .B1(new_n752), .B2(G283), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(G159), .A2(new_n766), .B1(new_n752), .B2(G128), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(new_n250), .B2(new_n741), .C1(new_n807), .C2(new_n747), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT54), .B(G143), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n804), .A2(G132), .B1(new_n805), .B2(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n740), .A2(new_n1162), .A3(G150), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1162), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n739), .B2(new_n245), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n276), .B1(new_n762), .B2(G125), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1161), .A2(new_n1163), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1156), .B1(new_n1158), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(KEYINPUT122), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n733), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1168), .A2(KEYINPUT122), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n730), .B1(new_n1023), .B2(new_n802), .C1(new_n1170), .C2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n1138), .B2(new_n775), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1173), .B(KEYINPUT123), .Z(new_n1174));
  NAND3_X1  g0974(.A1(new_n1128), .A2(new_n1142), .A3(new_n729), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1150), .A2(new_n1174), .A3(new_n1175), .ZN(G378));
  OAI21_X1  g0976(.A(new_n1109), .B1(new_n1101), .B2(new_n704), .ZN(new_n1177));
  OAI21_X1  g0977(.A(G330), .B1(new_n1177), .B2(new_n934), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n307), .A2(new_n653), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n311), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n311), .A2(new_n1181), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1180), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1184), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1186), .A2(new_n1182), .A3(new_n1179), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  NOR3_X1   g0988(.A1(new_n933), .A2(new_n1178), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT40), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n889), .A2(new_n890), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1191), .B1(new_n1192), .B2(new_n1177), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1116), .B1(new_n932), .B2(new_n935), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1190), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT108), .B1(new_n919), .B2(new_n904), .ZN(new_n1196));
  AND4_X1   g0996(.A1(KEYINPUT108), .A2(new_n891), .A3(new_n904), .A4(new_n906), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n1189), .A2(new_n1195), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1118), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1188), .B1(new_n933), .B2(new_n1178), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1193), .A2(new_n1194), .A3(new_n1190), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1200), .A2(new_n1201), .A3(new_n909), .A4(new_n920), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1198), .A2(new_n1199), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT57), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1198), .A2(new_n1199), .A3(KEYINPUT57), .A4(new_n1202), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(new_n672), .A3(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1198), .A2(new_n729), .A3(new_n1202), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1188), .A2(new_n775), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n730), .B1(G50), .B2(new_n802), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n753), .A2(new_n669), .B1(new_n741), .B2(new_n318), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G97), .B2(new_n746), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n276), .A2(new_n296), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G283), .B2(new_n762), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n804), .A2(G107), .B1(new_n805), .B2(new_n376), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n766), .A2(G68), .B1(new_n740), .B2(G77), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1212), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT58), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1213), .B(new_n250), .C1(G33), .C2(G41), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n746), .A2(G132), .ZN(new_n1222));
  INV_X1    g1022(.A(G125), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1222), .B1(new_n753), .B2(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n804), .A2(G128), .B1(new_n805), .B2(G137), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n739), .B2(new_n1159), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1224), .B(new_n1226), .C1(G150), .C2(new_n766), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n742), .A2(G159), .ZN(new_n1230));
  AOI211_X1 g1030(.A(G33), .B(G41), .C1(new_n762), .C2(G124), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1221), .B1(new_n1218), .B2(new_n1217), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1210), .B1(new_n1234), .B2(new_n733), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1209), .A2(new_n1235), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1208), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1207), .A2(new_n1237), .ZN(G375));
  NOR2_X1   g1038(.A1(new_n1126), .A2(new_n776), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(KEYINPUT124), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n730), .B1(G68), .B2(new_n802), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n756), .A2(new_n807), .B1(new_n755), .B2(new_n245), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n276), .B(new_n1242), .C1(G128), .C2(new_n762), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n764), .A2(G159), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n766), .A2(G50), .B1(new_n742), .B2(G58), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(G132), .A2(new_n752), .B1(new_n746), .B2(new_n1160), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .A4(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n756), .A2(new_n1028), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n276), .B1(new_n755), .B2(new_n452), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n1248), .B(new_n1249), .C1(G303), .C2(new_n762), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n764), .A2(G97), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n766), .A2(new_n376), .B1(new_n742), .B2(G77), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(G116), .A2(new_n746), .B1(new_n752), .B2(G294), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .A4(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1247), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1241), .B1(new_n1255), .B2(new_n733), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1240), .A2(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1257), .B1(new_n728), .B2(new_n1145), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1119), .A2(new_n1002), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1259), .A2(new_n1261), .ZN(G381));
  OR4_X1    g1062(.A1(G396), .A2(G393), .A3(G384), .A4(G381), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1150), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1089), .A2(new_n1264), .ZN(new_n1265));
  OR4_X1    g1065(.A1(G387), .A2(new_n1263), .A3(G375), .A4(new_n1265), .ZN(G407));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n654), .ZN(new_n1267));
  OAI211_X1 g1067(.A(G407), .B(G213), .C1(G375), .C2(new_n1267), .ZN(G409));
  XOR2_X1   g1068(.A(G393), .B(G396), .Z(new_n1269));
  NAND2_X1  g1069(.A1(G387), .A2(new_n1089), .ZN(new_n1270));
  OAI211_X1 g1070(.A(G390), .B(new_n974), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1269), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1270), .A2(new_n1269), .A3(new_n1271), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(G213), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1276), .A2(G343), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1198), .A2(KEYINPUT125), .A3(new_n1202), .ZN(new_n1278));
  AOI21_X1  g1078(.A(KEYINPUT125), .B1(new_n1198), .B2(new_n1202), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1278), .A2(new_n1279), .A3(new_n728), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1236), .B1(new_n1203), .B2(new_n1001), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1264), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1207), .A2(G378), .A3(new_n1237), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1277), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT126), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1145), .A2(new_n1147), .A3(KEYINPUT60), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n672), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT60), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1260), .B1(new_n1148), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(G384), .B1(new_n1291), .B2(new_n1259), .ZN(new_n1292));
  INV_X1    g1092(.A(G384), .ZN(new_n1293));
  AOI211_X1 g1093(.A(new_n1293), .B(new_n1258), .C1(new_n1288), .C2(new_n1290), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1285), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1119), .A2(KEYINPUT60), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1287), .B1(new_n1296), .B2(new_n1260), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1293), .B1(new_n1297), .B2(new_n1258), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1291), .A2(G384), .A3(new_n1259), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1298), .A2(KEYINPUT126), .A3(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1295), .A2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT62), .B1(new_n1284), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT127), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1277), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1303), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  AOI211_X1 g1106(.A(KEYINPUT127), .B(new_n1277), .C1(new_n1282), .C2(new_n1283), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  AND2_X1   g1108(.A1(new_n1301), .A2(KEYINPUT62), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1302), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1277), .A2(G2897), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1311), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1312), .B1(new_n1301), .B2(new_n1311), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1313), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT61), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1275), .B1(new_n1310), .B2(new_n1316), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1270), .A2(new_n1269), .A3(new_n1271), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1318), .A2(new_n1272), .ZN(new_n1319));
  AND2_X1   g1119(.A1(new_n1301), .A2(KEYINPUT63), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1308), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1284), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1313), .A2(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT63), .B1(new_n1284), .B2(new_n1301), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1324), .A2(KEYINPUT61), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1319), .A2(new_n1321), .A3(new_n1323), .A4(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1317), .A2(new_n1326), .ZN(G405));
  NAND2_X1  g1127(.A1(G375), .A2(new_n1264), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(new_n1283), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1329), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1330), .B1(new_n1301), .B2(new_n1329), .ZN(new_n1331));
  XNOR2_X1  g1131(.A(new_n1319), .B(new_n1331), .ZN(G402));
endmodule


