

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750;

  XNOR2_X1 U371 ( .A(n709), .B(n353), .ZN(n712) );
  XOR2_X1 U372 ( .A(KEYINPUT62), .B(n620), .Z(n621) );
  XOR2_X1 U373 ( .A(n703), .B(KEYINPUT59), .Z(n704) );
  XNOR2_X1 U374 ( .A(n370), .B(KEYINPUT32), .ZN(n368) );
  NOR2_X1 U375 ( .A1(n351), .A2(n572), .ZN(n514) );
  NOR2_X1 U376 ( .A1(n355), .A2(n645), .ZN(n678) );
  XNOR2_X1 U377 ( .A(n493), .B(KEYINPUT104), .ZN(n351) );
  OR2_X1 U378 ( .A1(n385), .A2(n532), .ZN(n413) );
  NOR2_X1 U379 ( .A1(n586), .A2(n530), .ZN(n522) );
  XNOR2_X1 U380 ( .A(n542), .B(KEYINPUT100), .ZN(n515) );
  OR2_X1 U381 ( .A1(n703), .A2(G902), .ZN(n381) );
  NAND2_X1 U382 ( .A1(n620), .A2(n473), .ZN(n471) );
  XNOR2_X1 U383 ( .A(n415), .B(n498), .ZN(n626) );
  XNOR2_X1 U384 ( .A(n448), .B(n469), .ZN(n699) );
  XNOR2_X1 U385 ( .A(n444), .B(n720), .ZN(n482) );
  XNOR2_X1 U386 ( .A(n728), .B(n350), .ZN(n445) );
  XNOR2_X1 U387 ( .A(n465), .B(KEYINPUT73), .ZN(n444) );
  XNOR2_X1 U388 ( .A(n439), .B(KEYINPUT89), .ZN(n728) );
  XNOR2_X1 U389 ( .A(n440), .B(n483), .ZN(n350) );
  BUF_X1 U390 ( .A(G140), .Z(n354) );
  BUF_X1 U391 ( .A(G143), .Z(n349) );
  INV_X1 U392 ( .A(KEYINPUT12), .ZN(n373) );
  XNOR2_X1 U393 ( .A(G137), .B(G140), .ZN(n439) );
  INV_X1 U394 ( .A(G143), .ZN(n446) );
  XNOR2_X1 U395 ( .A(n419), .B(G146), .ZN(n476) );
  XOR2_X2 U396 ( .A(KEYINPUT65), .B(n602), .Z(n603) );
  XNOR2_X2 U397 ( .A(n567), .B(n566), .ZN(n588) );
  XNOR2_X1 U398 ( .A(n372), .B(n507), .ZN(n509) );
  NAND2_X1 U399 ( .A1(n352), .A2(n603), .ZN(n390) );
  NAND2_X1 U400 ( .A1(n377), .A2(n379), .ZN(n352) );
  XNOR2_X1 U401 ( .A(n710), .B(KEYINPUT122), .ZN(n353) );
  NOR2_X2 U402 ( .A1(n587), .A2(n580), .ZN(n570) );
  XNOR2_X2 U403 ( .A(n410), .B(n409), .ZN(n748) );
  NOR2_X2 U404 ( .A1(n536), .A2(n535), .ZN(n538) );
  XNOR2_X2 U405 ( .A(n475), .B(n447), .ZN(n494) );
  XNOR2_X1 U406 ( .A(n476), .B(n397), .ZN(n727) );
  INV_X1 U407 ( .A(G953), .ZN(n738) );
  NOR2_X2 U408 ( .A1(n591), .A2(n402), .ZN(n547) );
  AND2_X2 U409 ( .A1(n608), .A2(n361), .ZN(n377) );
  NOR2_X2 U410 ( .A1(n745), .A2(n575), .ZN(n369) );
  NOR2_X1 U411 ( .A1(n744), .A2(n518), .ZN(n519) );
  XNOR2_X1 U412 ( .A(n519), .B(KEYINPUT79), .ZN(n536) );
  XNOR2_X1 U413 ( .A(n401), .B(n400), .ZN(n750) );
  OR2_X1 U414 ( .A1(n654), .A2(n546), .ZN(n401) );
  NOR2_X1 U415 ( .A1(n532), .A2(n387), .ZN(n384) );
  XNOR2_X1 U416 ( .A(n540), .B(KEYINPUT106), .ZN(n398) );
  XNOR2_X1 U417 ( .A(n434), .B(n433), .ZN(n568) );
  XNOR2_X1 U418 ( .A(n373), .B(KEYINPUT11), .ZN(n372) );
  INV_X1 U419 ( .A(G125), .ZN(n419) );
  XNOR2_X2 U420 ( .A(n469), .B(n468), .ZN(n620) );
  XOR2_X1 U421 ( .A(KEYINPUT69), .B(G131), .Z(n501) );
  INV_X1 U422 ( .A(n727), .ZN(n396) );
  INV_X1 U423 ( .A(KEYINPUT86), .ZN(n389) );
  XNOR2_X1 U424 ( .A(n371), .B(KEYINPUT22), .ZN(n578) );
  NOR2_X1 U425 ( .A1(n588), .A2(n356), .ZN(n371) );
  BUF_X1 U426 ( .A(n568), .Z(n660) );
  INV_X1 U427 ( .A(n750), .ZN(n551) );
  INV_X1 U428 ( .A(G237), .ZN(n472) );
  INV_X1 U429 ( .A(G134), .ZN(n447) );
  INV_X1 U430 ( .A(n520), .ZN(n403) );
  XNOR2_X1 U431 ( .A(n474), .B(n405), .ZN(n404) );
  OR2_X1 U432 ( .A1(n626), .A2(G902), .ZN(n414) );
  NOR2_X1 U433 ( .A1(n710), .A2(G902), .ZN(n434) );
  XNOR2_X1 U434 ( .A(n423), .B(n416), .ZN(n424) );
  XOR2_X1 U435 ( .A(G128), .B(G110), .Z(n416) );
  XNOR2_X1 U436 ( .A(n484), .B(n483), .ZN(n497) );
  XNOR2_X1 U437 ( .A(G122), .B(G116), .ZN(n484) );
  XOR2_X1 U438 ( .A(KEYINPUT98), .B(n354), .Z(n504) );
  XNOR2_X1 U439 ( .A(n349), .B(G122), .ZN(n503) );
  XNOR2_X1 U440 ( .A(n509), .B(n417), .ZN(n510) );
  XNOR2_X1 U441 ( .A(KEYINPUT97), .B(KEYINPUT99), .ZN(n507) );
  INV_X1 U442 ( .A(KEYINPUT10), .ZN(n397) );
  XNOR2_X1 U443 ( .A(G104), .B(G113), .ZN(n502) );
  INV_X1 U444 ( .A(KEYINPUT36), .ZN(n412) );
  OR2_X1 U445 ( .A1(n689), .A2(n693), .ZN(n408) );
  NAND2_X1 U446 ( .A1(n578), .A2(n579), .ZN(n370) );
  INV_X1 U447 ( .A(KEYINPUT44), .ZN(n392) );
  INV_X1 U448 ( .A(KEYINPUT70), .ZN(n537) );
  INV_X1 U449 ( .A(KEYINPUT30), .ZN(n405) );
  XOR2_X1 U450 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n457) );
  XNOR2_X1 U451 ( .A(G116), .B(G137), .ZN(n459) );
  NOR2_X1 U452 ( .A1(G953), .A2(G237), .ZN(n508) );
  NAND2_X1 U453 ( .A1(n673), .A2(n672), .ZN(n540) );
  NOR2_X1 U454 ( .A1(n541), .A2(n530), .ZN(n383) );
  XNOR2_X1 U455 ( .A(n438), .B(KEYINPUT68), .ZN(n656) );
  NOR2_X1 U456 ( .A1(n568), .A2(n661), .ZN(n438) );
  XNOR2_X1 U457 ( .A(G119), .B(G113), .ZN(n463) );
  INV_X1 U458 ( .A(KEYINPUT72), .ZN(n462) );
  XNOR2_X1 U459 ( .A(G104), .B(KEYINPUT75), .ZN(n443) );
  XNOR2_X1 U460 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n478) );
  XNOR2_X1 U461 ( .A(n395), .B(n394), .ZN(n710) );
  XNOR2_X1 U462 ( .A(n427), .B(n420), .ZN(n394) );
  XNOR2_X1 U463 ( .A(n424), .B(n396), .ZN(n395) );
  XNOR2_X1 U464 ( .A(n494), .B(n500), .ZN(n415) );
  XNOR2_X1 U465 ( .A(n382), .B(n511), .ZN(n703) );
  XNOR2_X1 U466 ( .A(n510), .B(n727), .ZN(n382) );
  INV_X1 U467 ( .A(n399), .ZN(n558) );
  XNOR2_X1 U468 ( .A(KEYINPUT42), .B(KEYINPUT107), .ZN(n400) );
  INV_X1 U469 ( .A(KEYINPUT108), .ZN(n409) );
  XNOR2_X1 U470 ( .A(n413), .B(n412), .ZN(n411) );
  XNOR2_X1 U471 ( .A(n367), .B(KEYINPUT35), .ZN(n745) );
  INV_X1 U472 ( .A(KEYINPUT77), .ZN(n366) );
  NOR2_X1 U473 ( .A1(n546), .A2(n561), .ZN(n525) );
  XNOR2_X1 U474 ( .A(n514), .B(n513), .ZN(n744) );
  NAND2_X1 U475 ( .A1(n578), .A2(n359), .ZN(n638) );
  NOR2_X1 U476 ( .A1(n406), .A2(G953), .ZN(n694) );
  XNOR2_X1 U477 ( .A(n407), .B(KEYINPUT118), .ZN(n406) );
  OR2_X1 U478 ( .A1(n690), .A2(n408), .ZN(n407) );
  XNOR2_X1 U479 ( .A(n368), .B(n363), .ZN(G21) );
  AND2_X1 U480 ( .A1(n515), .A2(n516), .ZN(n355) );
  OR2_X1 U481 ( .A1(n676), .A2(n661), .ZN(n356) );
  XNOR2_X1 U482 ( .A(n414), .B(G478), .ZN(n541) );
  XOR2_X1 U483 ( .A(KEYINPUT13), .B(G475), .Z(n357) );
  XOR2_X1 U484 ( .A(n655), .B(n389), .Z(n358) );
  AND2_X1 U485 ( .A1(n581), .A2(n569), .ZN(n359) );
  AND2_X1 U486 ( .A1(n581), .A2(n580), .ZN(n360) );
  AND2_X1 U487 ( .A1(n560), .A2(n378), .ZN(n361) );
  INV_X1 U488 ( .A(G107), .ZN(n483) );
  NAND2_X1 U489 ( .A1(n601), .A2(n600), .ZN(n362) );
  XOR2_X1 U490 ( .A(G119), .B(KEYINPUT125), .Z(n363) );
  NAND2_X1 U491 ( .A1(n411), .A2(n358), .ZN(n410) );
  BUF_X1 U492 ( .A(n604), .Z(n650) );
  INV_X1 U493 ( .A(n655), .ZN(n581) );
  XNOR2_X1 U494 ( .A(n524), .B(n539), .ZN(n673) );
  BUF_X1 U495 ( .A(n524), .Z(n399) );
  NAND2_X1 U496 ( .A1(n655), .A2(n656), .ZN(n364) );
  NAND2_X1 U497 ( .A1(n655), .A2(n656), .ZN(n587) );
  NAND2_X1 U498 ( .A1(n524), .A2(n672), .ZN(n388) );
  BUF_X1 U499 ( .A(n681), .Z(n691) );
  INV_X1 U500 ( .A(n586), .ZN(n365) );
  XNOR2_X1 U501 ( .A(n366), .B(n525), .ZN(n526) );
  NAND2_X1 U502 ( .A1(n574), .A2(n573), .ZN(n367) );
  NAND2_X1 U503 ( .A1(n578), .A2(n360), .ZN(n583) );
  NAND2_X1 U504 ( .A1(n369), .A2(n368), .ZN(n393) );
  NAND2_X1 U505 ( .A1(n391), .A2(n598), .ZN(n599) );
  NOR2_X2 U506 ( .A1(G902), .A2(n699), .ZN(n449) );
  NAND2_X1 U507 ( .A1(n404), .A2(n403), .ZN(n402) );
  NAND2_X1 U508 ( .A1(n376), .A2(n600), .ZN(n375) );
  NAND2_X1 U509 ( .A1(n375), .A2(n374), .ZN(n379) );
  NAND2_X1 U510 ( .A1(n604), .A2(n362), .ZN(n374) );
  INV_X1 U511 ( .A(n604), .ZN(n376) );
  NAND2_X1 U512 ( .A1(n608), .A2(n560), .ZN(n736) );
  NAND2_X1 U513 ( .A1(n489), .A2(KEYINPUT82), .ZN(n378) );
  XNOR2_X2 U514 ( .A(n381), .B(n357), .ZN(n542) );
  NAND2_X1 U515 ( .A1(n515), .A2(n383), .ZN(n387) );
  INV_X1 U516 ( .A(n387), .ZN(n386) );
  NAND2_X1 U517 ( .A1(n386), .A2(n399), .ZN(n385) );
  INV_X1 U518 ( .A(n565), .ZN(n561) );
  XNOR2_X2 U519 ( .A(n388), .B(KEYINPUT19), .ZN(n565) );
  XNOR2_X2 U520 ( .A(n492), .B(n491), .ZN(n524) );
  XNOR2_X2 U521 ( .A(n529), .B(KEYINPUT1), .ZN(n655) );
  XNOR2_X2 U522 ( .A(n449), .B(n450), .ZN(n529) );
  NAND2_X1 U523 ( .A1(n390), .A2(n609), .ZN(n611) );
  XNOR2_X1 U524 ( .A(n393), .B(n392), .ZN(n391) );
  NOR2_X1 U525 ( .A1(n398), .A2(n676), .ZN(n545) );
  NOR2_X1 U526 ( .A1(n398), .A2(n678), .ZN(n679) );
  NAND2_X1 U527 ( .A1(n547), .A2(n399), .ZN(n493) );
  XNOR2_X2 U528 ( .A(n729), .B(G146), .ZN(n469) );
  XNOR2_X2 U529 ( .A(n494), .B(n501), .ZN(n729) );
  XNOR2_X2 U530 ( .A(n442), .B(KEYINPUT4), .ZN(n465) );
  BUF_X1 U531 ( .A(n654), .Z(n692) );
  AND2_X1 U532 ( .A1(n508), .A2(G214), .ZN(n417) );
  OR2_X1 U533 ( .A1(n564), .A2(n563), .ZN(n418) );
  INV_X1 U534 ( .A(n743), .ZN(n550) );
  INV_X1 U535 ( .A(KEYINPUT82), .ZN(n600) );
  INV_X1 U536 ( .A(KEYINPUT5), .ZN(n458) );
  XNOR2_X1 U537 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U538 ( .A(n461), .B(n460), .ZN(n467) );
  XNOR2_X1 U539 ( .A(n487), .B(n486), .ZN(n722) );
  INV_X1 U540 ( .A(KEYINPUT105), .ZN(n513) );
  INV_X1 U541 ( .A(KEYINPUT63), .ZN(n624) );
  INV_X1 U542 ( .A(KEYINPUT121), .ZN(n629) );
  INV_X1 U543 ( .A(n439), .ZN(n420) );
  XOR2_X1 U544 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n422) );
  XNOR2_X1 U545 ( .A(G119), .B(KEYINPUT23), .ZN(n421) );
  XNOR2_X1 U546 ( .A(n422), .B(n421), .ZN(n423) );
  NAND2_X1 U547 ( .A1(n738), .A2(G234), .ZN(n426) );
  XNOR2_X1 U548 ( .A(KEYINPUT81), .B(KEYINPUT8), .ZN(n425) );
  XNOR2_X1 U549 ( .A(n426), .B(n425), .ZN(n499) );
  NAND2_X1 U550 ( .A1(G221), .A2(n499), .ZN(n427) );
  XOR2_X1 U551 ( .A(KEYINPUT25), .B(KEYINPUT76), .Z(n432) );
  XNOR2_X1 U552 ( .A(G902), .B(KEYINPUT87), .ZN(n429) );
  INV_X1 U553 ( .A(KEYINPUT15), .ZN(n428) );
  XNOR2_X1 U554 ( .A(n429), .B(n428), .ZN(n489) );
  NAND2_X1 U555 ( .A1(n489), .A2(G234), .ZN(n430) );
  XNOR2_X1 U556 ( .A(n430), .B(KEYINPUT20), .ZN(n435) );
  NAND2_X1 U557 ( .A1(n435), .A2(G217), .ZN(n431) );
  XNOR2_X1 U558 ( .A(n432), .B(n431), .ZN(n433) );
  AND2_X1 U559 ( .A1(n435), .A2(G221), .ZN(n437) );
  XNOR2_X1 U560 ( .A(KEYINPUT91), .B(KEYINPUT21), .ZN(n436) );
  XNOR2_X1 U561 ( .A(n437), .B(n436), .ZN(n661) );
  XNOR2_X1 U562 ( .A(KEYINPUT71), .B(G469), .ZN(n450) );
  NAND2_X1 U563 ( .A1(G227), .A2(n738), .ZN(n440) );
  XNOR2_X2 U564 ( .A(G101), .B(KEYINPUT67), .ZN(n442) );
  XNOR2_X1 U565 ( .A(n443), .B(G110), .ZN(n720) );
  XNOR2_X1 U566 ( .A(n482), .B(n445), .ZN(n448) );
  XNOR2_X2 U567 ( .A(n446), .B(G128), .ZN(n475) );
  NAND2_X1 U568 ( .A1(n656), .A2(n529), .ZN(n591) );
  NAND2_X1 U569 ( .A1(G237), .A2(G234), .ZN(n451) );
  XNOR2_X1 U570 ( .A(n451), .B(KEYINPUT14), .ZN(n452) );
  XNOR2_X1 U571 ( .A(KEYINPUT74), .B(n452), .ZN(n453) );
  NAND2_X1 U572 ( .A1(G952), .A2(n453), .ZN(n688) );
  NOR2_X1 U573 ( .A1(n688), .A2(G953), .ZN(n564) );
  NAND2_X1 U574 ( .A1(n453), .A2(G902), .ZN(n562) );
  OR2_X1 U575 ( .A1(n738), .A2(n562), .ZN(n454) );
  NOR2_X1 U576 ( .A1(G900), .A2(n454), .ZN(n455) );
  NOR2_X1 U577 ( .A1(n564), .A2(n455), .ZN(n520) );
  NAND2_X1 U578 ( .A1(n508), .A2(G210), .ZN(n456) );
  XNOR2_X1 U579 ( .A(n457), .B(n456), .ZN(n461) );
  XNOR2_X1 U580 ( .A(n462), .B(KEYINPUT3), .ZN(n464) );
  XNOR2_X1 U581 ( .A(n464), .B(n463), .ZN(n485) );
  XNOR2_X1 U582 ( .A(n465), .B(n485), .ZN(n466) );
  XNOR2_X1 U583 ( .A(n467), .B(n466), .ZN(n468) );
  INV_X1 U584 ( .A(G902), .ZN(n473) );
  XNOR2_X1 U585 ( .A(KEYINPUT94), .B(G472), .ZN(n470) );
  XNOR2_X2 U586 ( .A(n471), .B(n470), .ZN(n666) );
  NAND2_X1 U587 ( .A1(n473), .A2(n472), .ZN(n490) );
  NAND2_X1 U588 ( .A1(n490), .A2(G214), .ZN(n672) );
  NAND2_X1 U589 ( .A1(n666), .A2(n672), .ZN(n474) );
  XNOR2_X1 U590 ( .A(n475), .B(n476), .ZN(n480) );
  NAND2_X1 U591 ( .A1(n738), .A2(G224), .ZN(n477) );
  XNOR2_X1 U592 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U593 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U594 ( .A(n482), .B(n481), .ZN(n488) );
  XNOR2_X1 U595 ( .A(n497), .B(KEYINPUT16), .ZN(n487) );
  INV_X1 U596 ( .A(n485), .ZN(n486) );
  XNOR2_X1 U597 ( .A(n488), .B(n722), .ZN(n614) );
  INV_X1 U598 ( .A(n489), .ZN(n601) );
  OR2_X2 U599 ( .A1(n614), .A2(n601), .ZN(n492) );
  AND2_X1 U600 ( .A1(n490), .A2(G210), .ZN(n491) );
  XOR2_X1 U601 ( .A(KEYINPUT101), .B(KEYINPUT9), .Z(n495) );
  XNOR2_X1 U602 ( .A(n495), .B(KEYINPUT7), .ZN(n496) );
  XOR2_X1 U603 ( .A(n497), .B(n496), .Z(n498) );
  NAND2_X1 U604 ( .A1(G217), .A2(n499), .ZN(n500) );
  XNOR2_X1 U605 ( .A(n502), .B(n501), .ZN(n506) );
  XNOR2_X1 U606 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U607 ( .A(n506), .B(n505), .ZN(n511) );
  NAND2_X1 U608 ( .A1(n541), .A2(n542), .ZN(n572) );
  INV_X1 U609 ( .A(n541), .ZN(n516) );
  NOR2_X1 U610 ( .A1(n516), .A2(n515), .ZN(n645) );
  NAND2_X1 U611 ( .A1(n678), .A2(KEYINPUT47), .ZN(n517) );
  XOR2_X1 U612 ( .A(KEYINPUT80), .B(n517), .Z(n518) );
  INV_X1 U613 ( .A(n666), .ZN(n586) );
  NOR2_X1 U614 ( .A1(n520), .A2(n661), .ZN(n521) );
  NAND2_X1 U615 ( .A1(n521), .A2(n568), .ZN(n530) );
  XNOR2_X1 U616 ( .A(KEYINPUT28), .B(n522), .ZN(n523) );
  NAND2_X1 U617 ( .A1(n523), .A2(n529), .ZN(n546) );
  XOR2_X1 U618 ( .A(n526), .B(KEYINPUT47), .Z(n528) );
  NAND2_X1 U619 ( .A1(n526), .A2(n678), .ZN(n527) );
  NAND2_X1 U620 ( .A1(n528), .A2(n527), .ZN(n534) );
  XNOR2_X1 U621 ( .A(n666), .B(KEYINPUT6), .ZN(n580) );
  INV_X1 U622 ( .A(n580), .ZN(n531) );
  NAND2_X1 U623 ( .A1(n672), .A2(n531), .ZN(n532) );
  XNOR2_X1 U624 ( .A(n748), .B(KEYINPUT83), .ZN(n533) );
  NAND2_X1 U625 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U626 ( .A(n538), .B(n537), .ZN(n554) );
  INV_X1 U627 ( .A(KEYINPUT38), .ZN(n539) );
  NOR2_X1 U628 ( .A1(n542), .A2(n541), .ZN(n544) );
  INV_X1 U629 ( .A(KEYINPUT102), .ZN(n543) );
  XNOR2_X1 U630 ( .A(n544), .B(n543), .ZN(n676) );
  XNOR2_X1 U631 ( .A(n545), .B(KEYINPUT41), .ZN(n654) );
  NAND2_X1 U632 ( .A1(n547), .A2(n673), .ZN(n548) );
  XNOR2_X1 U633 ( .A(n548), .B(KEYINPUT39), .ZN(n556) );
  AND2_X1 U634 ( .A1(n556), .A2(n355), .ZN(n549) );
  XNOR2_X1 U635 ( .A(n549), .B(KEYINPUT40), .ZN(n743) );
  NAND2_X1 U636 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U637 ( .A(n552), .B(KEYINPUT46), .ZN(n553) );
  NOR2_X2 U638 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X2 U639 ( .A(n555), .B(KEYINPUT48), .ZN(n608) );
  NAND2_X1 U640 ( .A1(n556), .A2(n645), .ZN(n648) );
  NAND2_X1 U641 ( .A1(n581), .A2(n384), .ZN(n557) );
  XNOR2_X1 U642 ( .A(n557), .B(KEYINPUT43), .ZN(n559) );
  NAND2_X1 U643 ( .A1(n559), .A2(n558), .ZN(n631) );
  AND2_X1 U644 ( .A1(n648), .A2(n631), .ZN(n560) );
  XOR2_X1 U645 ( .A(G898), .B(KEYINPUT88), .Z(n717) );
  NAND2_X1 U646 ( .A1(G953), .A2(n717), .ZN(n723) );
  NOR2_X1 U647 ( .A1(n562), .A2(n723), .ZN(n563) );
  NAND2_X1 U648 ( .A1(n565), .A2(n418), .ZN(n567) );
  XNOR2_X1 U649 ( .A(KEYINPUT66), .B(KEYINPUT0), .ZN(n566) );
  AND2_X1 U650 ( .A1(n660), .A2(n586), .ZN(n569) );
  INV_X1 U651 ( .A(n638), .ZN(n575) );
  XNOR2_X1 U652 ( .A(n570), .B(KEYINPUT33), .ZN(n681) );
  NOR2_X1 U653 ( .A1(n681), .A2(n588), .ZN(n571) );
  XNOR2_X1 U654 ( .A(n571), .B(KEYINPUT34), .ZN(n574) );
  INV_X1 U655 ( .A(n572), .ZN(n573) );
  NAND2_X1 U656 ( .A1(n358), .A2(n660), .ZN(n576) );
  XNOR2_X1 U657 ( .A(n576), .B(KEYINPUT103), .ZN(n577) );
  AND2_X1 U658 ( .A1(n577), .A2(n580), .ZN(n579) );
  INV_X1 U659 ( .A(KEYINPUT84), .ZN(n582) );
  XNOR2_X1 U660 ( .A(n583), .B(n582), .ZN(n585) );
  INV_X1 U661 ( .A(n660), .ZN(n584) );
  AND2_X1 U662 ( .A1(n585), .A2(n584), .ZN(n632) );
  NOR2_X1 U663 ( .A1(n364), .A2(n586), .ZN(n668) );
  INV_X1 U664 ( .A(n588), .ZN(n593) );
  NAND2_X1 U665 ( .A1(n668), .A2(n593), .ZN(n590) );
  XNOR2_X1 U666 ( .A(KEYINPUT31), .B(KEYINPUT96), .ZN(n589) );
  XNOR2_X1 U667 ( .A(n590), .B(n589), .ZN(n646) );
  NOR2_X1 U668 ( .A1(n591), .A2(n365), .ZN(n592) );
  NAND2_X1 U669 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U670 ( .A(n594), .B(KEYINPUT95), .ZN(n634) );
  OR2_X1 U671 ( .A1(n646), .A2(n634), .ZN(n596) );
  INV_X1 U672 ( .A(n678), .ZN(n595) );
  AND2_X1 U673 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U674 ( .A1(n632), .A2(n597), .ZN(n598) );
  XNOR2_X2 U675 ( .A(n599), .B(KEYINPUT45), .ZN(n604) );
  NAND2_X1 U676 ( .A1(n601), .A2(KEYINPUT2), .ZN(n602) );
  NAND2_X1 U677 ( .A1(KEYINPUT2), .A2(n648), .ZN(n605) );
  XOR2_X1 U678 ( .A(KEYINPUT78), .B(n605), .Z(n606) );
  AND2_X1 U679 ( .A1(n606), .A2(n631), .ZN(n607) );
  AND2_X1 U680 ( .A1(n608), .A2(n607), .ZN(n649) );
  NAND2_X1 U681 ( .A1(n650), .A2(n649), .ZN(n609) );
  INV_X1 U682 ( .A(KEYINPUT64), .ZN(n610) );
  XNOR2_X2 U683 ( .A(n611), .B(n610), .ZN(n708) );
  NAND2_X1 U684 ( .A1(n708), .A2(G210), .ZN(n616) );
  XNOR2_X1 U685 ( .A(KEYINPUT55), .B(KEYINPUT85), .ZN(n612) );
  XNOR2_X1 U686 ( .A(n612), .B(KEYINPUT54), .ZN(n613) );
  XNOR2_X1 U687 ( .A(n614), .B(n613), .ZN(n615) );
  XNOR2_X1 U688 ( .A(n616), .B(n615), .ZN(n618) );
  INV_X1 U689 ( .A(G952), .ZN(n617) );
  AND2_X1 U690 ( .A1(n617), .A2(G953), .ZN(n713) );
  NOR2_X2 U691 ( .A1(n618), .A2(n713), .ZN(n619) );
  XNOR2_X1 U692 ( .A(n619), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U693 ( .A1(n708), .A2(G472), .ZN(n622) );
  XNOR2_X1 U694 ( .A(n622), .B(n621), .ZN(n623) );
  NOR2_X2 U695 ( .A1(n623), .A2(n713), .ZN(n625) );
  XNOR2_X1 U696 ( .A(n625), .B(n624), .ZN(G57) );
  NAND2_X1 U697 ( .A1(n708), .A2(G478), .ZN(n627) );
  XNOR2_X1 U698 ( .A(n627), .B(n626), .ZN(n628) );
  NOR2_X2 U699 ( .A1(n628), .A2(n713), .ZN(n630) );
  XNOR2_X1 U700 ( .A(n630), .B(n629), .ZN(G63) );
  XNOR2_X1 U701 ( .A(n631), .B(n354), .ZN(G42) );
  XOR2_X1 U702 ( .A(G101), .B(n632), .Z(G3) );
  NAND2_X1 U703 ( .A1(n634), .A2(n355), .ZN(n633) );
  XNOR2_X1 U704 ( .A(n633), .B(G104), .ZN(G6) );
  XOR2_X1 U705 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n636) );
  NAND2_X1 U706 ( .A1(n634), .A2(n645), .ZN(n635) );
  XNOR2_X1 U707 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U708 ( .A(G107), .B(n637), .ZN(G9) );
  XNOR2_X1 U709 ( .A(G110), .B(n638), .ZN(G12) );
  XOR2_X1 U710 ( .A(KEYINPUT110), .B(KEYINPUT29), .Z(n640) );
  NAND2_X1 U711 ( .A1(n526), .A2(n645), .ZN(n639) );
  XNOR2_X1 U712 ( .A(n640), .B(n639), .ZN(n642) );
  XOR2_X1 U713 ( .A(G128), .B(KEYINPUT109), .Z(n641) );
  XNOR2_X1 U714 ( .A(n642), .B(n641), .ZN(G30) );
  NAND2_X1 U715 ( .A1(n526), .A2(n355), .ZN(n643) );
  XNOR2_X1 U716 ( .A(n643), .B(G146), .ZN(G48) );
  NAND2_X1 U717 ( .A1(n646), .A2(n355), .ZN(n644) );
  XNOR2_X1 U718 ( .A(n644), .B(G113), .ZN(G15) );
  NAND2_X1 U719 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U720 ( .A(n647), .B(G116), .ZN(G18) );
  XNOR2_X1 U721 ( .A(G134), .B(n648), .ZN(G36) );
  AND2_X1 U722 ( .A1(n650), .A2(n649), .ZN(n653) );
  INV_X1 U723 ( .A(n650), .ZN(n714) );
  NOR2_X1 U724 ( .A1(n714), .A2(n736), .ZN(n651) );
  NOR2_X1 U725 ( .A1(n651), .A2(KEYINPUT2), .ZN(n652) );
  NOR2_X1 U726 ( .A1(n653), .A2(n652), .ZN(n690) );
  XOR2_X1 U727 ( .A(KEYINPUT113), .B(KEYINPUT50), .Z(n658) );
  OR2_X1 U728 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U729 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U730 ( .A(KEYINPUT112), .B(n659), .ZN(n664) );
  NAND2_X1 U731 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U732 ( .A(KEYINPUT49), .B(n662), .Z(n663) );
  NAND2_X1 U733 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U734 ( .A1(n365), .A2(n665), .ZN(n667) );
  NOR2_X1 U735 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U736 ( .A(n669), .B(KEYINPUT51), .Z(n670) );
  XNOR2_X1 U737 ( .A(KEYINPUT114), .B(n670), .ZN(n671) );
  NOR2_X1 U738 ( .A1(n692), .A2(n671), .ZN(n685) );
  NOR2_X1 U739 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U740 ( .A(KEYINPUT115), .B(n674), .Z(n675) );
  NOR2_X1 U741 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U742 ( .A(n677), .B(KEYINPUT116), .ZN(n680) );
  NOR2_X1 U743 ( .A1(n680), .A2(n679), .ZN(n682) );
  NOR2_X1 U744 ( .A1(n682), .A2(n691), .ZN(n683) );
  XOR2_X1 U745 ( .A(KEYINPUT117), .B(n683), .Z(n684) );
  NOR2_X1 U746 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U747 ( .A(n686), .B(KEYINPUT52), .ZN(n687) );
  NOR2_X1 U748 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U749 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U750 ( .A(KEYINPUT53), .B(n694), .ZN(G75) );
  BUF_X1 U751 ( .A(n708), .Z(n695) );
  NAND2_X1 U752 ( .A1(n695), .A2(G469), .ZN(n701) );
  XOR2_X1 U753 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n697) );
  XNOR2_X1 U754 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n696) );
  XNOR2_X1 U755 ( .A(n697), .B(n696), .ZN(n698) );
  XOR2_X1 U756 ( .A(n699), .B(n698), .Z(n700) );
  XNOR2_X1 U757 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U758 ( .A1(n713), .A2(n702), .ZN(G54) );
  NAND2_X1 U759 ( .A1(n708), .A2(G475), .ZN(n705) );
  XNOR2_X1 U760 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X2 U761 ( .A1(n706), .A2(n713), .ZN(n707) );
  XNOR2_X1 U762 ( .A(n707), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U763 ( .A1(n695), .A2(G217), .ZN(n709) );
  NOR2_X1 U764 ( .A1(n713), .A2(n712), .ZN(G66) );
  NOR2_X1 U765 ( .A1(n714), .A2(G953), .ZN(n719) );
  NAND2_X1 U766 ( .A1(G953), .A2(G224), .ZN(n715) );
  XOR2_X1 U767 ( .A(KEYINPUT61), .B(n715), .Z(n716) );
  NOR2_X1 U768 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U769 ( .A1(n719), .A2(n718), .ZN(n726) );
  XOR2_X1 U770 ( .A(n720), .B(G101), .Z(n721) );
  XNOR2_X1 U771 ( .A(n722), .B(n721), .ZN(n724) );
  NAND2_X1 U772 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U773 ( .A(n726), .B(n725), .ZN(G69) );
  XNOR2_X1 U774 ( .A(n728), .B(n727), .ZN(n730) );
  XNOR2_X1 U775 ( .A(n729), .B(n730), .ZN(n731) );
  XOR2_X1 U776 ( .A(KEYINPUT4), .B(n731), .Z(n735) );
  XOR2_X1 U777 ( .A(G227), .B(n735), .Z(n732) );
  NAND2_X1 U778 ( .A1(n732), .A2(G900), .ZN(n733) );
  XNOR2_X1 U779 ( .A(n733), .B(KEYINPUT123), .ZN(n734) );
  NAND2_X1 U780 ( .A1(n734), .A2(G953), .ZN(n740) );
  XNOR2_X1 U781 ( .A(n736), .B(n735), .ZN(n737) );
  NAND2_X1 U782 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U783 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U784 ( .A(KEYINPUT124), .B(n741), .Z(G72) );
  XOR2_X1 U785 ( .A(G131), .B(KEYINPUT126), .Z(n742) );
  XNOR2_X1 U786 ( .A(n743), .B(n742), .ZN(G33) );
  XOR2_X1 U787 ( .A(n744), .B(n349), .Z(G45) );
  BUF_X1 U788 ( .A(n745), .Z(n746) );
  XOR2_X1 U789 ( .A(G122), .B(n746), .Z(G24) );
  XOR2_X1 U790 ( .A(KEYINPUT111), .B(KEYINPUT37), .Z(n747) );
  XNOR2_X1 U791 ( .A(n748), .B(n747), .ZN(n749) );
  XNOR2_X1 U792 ( .A(G125), .B(n749), .ZN(G27) );
  XOR2_X1 U793 ( .A(G137), .B(n750), .Z(G39) );
endmodule

