//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0 1 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n551,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n607, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1189, new_n1190, new_n1191;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(G125), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n461), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  OAI211_X1 g044(.A(G137), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n466), .A2(new_n471), .ZN(G160));
  INV_X1    g047(.A(new_n462), .ZN(new_n473));
  INV_X1    g048(.A(new_n463), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n461), .B1(new_n473), .B2(new_n474), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n476), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  OAI211_X1 g057(.A(G138), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT4), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g062(.A(KEYINPUT3), .B(G2104), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n488), .A2(G138), .A3(new_n461), .A4(new_n485), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g065(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n492), .A2(new_n494), .A3(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT67), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT67), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n491), .A2(new_n498), .A3(new_n495), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n490), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  XNOR2_X1  g076(.A(KEYINPUT5), .B(G543), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OR2_X1    g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n509), .A2(new_n510), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n505), .A2(new_n517), .ZN(G166));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  INV_X1    g095(.A(G89), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n520), .B1(new_n521), .B2(new_n515), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n522), .A2(KEYINPUT69), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(KEYINPUT69), .ZN(new_n524));
  INV_X1    g099(.A(G543), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n525), .B1(new_n506), .B2(new_n507), .ZN(new_n526));
  AND2_X1   g101(.A1(G63), .A2(G651), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n526), .A2(G51), .B1(new_n502), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n523), .A2(new_n524), .A3(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(G168));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n512), .A2(new_n511), .ZN(new_n532));
  INV_X1    g107(.A(G64), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT70), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n504), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n536), .B1(new_n535), .B2(new_n534), .ZN(new_n537));
  INV_X1    g112(.A(new_n515), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n538), .A2(G90), .B1(G52), .B2(new_n526), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  AOI22_X1  g116(.A1(new_n502), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n504), .ZN(new_n543));
  INV_X1    g118(.A(G43), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n509), .A2(new_n544), .B1(new_n515), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n549));
  XOR2_X1   g124(.A(new_n549), .B(KEYINPUT71), .Z(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT72), .ZN(G188));
  INV_X1    g129(.A(KEYINPUT73), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n515), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n508), .A2(new_n502), .A3(KEYINPUT73), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n556), .A2(G91), .A3(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n526), .A2(new_n559), .A3(G53), .ZN(new_n560));
  OAI211_X1 g135(.A(G53), .B(G543), .C1(new_n513), .C2(new_n514), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n532), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G651), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n558), .A2(new_n563), .A3(new_n567), .ZN(G299));
  INV_X1    g143(.A(KEYINPUT74), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n529), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n523), .A2(KEYINPUT74), .A3(new_n524), .A4(new_n528), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G286));
  OR2_X1    g148(.A1(new_n505), .A2(new_n517), .ZN(G303));
  NAND3_X1  g149(.A1(new_n556), .A2(G87), .A3(new_n557), .ZN(new_n575));
  INV_X1    g150(.A(G74), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n532), .A2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G651), .B1(new_n526), .B2(G49), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n575), .A2(new_n578), .ZN(G288));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n532), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(G48), .B2(new_n526), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n556), .A2(G86), .A3(new_n557), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G305));
  AOI22_X1  g160(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(new_n504), .ZN(new_n587));
  INV_X1    g162(.A(G47), .ZN(new_n588));
  INV_X1    g163(.A(G85), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n509), .A2(new_n588), .B1(new_n515), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n556), .A2(G92), .A3(new_n557), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n532), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G651), .B1(G54), .B2(new_n526), .ZN(new_n600));
  AND2_X1   g175(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n593), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n593), .B1(new_n601), .B2(G868), .ZN(G321));
  NOR2_X1   g178(.A1(G299), .A2(G868), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n604), .B1(new_n572), .B2(G868), .ZN(G297));
  AOI21_X1  g180(.A(new_n604), .B1(new_n572), .B2(G868), .ZN(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n601), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND2_X1  g183(.A1(new_n596), .A2(new_n600), .ZN(new_n609));
  OAI21_X1  g184(.A(G868), .B1(new_n609), .B2(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n488), .A2(new_n468), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT13), .Z(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G2100), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT75), .Z(new_n617));
  NAND2_X1  g192(.A1(new_n477), .A2(G123), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n475), .A2(G135), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT76), .ZN(new_n620));
  NOR3_X1   g195(.A1(new_n620), .A2(new_n461), .A3(G111), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n461), .B2(G111), .ZN(new_n622));
  OR2_X1    g197(.A1(G99), .A2(G2105), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n622), .A2(G2104), .A3(new_n623), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n618), .B(new_n619), .C1(new_n621), .C2(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(G2096), .Z(new_n626));
  OAI211_X1 g201(.A(new_n617), .B(new_n626), .C1(G2100), .C2(new_n615), .ZN(G156));
  XNOR2_X1  g202(.A(G2427), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2430), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n631), .A2(KEYINPUT14), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n635), .A2(new_n637), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2451), .B(G2454), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT77), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n638), .A2(new_n643), .A3(new_n639), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(G14), .A3(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(G401));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2072), .B(G2078), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(KEYINPUT78), .B(KEYINPUT18), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n650), .A2(new_n651), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n655), .A2(new_n649), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT79), .Z(new_n657));
  XOR2_X1   g232(.A(new_n651), .B(KEYINPUT17), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n654), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n649), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n650), .B1(new_n657), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2096), .B(G2100), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT19), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  AND2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n669), .A2(new_n670), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  MUX2_X1   g251(.A(new_n676), .B(new_n675), .S(new_n668), .Z(new_n677));
  NOR2_X1   g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(G1981), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n678), .B(G1981), .ZN(new_n685));
  INV_X1    g260(.A(new_n683), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  INV_X1    g263(.A(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  AND3_X1   g265(.A1(new_n684), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n690), .B1(new_n684), .B2(new_n687), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(G229));
  NAND2_X1  g268(.A1(new_n475), .A2(G139), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT91), .B(KEYINPUT25), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n694), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT92), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n488), .A2(G127), .ZN(new_n701));
  AND2_X1   g276(.A1(G115), .A2(G2104), .ZN(new_n702));
  OAI21_X1  g277(.A(G2105), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  MUX2_X1   g279(.A(G33), .B(new_n704), .S(G29), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G2072), .ZN(new_n706));
  INV_X1    g281(.A(new_n547), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT82), .B(G16), .Z(new_n708));
  MUX2_X1   g283(.A(new_n707), .B(G19), .S(new_n708), .Z(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G1341), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G26), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT28), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n475), .A2(G140), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n477), .A2(G128), .ZN(new_n715));
  OR2_X1    g290(.A1(G104), .A2(G2105), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n716), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n714), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n713), .B1(new_n719), .B2(new_n711), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT90), .B(G2067), .Z(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT31), .B(G11), .Z(new_n723));
  NOR2_X1   g298(.A1(new_n625), .A2(new_n711), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT30), .B(G28), .ZN(new_n725));
  AOI211_X1 g300(.A(new_n723), .B(new_n724), .C1(new_n711), .C2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT24), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n711), .B1(new_n727), .B2(G34), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n727), .B2(G34), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G160), .B2(G29), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G2084), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n710), .A2(new_n722), .A3(new_n726), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n720), .A2(new_n721), .ZN(new_n733));
  OAI221_X1 g308(.A(new_n733), .B1(G2084), .B2(new_n730), .C1(new_n709), .C2(G1341), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(G29), .A2(G35), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G162), .B2(G29), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G2090), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n741), .A2(KEYINPUT95), .ZN(new_n742));
  MUX2_X1   g317(.A(G21), .B(new_n529), .S(G16), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G1966), .ZN(new_n744));
  NOR4_X1   g319(.A1(new_n706), .A2(new_n735), .A3(new_n742), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n711), .A2(G32), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n475), .A2(G141), .ZN(new_n747));
  INV_X1    g322(.A(G105), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(new_n467), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n477), .A2(G129), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT26), .Z(new_n752));
  NAND2_X1  g327(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n746), .B1(new_n754), .B2(new_n711), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT93), .Z(new_n756));
  XOR2_X1   g331(.A(KEYINPUT27), .B(G1996), .Z(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(G164), .A2(new_n711), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G27), .B2(new_n711), .ZN(new_n760));
  INV_X1    g335(.A(G2078), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  INV_X1    g338(.A(G5), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(G16), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G301), .B2(G16), .ZN(new_n766));
  INV_X1    g341(.A(G1961), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n758), .A2(new_n762), .A3(new_n763), .A4(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n766), .A2(new_n767), .ZN(new_n770));
  OAI221_X1 g345(.A(new_n770), .B1(new_n740), .B2(new_n739), .C1(new_n756), .C2(new_n757), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(G299), .A2(G16), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n708), .A2(G20), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT23), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT96), .ZN(new_n777));
  INV_X1    g352(.A(G1956), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G4), .A2(G16), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT87), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n601), .B2(G16), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT89), .B(G1348), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT88), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n782), .A2(new_n784), .ZN(new_n786));
  AOI211_X1 g361(.A(new_n785), .B(new_n786), .C1(KEYINPUT95), .C2(new_n741), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n745), .A2(new_n772), .A3(new_n779), .A4(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(G6), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n789), .A2(G16), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G305), .B2(G16), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT32), .B(G1981), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n791), .B(new_n792), .Z(new_n793));
  INV_X1    g368(.A(G22), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n708), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G303), .B2(new_n708), .ZN(new_n796));
  INV_X1    g371(.A(G1971), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  MUX2_X1   g374(.A(G23), .B(G288), .S(G16), .Z(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(KEYINPUT85), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(KEYINPUT85), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT33), .B(G1976), .Z(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n801), .A2(new_n804), .A3(new_n802), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n799), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(KEYINPUT86), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT86), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n799), .A2(new_n806), .A3(new_n810), .A4(new_n807), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT84), .B(KEYINPUT34), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n813), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n809), .A2(new_n811), .A3(new_n815), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n591), .B(KEYINPUT83), .Z(new_n817));
  MUX2_X1   g392(.A(new_n817), .B(G24), .S(new_n708), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(G1986), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n711), .A2(G25), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n475), .A2(G131), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n477), .A2(G119), .ZN(new_n822));
  OR2_X1    g397(.A1(G95), .A2(G2105), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n823), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n821), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n820), .B1(new_n826), .B2(new_n711), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT35), .B(G1991), .Z(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n827), .B(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n819), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n814), .A2(new_n816), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(KEYINPUT36), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT36), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n814), .A2(new_n834), .A3(new_n816), .A4(new_n831), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n788), .B1(new_n833), .B2(new_n835), .ZN(G311));
  INV_X1    g411(.A(KEYINPUT97), .ZN(new_n837));
  XNOR2_X1  g412(.A(G311), .B(new_n837), .ZN(G150));
  AOI22_X1  g413(.A1(new_n502), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n839), .A2(new_n504), .ZN(new_n840));
  INV_X1    g415(.A(G55), .ZN(new_n841));
  INV_X1    g416(.A(G93), .ZN(new_n842));
  OAI22_X1  g417(.A1(new_n509), .A2(new_n841), .B1(new_n515), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(G860), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT37), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n601), .A2(G559), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT38), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n840), .A2(new_n843), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n547), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n847), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT98), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(KEYINPUT98), .B1(new_n850), .B2(new_n851), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(G860), .B1(new_n850), .B2(new_n851), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n845), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(G145));
  XNOR2_X1  g435(.A(new_n754), .B(new_n718), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n496), .B1(new_n489), .B2(new_n487), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n700), .A2(new_n703), .A3(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n862), .B1(new_n700), .B2(new_n703), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n861), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n865), .ZN(new_n867));
  INV_X1    g442(.A(new_n861), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(new_n868), .A3(new_n863), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n475), .A2(G142), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n477), .A2(G130), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n461), .A2(G118), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n871), .B(new_n872), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n614), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n876), .A2(new_n826), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n826), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT100), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n877), .A2(KEYINPUT100), .A3(new_n878), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n870), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n481), .B(G160), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n625), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n866), .A2(new_n869), .A3(new_n880), .A4(new_n879), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n883), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n885), .B1(new_n883), .B2(new_n886), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g467(.A(KEYINPUT103), .ZN(new_n893));
  NAND2_X1  g468(.A1(G303), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(G166), .A2(KEYINPUT103), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(G290), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(G290), .B1(new_n894), .B2(new_n895), .ZN(new_n898));
  AOI21_X1  g473(.A(G288), .B1(new_n584), .B2(new_n583), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n575), .A2(new_n578), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n900), .A2(G305), .ZN(new_n901));
  OAI22_X1  g476(.A1(new_n897), .A2(new_n898), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n898), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n901), .A2(new_n899), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(new_n904), .A3(new_n896), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT104), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n902), .A2(new_n905), .A3(KEYINPUT104), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(KEYINPUT105), .A3(KEYINPUT42), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT42), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT105), .B1(new_n906), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n914), .B1(new_n910), .B2(new_n913), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n609), .A2(G559), .ZN(new_n916));
  INV_X1    g491(.A(new_n849), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n916), .B(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT101), .ZN(new_n919));
  NAND2_X1  g494(.A1(G299), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g495(.A1(G299), .A2(new_n919), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n601), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n609), .A2(new_n919), .A3(G299), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n918), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g500(.A(KEYINPUT102), .B(KEYINPUT41), .Z(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(KEYINPUT41), .B2(new_n924), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n925), .B1(new_n929), .B2(new_n918), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n912), .A2(new_n915), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n930), .B1(new_n912), .B2(new_n915), .ZN(new_n932));
  OAI21_X1  g507(.A(G868), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(G868), .B2(new_n848), .ZN(G295));
  OAI21_X1  g509(.A(new_n933), .B1(G868), .B2(new_n848), .ZN(G331));
  AOI21_X1  g510(.A(G301), .B1(new_n570), .B2(new_n571), .ZN(new_n936));
  NOR2_X1   g511(.A1(G168), .A2(G171), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n849), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n939), .A2(new_n924), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n936), .A2(new_n937), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n917), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n924), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n927), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(KEYINPUT41), .B2(new_n944), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT106), .B1(new_n941), .B2(new_n917), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n948));
  NOR4_X1   g523(.A1(new_n936), .A2(new_n937), .A3(new_n948), .A4(new_n849), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n947), .A2(new_n939), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n943), .B1(new_n946), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n910), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n947), .A2(new_n949), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n940), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n942), .A2(new_n938), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n929), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n954), .A2(new_n911), .A3(new_n956), .ZN(new_n957));
  AND4_X1   g532(.A1(KEYINPUT43), .A2(new_n952), .A3(new_n888), .A4(new_n957), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n953), .A2(new_n940), .B1(new_n929), .B2(new_n955), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(new_n911), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(G37), .B1(new_n959), .B2(new_n911), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT43), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT44), .B1(new_n958), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n957), .A2(new_n888), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT43), .B1(new_n965), .B2(new_n960), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT43), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n962), .A2(new_n952), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n964), .B1(new_n970), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n972), .B1(new_n862), .B2(G1384), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n464), .A2(new_n465), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(G2105), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n975), .A2(G40), .A3(new_n469), .A4(new_n470), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G2067), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n718), .B(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G1996), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(G1996), .B1(new_n749), .B2(new_n753), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n980), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n977), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n985), .B(KEYINPUT107), .Z(new_n986));
  NOR2_X1   g561(.A1(new_n825), .A2(new_n829), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n719), .A2(new_n979), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n978), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT126), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n990), .A2(new_n991), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n978), .B1(new_n754), .B2(new_n980), .ZN(new_n994));
  OR3_X1    g569(.A1(new_n978), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT46), .B1(new_n978), .B2(G1996), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  XOR2_X1   g572(.A(new_n997), .B(KEYINPUT47), .Z(new_n998));
  NOR2_X1   g573(.A1(new_n826), .A2(new_n828), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n977), .B1(new_n987), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n986), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n977), .A2(new_n689), .A3(new_n591), .ZN(new_n1002));
  XOR2_X1   g577(.A(new_n1002), .B(KEYINPUT48), .Z(new_n1003));
  OAI21_X1  g578(.A(new_n998), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n992), .A2(new_n993), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n1006));
  INV_X1    g581(.A(G1384), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n500), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G40), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n466), .A2(new_n471), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n496), .ZN(new_n1011));
  AOI21_X1  g586(.A(G1384), .B1(new_n490), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1010), .B1(new_n1012), .B2(new_n1006), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n778), .B1(new_n1008), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n976), .B1(new_n1012), .B2(KEYINPUT45), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT56), .B(G2072), .ZN(new_n1016));
  AOI22_X1  g591(.A1(new_n489), .A2(new_n487), .B1(new_n496), .B2(KEYINPUT67), .ZN(new_n1017));
  AOI21_X1  g592(.A(G1384), .B1(new_n1017), .B2(new_n499), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1015), .B(new_n1016), .C1(KEYINPUT45), .C2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT118), .ZN(new_n1020));
  OR2_X1    g595(.A1(new_n1020), .A2(KEYINPUT57), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n558), .A2(new_n563), .A3(new_n567), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1020), .A2(KEYINPUT57), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1014), .A2(new_n1019), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  AOI211_X1 g601(.A(KEYINPUT50), .B(G1384), .C1(new_n490), .C2(new_n1011), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n1028));
  OAI22_X1  g603(.A1(new_n1018), .A2(new_n1006), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n500), .A2(new_n1007), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1030), .A2(KEYINPUT109), .A3(KEYINPUT50), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(new_n1010), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n783), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1012), .A2(new_n979), .A3(new_n1010), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n609), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1024), .B1(new_n1014), .B2(new_n1019), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1026), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(new_n1025), .B2(new_n1036), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT61), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT61), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1038), .B(new_n1041), .C1(new_n1025), .C2(new_n1036), .ZN(new_n1042));
  OR2_X1    g617(.A1(new_n601), .A2(KEYINPUT60), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1033), .A2(new_n1043), .A3(new_n1034), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n596), .A2(KEYINPUT60), .A3(new_n600), .ZN(new_n1045));
  XOR2_X1   g620(.A(new_n1045), .B(KEYINPUT121), .Z(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1040), .A2(new_n1042), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1030), .A2(new_n972), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1050), .A2(new_n981), .A3(new_n1015), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1012), .A2(new_n1010), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1053), .B(G1341), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1049), .B1(new_n1056), .B2(new_n547), .ZN(new_n1057));
  AOI211_X1 g632(.A(KEYINPUT59), .B(new_n707), .C1(new_n1051), .C2(new_n1055), .ZN(new_n1058));
  OAI22_X1  g633(.A1(new_n1044), .A2(new_n1046), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1037), .B1(new_n1048), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1032), .A2(new_n767), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT116), .B1(new_n1018), .B2(KEYINPUT45), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n973), .A2(new_n1010), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n500), .A2(KEYINPUT116), .A3(KEYINPUT45), .A4(new_n1007), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1066), .A2(G2078), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .A4(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1050), .A2(new_n1015), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1066), .B1(new_n1069), .B2(G2078), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1061), .A2(new_n1068), .A3(G301), .A4(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT123), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n1071), .B(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1012), .A2(KEYINPUT45), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1064), .A2(new_n1075), .A3(new_n1067), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1061), .A2(new_n1070), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1074), .B1(new_n1077), .B2(G171), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1073), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1966), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1065), .A2(new_n1010), .A3(new_n973), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(new_n1081), .B2(new_n1062), .ZN(new_n1082));
  INV_X1    g657(.A(G2084), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1029), .A2(new_n1083), .A3(new_n1010), .A4(new_n1031), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n529), .A2(G8), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT51), .B1(new_n1087), .B2(KEYINPUT122), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1085), .A2(G8), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1089), .B1(new_n1090), .B2(new_n1086), .ZN(new_n1091));
  INV_X1    g666(.A(G8), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1092), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1089), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1093), .A2(new_n1094), .A3(new_n1087), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1088), .B1(new_n1091), .B2(new_n1095), .ZN(new_n1096));
  XOR2_X1   g671(.A(KEYINPUT110), .B(G2090), .Z(new_n1097));
  NAND4_X1  g672(.A1(new_n1029), .A2(new_n1010), .A3(new_n1031), .A4(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(G1971), .B1(new_n1050), .B2(new_n1015), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1092), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(G303), .A2(G8), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(KEYINPUT55), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1092), .B1(new_n1012), .B2(new_n1010), .ZN(new_n1106));
  INV_X1    g681(.A(G1976), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT52), .B1(G288), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n575), .A2(G1976), .A3(new_n578), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1106), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT112), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT112), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1106), .A2(new_n1108), .A3(new_n1112), .A4(new_n1109), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1052), .A2(G8), .A3(new_n1109), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT111), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1106), .A2(KEYINPUT111), .A3(new_n1109), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1117), .A2(KEYINPUT52), .A3(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT113), .B(G1981), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n583), .A2(new_n584), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n526), .A2(G48), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n508), .A2(new_n502), .A3(G86), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n502), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1122), .B(new_n1123), .C1(new_n1124), .C2(new_n504), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(G1981), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1121), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT49), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1121), .A2(new_n1126), .A3(KEYINPUT49), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1129), .A2(new_n1106), .A3(new_n1130), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1114), .A2(new_n1119), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1097), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1008), .A2(new_n1013), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(G8), .B1(new_n1134), .B2(new_n1099), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n1103), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1105), .A2(new_n1132), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1061), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(G171), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1061), .A2(G301), .A3(new_n1070), .A4(new_n1076), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1137), .B1(new_n1141), .B2(new_n1074), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1060), .A2(new_n1079), .A3(new_n1096), .A4(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT117), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1114), .A2(new_n1119), .A3(new_n1131), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1144), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1132), .B(KEYINPUT117), .C1(new_n1104), .C2(new_n1101), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1093), .A2(new_n572), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT63), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1151), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .A4(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1151), .B1(new_n1137), .B2(new_n1149), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1131), .A2(new_n1107), .A3(new_n900), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n1121), .ZN(new_n1156));
  XOR2_X1   g731(.A(new_n1106), .B(KEYINPUT114), .Z(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1158), .B1(new_n1105), .B2(new_n1146), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT115), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1158), .B(KEYINPUT115), .C1(new_n1105), .C2(new_n1146), .ZN(new_n1162));
  AOI22_X1  g737(.A1(new_n1153), .A2(new_n1154), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1143), .A2(new_n1163), .A3(KEYINPUT124), .ZN(new_n1164));
  AOI21_X1  g739(.A(KEYINPUT124), .B1(new_n1143), .B2(new_n1163), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT62), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1088), .B(new_n1166), .C1(new_n1091), .C2(new_n1095), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT125), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1168), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n1096), .A2(KEYINPUT62), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NOR3_X1   g748(.A1(new_n1164), .A2(new_n1165), .A3(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n591), .B(new_n689), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1001), .B1(new_n977), .B2(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT108), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1005), .B1(new_n1174), .B2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g753(.A(G229), .ZN(new_n1180));
  NOR2_X1   g754(.A1(G227), .A2(new_n459), .ZN(new_n1181));
  AND2_X1   g755(.A1(new_n647), .A2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g756(.A(new_n1180), .B(new_n1182), .C1(new_n890), .C2(new_n889), .ZN(new_n1183));
  AOI211_X1 g757(.A(KEYINPUT127), .B(new_n1183), .C1(new_n966), .C2(new_n968), .ZN(new_n1184));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n1185));
  INV_X1    g759(.A(new_n1183), .ZN(new_n1186));
  AOI21_X1  g760(.A(new_n1185), .B1(new_n969), .B2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g761(.A1(new_n1184), .A2(new_n1187), .ZN(G308));
  NAND2_X1  g762(.A1(new_n969), .A2(new_n1186), .ZN(new_n1189));
  NAND2_X1  g763(.A1(new_n1189), .A2(KEYINPUT127), .ZN(new_n1190));
  NAND3_X1  g764(.A1(new_n969), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1191));
  NAND2_X1  g765(.A1(new_n1190), .A2(new_n1191), .ZN(G225));
endmodule


