//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n801, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1029, new_n1030, new_n1031, new_n1032;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n203), .A2(KEYINPUT91), .ZN(new_n204));
  OAI21_X1  g003(.A(KEYINPUT92), .B1(new_n202), .B2(KEYINPUT15), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(KEYINPUT91), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n208));
  INV_X1    g007(.A(G36gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT93), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n212), .A2(new_n213), .B1(G29gat), .B2(G36gat), .ZN(new_n214));
  OR3_X1    g013(.A1(new_n202), .A2(KEYINPUT92), .A3(KEYINPUT15), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n210), .A2(KEYINPUT93), .A3(new_n211), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n211), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n218), .B1(KEYINPUT90), .B2(new_n210), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n210), .A2(KEYINPUT90), .ZN(new_n220));
  AOI22_X1  g019(.A1(new_n219), .A2(new_n220), .B1(G29gat), .B2(G36gat), .ZN(new_n221));
  OAI22_X1  g020(.A1(new_n207), .A2(new_n217), .B1(new_n203), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT17), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G15gat), .B(G22gat), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n225), .A2(G1gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT16), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n225), .B1(new_n227), .B2(G1gat), .ZN(new_n228));
  INV_X1    g027(.A(G8gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n230), .B(KEYINPUT96), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n226), .A2(new_n228), .A3(KEYINPUT95), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n232), .B(G8gat), .C1(KEYINPUT95), .C2(new_n226), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n224), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT94), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n222), .A2(new_n236), .ZN(new_n237));
  OAI221_X1 g036(.A(KEYINPUT94), .B1(new_n203), .B2(new_n221), .C1(new_n207), .C2(new_n217), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(new_n223), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G229gat), .A2(G233gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n237), .A2(new_n234), .A3(new_n238), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT18), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n240), .A2(KEYINPUT18), .A3(new_n241), .A4(new_n242), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n237), .A2(new_n238), .ZN(new_n247));
  INV_X1    g046(.A(new_n234), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(new_n242), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n241), .B(KEYINPUT13), .Z(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n245), .A2(new_n246), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G113gat), .B(G141gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT89), .B(G197gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XOR2_X1   g055(.A(KEYINPUT11), .B(G169gat), .Z(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT12), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n253), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n245), .A2(new_n246), .A3(new_n252), .A4(new_n259), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n261), .A2(KEYINPUT97), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT97), .B1(new_n261), .B2(new_n262), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT22), .ZN(new_n267));
  INV_X1    g066(.A(G211gat), .ZN(new_n268));
  INV_X1    g067(.A(G218gat), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT74), .B(G197gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n271), .A2(G204gat), .ZN(new_n272));
  INV_X1    g071(.A(G197gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT74), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT74), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(G197gat), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n274), .A2(new_n276), .A3(G204gat), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n270), .B1(new_n272), .B2(new_n277), .ZN(new_n278));
  XOR2_X1   g077(.A(G211gat), .B(G218gat), .Z(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n279), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n274), .A2(new_n276), .ZN(new_n282));
  INV_X1    g081(.A(G204gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n271), .A2(G204gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n281), .B1(new_n286), .B2(new_n270), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n280), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT75), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT29), .ZN(new_n290));
  NOR2_X1   g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT65), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT23), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n292), .A2(new_n293), .B1(G169gat), .B2(G176gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n291), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G176gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT23), .ZN(new_n298));
  AND2_X1   g097(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n300));
  NOR3_X1   g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT66), .B1(new_n296), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G169gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(new_n297), .ZN(new_n304));
  NAND2_X1  g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n305), .B1(KEYINPUT65), .B2(KEYINPUT23), .ZN(new_n306));
  INV_X1    g105(.A(new_n295), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT66), .ZN(new_n309));
  INV_X1    g108(.A(new_n300), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n293), .A2(G176gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n308), .A2(new_n309), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G190gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n315), .A2(G183gat), .ZN(new_n316));
  INV_X1    g115(.A(G183gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(G190gat), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT24), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G183gat), .A2(G190gat), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n320), .A2(KEYINPUT24), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n302), .A2(new_n314), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT25), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT67), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n325), .B1(new_n319), .B2(new_n321), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n324), .B1(new_n311), .B2(new_n303), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n308), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n319), .A2(new_n325), .A3(new_n321), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n323), .A2(new_n324), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n303), .A2(new_n297), .A3(KEYINPUT26), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT26), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n333), .B1(G169gat), .B2(G176gat), .ZN(new_n334));
  INV_X1    g133(.A(new_n305), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n332), .B(new_n320), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n317), .A2(KEYINPUT27), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT27), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(G183gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n337), .A2(new_n339), .A3(new_n315), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT28), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n337), .A2(new_n339), .A3(KEYINPUT28), .A4(new_n315), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n336), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(KEYINPUT68), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n290), .B1(new_n331), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G226gat), .A2(G233gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n347), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n349), .B1(new_n331), .B2(new_n344), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n289), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT68), .ZN(new_n352));
  AOI211_X1 g151(.A(new_n352), .B(new_n336), .C1(new_n342), .C2(new_n343), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n342), .A2(new_n343), .ZN(new_n354));
  INV_X1    g153(.A(new_n336), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT68), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n319), .A2(new_n321), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n308), .A2(new_n313), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n358), .B1(new_n359), .B2(KEYINPUT66), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT25), .B1(new_n360), .B2(new_n314), .ZN(new_n361));
  INV_X1    g160(.A(new_n330), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n362), .A2(new_n326), .A3(new_n328), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n357), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n349), .B1(new_n364), .B2(new_n290), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n365), .A2(KEYINPUT75), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n288), .B1(new_n351), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT76), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n290), .B1(new_n331), .B2(new_n344), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n368), .B1(new_n369), .B2(new_n347), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n288), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n364), .A2(new_n349), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n323), .A2(new_n324), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n329), .A2(new_n330), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n344), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n368), .B(new_n347), .C1(new_n376), .C2(KEYINPUT29), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n371), .A2(new_n372), .A3(new_n373), .A4(new_n377), .ZN(new_n378));
  XOR2_X1   g177(.A(G8gat), .B(G36gat), .Z(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT77), .ZN(new_n380));
  XNOR2_X1  g179(.A(G64gat), .B(G92gat), .ZN(new_n381));
  XOR2_X1   g180(.A(new_n380), .B(new_n381), .Z(new_n382));
  NAND4_X1  g181(.A1(new_n367), .A2(new_n378), .A3(KEYINPUT30), .A4(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n382), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n376), .A2(new_n347), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT75), .B1(new_n365), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n348), .A2(new_n289), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n372), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n377), .A2(new_n373), .ZN(new_n389));
  NOR3_X1   g188(.A1(new_n389), .A2(new_n288), .A3(new_n370), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n384), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT78), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n383), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n388), .A2(new_n390), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n394), .A2(KEYINPUT78), .A3(KEYINPUT30), .A4(new_n382), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT79), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n367), .A2(new_n378), .A3(new_n382), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT30), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G1gat), .B(G29gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(KEYINPUT0), .ZN(new_n404));
  XNOR2_X1  g203(.A(G57gat), .B(G85gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n404), .B(new_n405), .Z(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  XOR2_X1   g206(.A(G141gat), .B(G148gat), .Z(new_n408));
  INV_X1    g207(.A(G155gat), .ZN(new_n409));
  INV_X1    g208(.A(G162gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(G155gat), .A2(G162gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(KEYINPUT2), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n408), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G141gat), .B(G148gat), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n412), .B(new_n411), .C1(new_n416), .C2(KEYINPUT2), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT3), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G127gat), .B(G134gat), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT69), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G113gat), .B(G120gat), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  OR2_X1    g224(.A1(G127gat), .A2(G134gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(G127gat), .A2(G134gat), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(KEYINPUT69), .A3(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n423), .A2(new_n425), .A3(new_n428), .A4(new_n429), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n426), .B(new_n427), .C1(new_n424), .C2(KEYINPUT1), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n420), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n415), .A2(new_n417), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT80), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n415), .A2(new_n417), .A3(KEYINPUT80), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n433), .B1(new_n439), .B2(KEYINPUT3), .ZN(new_n440));
  NAND2_X1  g239(.A1(G225gat), .A2(G233gat), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n442), .A2(KEYINPUT5), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n432), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT83), .ZN(new_n446));
  XNOR2_X1  g245(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n445), .A2(new_n446), .A3(new_n418), .A4(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n430), .A2(new_n417), .A3(new_n415), .A4(new_n431), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT4), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n447), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT83), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n448), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT84), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n450), .B(KEYINPUT83), .C1(new_n449), .C2(new_n452), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT84), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n457), .A3(new_n448), .ZN(new_n458));
  AOI211_X1 g257(.A(new_n440), .B(new_n444), .C1(new_n455), .C2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n449), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n460), .B1(new_n439), .B2(new_n432), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT5), .B1(new_n461), .B2(new_n441), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT82), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n460), .A2(KEYINPUT4), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n442), .B1(new_n449), .B2(new_n447), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n463), .B1(new_n440), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n432), .B(new_n420), .C1(new_n438), .C2(new_n419), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n468), .A2(KEYINPUT82), .A3(new_n464), .A4(new_n465), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n462), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g269(.A(KEYINPUT6), .B(new_n407), .C1(new_n459), .C2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n407), .B1(new_n459), .B2(new_n470), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n454), .A2(KEYINPUT84), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n457), .B1(new_n456), .B2(new_n448), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n468), .B(new_n443), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n467), .A2(new_n469), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n406), .B(new_n475), .C1(new_n476), .C2(new_n462), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n472), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n402), .B1(new_n471), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n393), .A2(new_n395), .A3(KEYINPUT79), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n398), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n445), .B1(new_n331), .B2(new_n345), .ZN(new_n483));
  INV_X1    g282(.A(G227gat), .ZN(new_n484));
  INV_X1    g283(.A(G233gat), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n357), .B(new_n432), .C1(new_n361), .C2(new_n363), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n483), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  XOR2_X1   g287(.A(G15gat), .B(G43gat), .Z(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(KEYINPUT71), .ZN(new_n490));
  XNOR2_X1  g289(.A(G71gat), .B(G99gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT33), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n488), .A2(KEYINPUT32), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT72), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT72), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n488), .A2(new_n496), .A3(KEYINPUT32), .A4(new_n493), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT34), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n487), .ZN(new_n500));
  INV_X1    g299(.A(new_n486), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AOI211_X1 g301(.A(KEYINPUT34), .B(new_n486), .C1(new_n483), .C2(new_n487), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n488), .A2(KEYINPUT32), .ZN(new_n505));
  INV_X1    g304(.A(new_n488), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n505), .B(new_n492), .C1(new_n506), .C2(KEYINPUT33), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n498), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n504), .B1(new_n498), .B2(new_n507), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G78gat), .B(G106gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(G22gat), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G228gat), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n514), .A2(new_n485), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n290), .B1(new_n280), .B2(new_n287), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n438), .B1(new_n516), .B2(new_n419), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n290), .B1(new_n434), .B2(KEYINPUT3), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n278), .A2(new_n279), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n286), .A2(new_n281), .A3(new_n270), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n515), .B1(new_n517), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n515), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT29), .B1(new_n287), .B2(KEYINPUT85), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT85), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n519), .A2(new_n526), .A3(new_n520), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT3), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n524), .B(new_n521), .C1(new_n528), .C2(new_n418), .ZN(new_n529));
  XNOR2_X1  g328(.A(KEYINPUT31), .B(G50gat), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n523), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n531), .B1(new_n523), .B2(new_n529), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n513), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n523), .A2(new_n529), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n530), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n523), .A2(new_n529), .A3(new_n531), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n536), .A2(new_n512), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n510), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT35), .B1(new_n482), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT35), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n534), .A2(new_n538), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n544), .B1(new_n479), .B2(new_n471), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n396), .A2(new_n545), .A3(new_n401), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT73), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n498), .A2(new_n507), .ZN(new_n548));
  INV_X1    g347(.A(new_n504), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n498), .A2(new_n504), .A3(new_n507), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n547), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n548), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT73), .B1(new_n553), .B2(new_n504), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT87), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT73), .B1(new_n508), .B2(new_n509), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT87), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI211_X1 g358(.A(KEYINPUT88), .B(new_n546), .C1(new_n555), .C2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT88), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n555), .A2(new_n559), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n396), .A2(new_n545), .A3(new_n401), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n542), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n396), .A2(new_n401), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n468), .B1(new_n473), .B2(new_n474), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(new_n442), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT39), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n569), .B1(new_n461), .B2(new_n441), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n567), .A2(new_n569), .A3(new_n442), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(new_n406), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT40), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n571), .A2(KEYINPUT40), .A3(new_n406), .A4(new_n572), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n575), .A2(new_n472), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n539), .B1(new_n566), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n367), .A2(new_n378), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n384), .B1(new_n579), .B2(KEYINPUT37), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT37), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n394), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(KEYINPUT38), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n479), .A2(new_n471), .A3(new_n399), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n382), .B1(new_n394), .B2(new_n581), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n386), .A2(new_n372), .A3(new_n387), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n288), .B1(new_n389), .B2(new_n370), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT86), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT86), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n589), .B(new_n288), .C1(new_n389), .C2(new_n370), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(KEYINPUT37), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT38), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n585), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n583), .A2(new_n584), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT36), .B1(new_n556), .B2(new_n558), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n510), .A2(KEYINPUT36), .ZN(new_n597));
  AOI22_X1  g396(.A1(new_n578), .A2(new_n594), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n482), .A2(new_n539), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n266), .B1(new_n565), .B2(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(G190gat), .B(G218gat), .Z(new_n602));
  XNOR2_X1  g401(.A(KEYINPUT103), .B(G85gat), .ZN(new_n603));
  INV_X1    g402(.A(G92gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(G99gat), .A2(G106gat), .ZN(new_n605));
  AOI22_X1  g404(.A1(new_n603), .A2(new_n604), .B1(KEYINPUT8), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT102), .ZN(new_n607));
  INV_X1    g406(.A(G85gat), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n607), .B1(new_n608), .B2(new_n604), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n609), .A2(KEYINPUT7), .ZN(new_n610));
  NAND3_X1  g409(.A1(KEYINPUT102), .A2(G85gat), .A3(G92gat), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n609), .A2(KEYINPUT7), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n606), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G99gat), .B(G106gat), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n606), .A2(new_n610), .A3(new_n614), .A4(new_n612), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n224), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(new_n239), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  AND2_X1   g420(.A1(G232gat), .A2(G233gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT41), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n616), .A2(new_n617), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n623), .B1(new_n247), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n602), .B1(new_n621), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n622), .A2(KEYINPUT41), .ZN(new_n627));
  XNOR2_X1  g426(.A(G134gat), .B(G162gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n625), .ZN(new_n630));
  INV_X1    g429(.A(new_n602), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(new_n620), .A3(new_n631), .ZN(new_n632));
  AND3_X1   g431(.A1(new_n626), .A2(new_n629), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n629), .B1(new_n626), .B2(new_n632), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT98), .ZN(new_n637));
  AOI22_X1  g436(.A1(new_n637), .A2(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(G71gat), .B2(G78gat), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n640));
  AND2_X1   g439(.A1(G57gat), .A2(G64gat), .ZN(new_n641));
  NOR2_X1   g440(.A1(G57gat), .A2(G64gat), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n639), .B(new_n643), .Z(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(KEYINPUT99), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n639), .B(new_n643), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT99), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT100), .B(KEYINPUT21), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g450(.A(G127gat), .B(G155gat), .Z(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT21), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n248), .B1(new_n654), .B2(new_n649), .ZN(new_n655));
  OR2_X1    g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n653), .A2(new_n655), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(G231gat), .A2(G233gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT101), .ZN(new_n660));
  XOR2_X1   g459(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G183gat), .B(G211gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n658), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n656), .A2(new_n657), .A3(new_n664), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(G230gat), .A2(G233gat), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT104), .B(KEYINPUT10), .Z(new_n670));
  NAND2_X1  g469(.A1(new_n618), .A2(new_n646), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n645), .A2(new_n648), .A3(new_n624), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT10), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n649), .A2(new_n674), .A3(new_n624), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n669), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n624), .A2(new_n644), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n646), .B(KEYINPUT99), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n677), .B1(new_n678), .B2(new_n624), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n676), .B1(new_n669), .B2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(G120gat), .B(G148gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(G176gat), .B(G204gat), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n682), .B(new_n683), .Z(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n676), .B(new_n684), .C1(new_n669), .C2(new_n680), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n636), .A2(new_n668), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(KEYINPUT105), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n636), .A2(new_n692), .A3(new_n668), .A4(new_n689), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n601), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n479), .A2(new_n471), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT106), .B(G1gat), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1324gat));
  XNOR2_X1  g498(.A(KEYINPUT16), .B(G8gat), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT42), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n601), .A2(new_n566), .A3(new_n694), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT108), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n402), .B1(new_n393), .B2(new_n395), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n705), .B1(new_n695), .B2(new_n706), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n601), .A2(KEYINPUT107), .A3(new_n566), .A4(new_n694), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(G8gat), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n700), .B1(new_n707), .B2(new_n708), .ZN(new_n710));
  OAI211_X1 g509(.A(new_n704), .B(new_n709), .C1(new_n710), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g510(.A(new_n597), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n595), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(G15gat), .B1(new_n695), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n562), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n716), .A2(G15gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(new_n695), .B2(new_n717), .ZN(G1326gat));
  NOR2_X1   g517(.A1(new_n695), .A2(new_n540), .ZN(new_n719));
  XOR2_X1   g518(.A(KEYINPUT43), .B(G22gat), .Z(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1327gat));
  AND3_X1   g520(.A1(new_n393), .A2(KEYINPUT79), .A3(new_n395), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT79), .B1(new_n393), .B2(new_n395), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n696), .A2(new_n401), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n541), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n543), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n557), .B1(new_n556), .B2(new_n558), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n563), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(KEYINPUT88), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n562), .A2(new_n561), .A3(new_n563), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n727), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n599), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n575), .A2(new_n472), .A3(new_n576), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n540), .B1(new_n706), .B2(new_n735), .ZN(new_n736));
  AND3_X1   g535(.A1(new_n583), .A2(new_n584), .A3(new_n593), .ZN(new_n737));
  OAI22_X1  g536(.A1(new_n736), .A2(new_n737), .B1(new_n595), .B2(new_n712), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  OAI211_X1 g538(.A(KEYINPUT44), .B(new_n635), .C1(new_n733), .C2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n668), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n689), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n742), .B1(new_n261), .B2(new_n262), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n599), .A2(KEYINPUT110), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n482), .A2(new_n745), .A3(new_n539), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n744), .A2(new_n598), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n636), .B1(new_n565), .B2(new_n747), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n740), .B(new_n743), .C1(new_n748), .C2(KEYINPUT44), .ZN(new_n749));
  OAI21_X1  g548(.A(G29gat), .B1(new_n749), .B2(new_n696), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n742), .A2(new_n636), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n601), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n696), .A2(G29gat), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT109), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT109), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n601), .A2(new_n757), .A3(new_n751), .A4(new_n753), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n756), .B1(new_n755), .B2(new_n758), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n750), .B1(new_n759), .B2(new_n760), .ZN(G1328gat));
  NOR3_X1   g560(.A1(new_n752), .A2(G36gat), .A3(new_n706), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT46), .ZN(new_n763));
  OAI21_X1  g562(.A(G36gat), .B1(new_n749), .B2(new_n706), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(G1329gat));
  INV_X1    g564(.A(G43gat), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n752), .B2(new_n716), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n713), .A2(G43gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n749), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(KEYINPUT47), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT47), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n767), .B(new_n771), .C1(new_n749), .C2(new_n768), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(G1330gat));
  INV_X1    g572(.A(G50gat), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(new_n752), .B2(new_n540), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n539), .A2(G50gat), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n775), .B1(new_n749), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT48), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT48), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n775), .B(new_n779), .C1(new_n749), .C2(new_n776), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(G1331gat));
  NAND2_X1  g580(.A1(new_n565), .A2(new_n747), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n261), .A2(new_n262), .ZN(new_n783));
  NOR4_X1   g582(.A1(new_n741), .A2(new_n783), .A3(new_n635), .A4(new_n689), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n696), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g587(.A1(new_n782), .A2(new_n784), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(new_n706), .ZN(new_n790));
  NOR2_X1   g589(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n791));
  AND2_X1   g590(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(new_n790), .B2(new_n791), .ZN(G1333gat));
  INV_X1    g593(.A(G71gat), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n785), .A2(new_n795), .A3(new_n562), .ZN(new_n796));
  OAI21_X1  g595(.A(G71gat), .B1(new_n789), .B2(new_n714), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n798), .B(new_n799), .ZN(G1334gat));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n539), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g601(.A1(new_n783), .A2(new_n668), .ZN(new_n803));
  INV_X1    g602(.A(new_n746), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n745), .B1(new_n482), .B2(new_n539), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n804), .A2(new_n738), .A3(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n635), .B(new_n803), .C1(new_n806), .C2(new_n733), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT51), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n782), .A2(KEYINPUT51), .A3(new_n635), .A4(new_n803), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n809), .A2(KEYINPUT112), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT51), .B1(new_n748), .B2(new_n803), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n696), .A2(new_n689), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n811), .A2(new_n814), .A3(new_n603), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n803), .A2(new_n688), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(KEYINPUT111), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n740), .B(new_n818), .C1(new_n748), .C2(KEYINPUT44), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n819), .A2(new_n696), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n816), .B1(new_n603), .B2(new_n820), .ZN(G1336gat));
  OAI21_X1  g620(.A(G92gat), .B1(new_n819), .B2(new_n706), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n706), .A2(G92gat), .A3(new_n689), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n823), .B1(new_n824), .B2(new_n812), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT52), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n811), .A2(new_n814), .A3(new_n823), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n828), .A2(new_n829), .A3(new_n822), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n827), .A2(new_n830), .ZN(G1337gat));
  NOR3_X1   g630(.A1(new_n716), .A2(G99gat), .A3(new_n689), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(KEYINPUT113), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n811), .A2(new_n814), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(G99gat), .B1(new_n819), .B2(new_n714), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(G1338gat));
  OAI21_X1  g635(.A(G106gat), .B1(new_n819), .B2(new_n540), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n689), .A2(new_n540), .A3(G106gat), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n838), .B1(new_n824), .B2(new_n812), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT53), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n811), .A2(new_n814), .A3(new_n838), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n843), .A3(new_n837), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n841), .A2(new_n844), .ZN(G1339gat));
  NOR2_X1   g644(.A1(new_n690), .A2(new_n783), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT55), .ZN(new_n847));
  INV_X1    g646(.A(new_n669), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n678), .A2(KEYINPUT10), .A3(new_n618), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n848), .B(new_n849), .C1(new_n679), .C2(new_n670), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n850), .A2(new_n676), .A3(KEYINPUT54), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n852), .B(new_n669), .C1(new_n673), .C2(new_n675), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n685), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n847), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n850), .A2(new_n676), .A3(KEYINPUT54), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n856), .A2(KEYINPUT55), .A3(new_n685), .A4(new_n853), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n855), .A2(new_n687), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n250), .A2(new_n251), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n241), .B1(new_n240), .B2(new_n242), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n258), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n262), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n858), .A2(new_n635), .A3(new_n862), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n688), .A2(new_n262), .A3(new_n861), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n864), .B1(new_n783), .B2(new_n858), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n863), .B1(new_n865), .B2(new_n635), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n846), .B1(new_n866), .B2(new_n741), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n867), .A2(new_n696), .A3(new_n566), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n716), .A2(new_n539), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(G113gat), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n870), .A2(new_n871), .A3(new_n266), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n866), .A2(new_n741), .ZN(new_n873));
  INV_X1    g672(.A(new_n846), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n875), .A2(new_n786), .A3(new_n706), .A4(new_n726), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(G113gat), .B1(new_n877), .B2(new_n783), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n872), .A2(new_n878), .ZN(G1340gat));
  OR3_X1    g678(.A1(new_n876), .A2(G120gat), .A3(new_n689), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n868), .A2(new_n688), .A3(new_n869), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT114), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(new_n882), .A3(G120gat), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n882), .B1(new_n881), .B2(G120gat), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n880), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT115), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n886), .B(new_n887), .ZN(G1341gat));
  INV_X1    g687(.A(G127gat), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n870), .A2(new_n889), .A3(new_n741), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n876), .A2(KEYINPUT116), .A3(new_n741), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(G127gat), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT116), .B1(new_n876), .B2(new_n741), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n890), .B1(new_n892), .B2(new_n893), .ZN(G1342gat));
  OR2_X1    g693(.A1(new_n636), .A2(G134gat), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n876), .A2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT56), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n868), .A2(new_n635), .A3(new_n869), .ZN(new_n898));
  AOI22_X1  g697(.A1(new_n896), .A2(new_n897), .B1(new_n898), .B2(G134gat), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT117), .ZN(new_n900));
  INV_X1    g699(.A(new_n896), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(KEYINPUT56), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n900), .B(KEYINPUT56), .C1(new_n876), .C2(new_n895), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n899), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT118), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT118), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n907), .B(new_n899), .C1(new_n902), .C2(new_n904), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(G1343gat));
  NAND4_X1  g708(.A1(new_n875), .A2(new_n786), .A3(new_n539), .A4(new_n714), .ZN(new_n910));
  INV_X1    g709(.A(new_n266), .ZN(new_n911));
  INV_X1    g710(.A(G141gat), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n910), .A2(new_n566), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n867), .A2(new_n540), .ZN(new_n915));
  XOR2_X1   g714(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT57), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n540), .A2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n922), .B1(new_n851), .B2(new_n854), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n856), .A2(KEYINPUT120), .A3(new_n685), .A4(new_n853), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n923), .A2(new_n847), .A3(new_n924), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n857), .A2(new_n687), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n927), .B1(new_n264), .B2(new_n265), .ZN(new_n928));
  INV_X1    g727(.A(new_n864), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n635), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n863), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n741), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n921), .B1(new_n932), .B2(new_n874), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n918), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n713), .A2(new_n566), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n786), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n783), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n914), .B1(new_n938), .B2(G141gat), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT58), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT121), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n910), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n566), .B1(new_n910), .B2(new_n941), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n940), .B1(new_n944), .B2(new_n913), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n912), .B1(new_n937), .B2(new_n911), .ZN(new_n946));
  OAI22_X1  g745(.A1(new_n939), .A2(new_n940), .B1(new_n945), .B2(new_n946), .ZN(G1344gat));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n867), .A2(new_n540), .A3(new_n916), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n925), .A2(new_n926), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT97), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n783), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n950), .B1(new_n952), .B2(new_n263), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n636), .B1(new_n953), .B2(new_n864), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n668), .B1(new_n954), .B2(new_n863), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n691), .A2(new_n266), .A3(new_n693), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n539), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n949), .B1(new_n957), .B2(new_n919), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n935), .A2(new_n815), .ZN(new_n959));
  OAI21_X1  g758(.A(G148gat), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(new_n936), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n688), .B(new_n961), .C1(new_n918), .C2(new_n933), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT59), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n963), .A2(G148gat), .ZN(new_n964));
  AOI22_X1  g763(.A1(new_n960), .A2(KEYINPUT59), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n944), .A2(G148gat), .A3(new_n689), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n948), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n942), .A2(new_n943), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n689), .A2(G148gat), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n915), .A2(new_n917), .ZN(new_n971));
  INV_X1    g770(.A(new_n956), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n540), .B1(new_n932), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n971), .B1(new_n973), .B2(KEYINPUT57), .ZN(new_n974));
  INV_X1    g773(.A(new_n959), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n963), .B1(new_n976), .B2(G148gat), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n962), .A2(new_n964), .ZN(new_n978));
  OAI211_X1 g777(.A(new_n970), .B(KEYINPUT122), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n967), .A2(new_n979), .ZN(G1345gat));
  NOR2_X1   g779(.A1(new_n944), .A2(new_n741), .ZN(new_n981));
  AOI21_X1  g780(.A(G155gat), .B1(new_n981), .B2(KEYINPUT123), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT123), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n983), .B1(new_n944), .B2(new_n741), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n741), .A2(new_n409), .ZN(new_n985));
  AOI22_X1  g784(.A1(new_n982), .A2(new_n984), .B1(new_n937), .B2(new_n985), .ZN(G1346gat));
  AOI21_X1  g785(.A(G162gat), .B1(new_n968), .B2(new_n635), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n636), .A2(new_n410), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n987), .B1(new_n937), .B2(new_n988), .ZN(G1347gat));
  NOR3_X1   g788(.A1(new_n867), .A2(new_n786), .A3(new_n706), .ZN(new_n990));
  AND2_X1   g789(.A1(new_n990), .A2(new_n869), .ZN(new_n991));
  INV_X1    g790(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g791(.A(G169gat), .B1(new_n992), .B2(new_n266), .ZN(new_n993));
  AND2_X1   g792(.A1(new_n990), .A2(new_n726), .ZN(new_n994));
  NAND4_X1  g793(.A1(new_n994), .A2(new_n310), .A3(new_n312), .A4(new_n783), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n993), .A2(new_n995), .ZN(G1348gat));
  OAI21_X1  g795(.A(G176gat), .B1(new_n992), .B2(new_n689), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n994), .A2(new_n297), .A3(new_n688), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(new_n998), .ZN(G1349gat));
  NAND2_X1  g798(.A1(new_n991), .A2(new_n668), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n1000), .A2(G183gat), .ZN(new_n1001));
  NAND4_X1  g800(.A1(new_n994), .A2(new_n337), .A3(new_n339), .A4(new_n668), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n1001), .A2(KEYINPUT124), .A3(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g802(.A(new_n1003), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g803(.A1(new_n994), .A2(new_n315), .A3(new_n635), .ZN(new_n1005));
  OAI21_X1  g804(.A(G190gat), .B1(new_n992), .B2(new_n636), .ZN(new_n1006));
  AND2_X1   g805(.A1(new_n1006), .A2(KEYINPUT61), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n1006), .A2(KEYINPUT61), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1005), .B1(new_n1007), .B2(new_n1008), .ZN(G1351gat));
  NOR3_X1   g808(.A1(new_n713), .A2(new_n786), .A3(new_n706), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n915), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g810(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g811(.A(G197gat), .B1(new_n1012), .B2(new_n783), .ZN(new_n1013));
  AND2_X1   g812(.A1(new_n974), .A2(new_n1010), .ZN(new_n1014));
  NOR2_X1   g813(.A1(new_n266), .A2(new_n273), .ZN(new_n1015));
  AOI21_X1  g814(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(G1352gat));
  XOR2_X1   g815(.A(KEYINPUT125), .B(G204gat), .Z(new_n1017));
  NOR3_X1   g816(.A1(new_n1011), .A2(new_n689), .A3(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g817(.A(new_n1018), .B(KEYINPUT62), .ZN(new_n1019));
  NAND3_X1  g818(.A1(new_n1014), .A2(KEYINPUT126), .A3(new_n688), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1020), .A2(new_n1017), .ZN(new_n1021));
  AOI21_X1  g820(.A(KEYINPUT126), .B1(new_n1014), .B2(new_n688), .ZN(new_n1022));
  OAI21_X1  g821(.A(new_n1019), .B1(new_n1021), .B2(new_n1022), .ZN(G1353gat));
  NAND3_X1  g822(.A1(new_n1012), .A2(new_n268), .A3(new_n668), .ZN(new_n1024));
  NAND3_X1  g823(.A1(new_n974), .A2(new_n668), .A3(new_n1010), .ZN(new_n1025));
  AND3_X1   g824(.A1(new_n1025), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1026));
  AOI21_X1  g825(.A(KEYINPUT63), .B1(new_n1025), .B2(G211gat), .ZN(new_n1027));
  OAI21_X1  g826(.A(new_n1024), .B1(new_n1026), .B2(new_n1027), .ZN(G1354gat));
  OAI21_X1  g827(.A(new_n635), .B1(new_n1014), .B2(KEYINPUT127), .ZN(new_n1029));
  AND3_X1   g828(.A1(new_n974), .A2(KEYINPUT127), .A3(new_n1010), .ZN(new_n1030));
  OAI21_X1  g829(.A(G218gat), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g830(.A1(new_n1012), .A2(new_n269), .A3(new_n635), .ZN(new_n1032));
  NAND2_X1  g831(.A1(new_n1031), .A2(new_n1032), .ZN(G1355gat));
endmodule


