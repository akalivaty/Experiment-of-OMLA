

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U554 ( .A1(n690), .A2(n802), .ZN(n733) );
  XOR2_X1 U555 ( .A(KEYINPUT14), .B(n561), .Z(n520) );
  INV_X1 U556 ( .A(KEYINPUT29), .ZN(n717) );
  XNOR2_X1 U557 ( .A(n562), .B(KEYINPUT72), .ZN(n563) );
  NOR2_X1 U558 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U559 ( .A(n564), .B(n563), .ZN(n566) );
  XNOR2_X1 U560 ( .A(KEYINPUT102), .B(n762), .ZN(n763) );
  INV_X1 U561 ( .A(G651), .ZN(n525) );
  NOR2_X1 U562 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U563 ( .A1(G651), .A2(G543), .ZN(n641) );
  XNOR2_X1 U564 ( .A(KEYINPUT1), .B(n527), .ZN(n645) );
  AND2_X1 U565 ( .A1(n827), .A2(n826), .ZN(n828) );
  XOR2_X1 U566 ( .A(KEYINPUT64), .B(n543), .Z(G160) );
  NAND2_X1 U567 ( .A1(n641), .A2(G89), .ZN(n521) );
  XNOR2_X1 U568 ( .A(n521), .B(KEYINPUT4), .ZN(n523) );
  XOR2_X1 U569 ( .A(KEYINPUT0), .B(G543), .Z(n623) );
  NOR2_X1 U570 ( .A1(n623), .A2(n525), .ZN(n638) );
  NAND2_X1 U571 ( .A1(G76), .A2(n638), .ZN(n522) );
  NAND2_X1 U572 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U573 ( .A(n524), .B(KEYINPUT5), .ZN(n532) );
  NOR2_X2 U574 ( .A1(G651), .A2(n623), .ZN(n642) );
  NAND2_X1 U575 ( .A1(n642), .A2(G51), .ZN(n529) );
  NOR2_X1 U576 ( .A1(G543), .A2(n525), .ZN(n526) );
  XOR2_X1 U577 ( .A(KEYINPUT66), .B(n526), .Z(n527) );
  NAND2_X1 U578 ( .A1(G63), .A2(n645), .ZN(n528) );
  NAND2_X1 U579 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U580 ( .A(KEYINPUT6), .B(n530), .Z(n531) );
  NAND2_X1 U581 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U582 ( .A(n533), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U583 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U584 ( .A(G2105), .ZN(n537) );
  NOR2_X1 U585 ( .A1(G2104), .A2(n537), .ZN(n883) );
  NAND2_X1 U586 ( .A1(n883), .A2(G125), .ZN(n542) );
  AND2_X1 U587 ( .A1(G2104), .A2(G2105), .ZN(n882) );
  NAND2_X1 U588 ( .A1(G113), .A2(n882), .ZN(n536) );
  NOR2_X1 U589 ( .A1(G2104), .A2(G2105), .ZN(n534) );
  XOR2_X2 U590 ( .A(KEYINPUT17), .B(n534), .Z(n887) );
  NAND2_X1 U591 ( .A1(G137), .A2(n887), .ZN(n535) );
  NAND2_X1 U592 ( .A1(n536), .A2(n535), .ZN(n540) );
  AND2_X1 U593 ( .A1(n537), .A2(G2104), .ZN(n886) );
  NAND2_X1 U594 ( .A1(G101), .A2(n886), .ZN(n538) );
  XNOR2_X1 U595 ( .A(KEYINPUT23), .B(n538), .ZN(n539) );
  NOR2_X1 U596 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U597 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U598 ( .A1(n642), .A2(G52), .ZN(n545) );
  NAND2_X1 U599 ( .A1(G64), .A2(n645), .ZN(n544) );
  NAND2_X1 U600 ( .A1(n545), .A2(n544), .ZN(n551) );
  NAND2_X1 U601 ( .A1(G90), .A2(n641), .ZN(n547) );
  NAND2_X1 U602 ( .A1(G77), .A2(n638), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U604 ( .A(KEYINPUT9), .B(n548), .Z(n549) );
  XNOR2_X1 U605 ( .A(KEYINPUT68), .B(n549), .ZN(n550) );
  NOR2_X1 U606 ( .A1(n551), .A2(n550), .ZN(G171) );
  AND2_X1 U607 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U608 ( .A(G132), .ZN(G219) );
  INV_X1 U609 ( .A(G82), .ZN(G220) );
  NAND2_X1 U610 ( .A1(G88), .A2(n641), .ZN(n553) );
  NAND2_X1 U611 ( .A1(G75), .A2(n638), .ZN(n552) );
  NAND2_X1 U612 ( .A1(n553), .A2(n552), .ZN(n557) );
  NAND2_X1 U613 ( .A1(n642), .A2(G50), .ZN(n555) );
  NAND2_X1 U614 ( .A1(G62), .A2(n645), .ZN(n554) );
  NAND2_X1 U615 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U616 ( .A1(n557), .A2(n556), .ZN(G166) );
  NAND2_X1 U617 ( .A1(G7), .A2(G661), .ZN(n558) );
  XNOR2_X1 U618 ( .A(n558), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U619 ( .A(G223), .ZN(n829) );
  NAND2_X1 U620 ( .A1(n829), .A2(G567), .ZN(n559) );
  XNOR2_X1 U621 ( .A(n559), .B(KEYINPUT11), .ZN(n560) );
  XNOR2_X1 U622 ( .A(KEYINPUT71), .B(n560), .ZN(G234) );
  NAND2_X1 U623 ( .A1(G56), .A2(n645), .ZN(n561) );
  NAND2_X1 U624 ( .A1(G81), .A2(n641), .ZN(n564) );
  XOR2_X1 U625 ( .A(KEYINPUT12), .B(KEYINPUT73), .Z(n562) );
  NAND2_X1 U626 ( .A1(n638), .A2(G68), .ZN(n565) );
  NAND2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U628 ( .A(KEYINPUT13), .B(n567), .Z(n568) );
  NOR2_X1 U629 ( .A1(n520), .A2(n568), .ZN(n569) );
  XNOR2_X1 U630 ( .A(KEYINPUT74), .B(n569), .ZN(n571) );
  NAND2_X1 U631 ( .A1(G43), .A2(n642), .ZN(n570) );
  NAND2_X1 U632 ( .A1(n571), .A2(n570), .ZN(n599) );
  INV_X2 U633 ( .A(n599), .ZN(n694) );
  NAND2_X1 U634 ( .A1(n694), .A2(G860), .ZN(G153) );
  INV_X1 U635 ( .A(G171), .ZN(G301) );
  NAND2_X1 U636 ( .A1(G868), .A2(G301), .ZN(n583) );
  NAND2_X1 U637 ( .A1(n641), .A2(G92), .ZN(n573) );
  NAND2_X1 U638 ( .A1(G66), .A2(n645), .ZN(n572) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n580) );
  NAND2_X1 U640 ( .A1(n638), .A2(G79), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n574), .B(KEYINPUT75), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n642), .A2(G54), .ZN(n575) );
  XOR2_X1 U643 ( .A(KEYINPUT76), .B(n575), .Z(n576) );
  NOR2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n578), .B(KEYINPUT77), .ZN(n579) );
  XOR2_X1 U646 ( .A(KEYINPUT15), .B(n581), .Z(n941) );
  OR2_X1 U647 ( .A1(n941), .A2(G868), .ZN(n582) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(G284) );
  NAND2_X1 U649 ( .A1(n642), .A2(G53), .ZN(n585) );
  NAND2_X1 U650 ( .A1(G65), .A2(n645), .ZN(n584) );
  NAND2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n589) );
  NAND2_X1 U652 ( .A1(G91), .A2(n641), .ZN(n587) );
  NAND2_X1 U653 ( .A1(G78), .A2(n638), .ZN(n586) );
  NAND2_X1 U654 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U655 ( .A1(n589), .A2(n588), .ZN(n922) );
  XNOR2_X1 U656 ( .A(n922), .B(KEYINPUT69), .ZN(G299) );
  NOR2_X1 U657 ( .A1(G868), .A2(G299), .ZN(n590) );
  XNOR2_X1 U658 ( .A(n590), .B(KEYINPUT78), .ZN(n592) );
  INV_X1 U659 ( .A(G868), .ZN(n661) );
  NOR2_X1 U660 ( .A1(n661), .A2(G286), .ZN(n591) );
  NOR2_X1 U661 ( .A1(n592), .A2(n591), .ZN(G297) );
  INV_X1 U662 ( .A(G860), .ZN(n593) );
  NAND2_X1 U663 ( .A1(n593), .A2(G559), .ZN(n594) );
  NAND2_X1 U664 ( .A1(n594), .A2(n941), .ZN(n595) );
  XNOR2_X1 U665 ( .A(n595), .B(KEYINPUT16), .ZN(n596) );
  XOR2_X1 U666 ( .A(KEYINPUT79), .B(n596), .Z(G148) );
  NAND2_X1 U667 ( .A1(n941), .A2(G868), .ZN(n597) );
  NOR2_X1 U668 ( .A1(G559), .A2(n597), .ZN(n598) );
  XNOR2_X1 U669 ( .A(n598), .B(KEYINPUT80), .ZN(n601) );
  NOR2_X1 U670 ( .A1(n599), .A2(G868), .ZN(n600) );
  NOR2_X1 U671 ( .A1(n601), .A2(n600), .ZN(G282) );
  NAND2_X1 U672 ( .A1(G111), .A2(n882), .ZN(n603) );
  NAND2_X1 U673 ( .A1(G99), .A2(n886), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U675 ( .A(n604), .B(KEYINPUT81), .ZN(n606) );
  NAND2_X1 U676 ( .A1(G135), .A2(n887), .ZN(n605) );
  NAND2_X1 U677 ( .A1(n606), .A2(n605), .ZN(n609) );
  NAND2_X1 U678 ( .A1(n883), .A2(G123), .ZN(n607) );
  XOR2_X1 U679 ( .A(KEYINPUT18), .B(n607), .Z(n608) );
  NOR2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n996) );
  XNOR2_X1 U681 ( .A(n996), .B(G2096), .ZN(n611) );
  INV_X1 U682 ( .A(G2100), .ZN(n610) );
  NAND2_X1 U683 ( .A1(n611), .A2(n610), .ZN(G156) );
  NAND2_X1 U684 ( .A1(n642), .A2(G55), .ZN(n613) );
  NAND2_X1 U685 ( .A1(G67), .A2(n645), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n614) );
  XOR2_X1 U687 ( .A(KEYINPUT84), .B(n614), .Z(n616) );
  NAND2_X1 U688 ( .A1(n641), .A2(G93), .ZN(n615) );
  NAND2_X1 U689 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U690 ( .A1(G80), .A2(n638), .ZN(n617) );
  XNOR2_X1 U691 ( .A(KEYINPUT83), .B(n617), .ZN(n618) );
  OR2_X1 U692 ( .A1(n619), .A2(n618), .ZN(n662) );
  NAND2_X1 U693 ( .A1(n941), .A2(G559), .ZN(n658) );
  XOR2_X1 U694 ( .A(n694), .B(KEYINPUT82), .Z(n620) );
  XNOR2_X1 U695 ( .A(n658), .B(n620), .ZN(n621) );
  NOR2_X1 U696 ( .A1(G860), .A2(n621), .ZN(n622) );
  XOR2_X1 U697 ( .A(n662), .B(n622), .Z(G145) );
  NAND2_X1 U698 ( .A1(G87), .A2(n623), .ZN(n625) );
  NAND2_X1 U699 ( .A1(G74), .A2(G651), .ZN(n624) );
  NAND2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U701 ( .A1(n645), .A2(n626), .ZN(n629) );
  NAND2_X1 U702 ( .A1(G49), .A2(n642), .ZN(n627) );
  XOR2_X1 U703 ( .A(KEYINPUT85), .B(n627), .Z(n628) );
  NAND2_X1 U704 ( .A1(n629), .A2(n628), .ZN(G288) );
  NAND2_X1 U705 ( .A1(n638), .A2(G72), .ZN(n632) );
  NAND2_X1 U706 ( .A1(G60), .A2(n645), .ZN(n630) );
  XOR2_X1 U707 ( .A(KEYINPUT67), .B(n630), .Z(n631) );
  NAND2_X1 U708 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U709 ( .A1(G85), .A2(n641), .ZN(n633) );
  XNOR2_X1 U710 ( .A(KEYINPUT65), .B(n633), .ZN(n634) );
  NOR2_X1 U711 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U712 ( .A1(n642), .A2(G47), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n637), .A2(n636), .ZN(G290) );
  XOR2_X1 U714 ( .A(KEYINPUT87), .B(KEYINPUT2), .Z(n640) );
  NAND2_X1 U715 ( .A1(G73), .A2(n638), .ZN(n639) );
  XNOR2_X1 U716 ( .A(n640), .B(n639), .ZN(n650) );
  NAND2_X1 U717 ( .A1(G86), .A2(n641), .ZN(n644) );
  NAND2_X1 U718 ( .A1(G48), .A2(n642), .ZN(n643) );
  NAND2_X1 U719 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U720 ( .A1(n645), .A2(G61), .ZN(n646) );
  XOR2_X1 U721 ( .A(KEYINPUT86), .B(n646), .Z(n647) );
  NOR2_X1 U722 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U723 ( .A1(n650), .A2(n649), .ZN(G305) );
  XNOR2_X1 U724 ( .A(KEYINPUT88), .B(KEYINPUT19), .ZN(n652) );
  XOR2_X1 U725 ( .A(G288), .B(n662), .Z(n651) );
  XNOR2_X1 U726 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U727 ( .A(G166), .B(n653), .ZN(n655) );
  XNOR2_X1 U728 ( .A(G290), .B(n694), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U730 ( .A(n656), .B(G305), .ZN(n657) );
  XNOR2_X1 U731 ( .A(n657), .B(G299), .ZN(n900) );
  XNOR2_X1 U732 ( .A(n900), .B(n658), .ZN(n659) );
  NAND2_X1 U733 ( .A1(n659), .A2(G868), .ZN(n660) );
  XOR2_X1 U734 ( .A(KEYINPUT89), .B(n660), .Z(n664) );
  NAND2_X1 U735 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U736 ( .A1(n664), .A2(n663), .ZN(G295) );
  NAND2_X1 U737 ( .A1(G2078), .A2(G2084), .ZN(n666) );
  XOR2_X1 U738 ( .A(KEYINPUT90), .B(KEYINPUT20), .Z(n665) );
  XNOR2_X1 U739 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U740 ( .A1(G2090), .A2(n667), .ZN(n668) );
  XNOR2_X1 U741 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U742 ( .A1(n669), .A2(G2072), .ZN(G158) );
  XOR2_X1 U743 ( .A(KEYINPUT70), .B(G57), .Z(G237) );
  XNOR2_X1 U744 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U745 ( .A1(G108), .A2(G120), .ZN(n670) );
  NOR2_X1 U746 ( .A1(G237), .A2(n670), .ZN(n671) );
  NAND2_X1 U747 ( .A1(G69), .A2(n671), .ZN(n836) );
  NAND2_X1 U748 ( .A1(n836), .A2(G567), .ZN(n676) );
  NOR2_X1 U749 ( .A1(G220), .A2(G219), .ZN(n672) );
  XOR2_X1 U750 ( .A(KEYINPUT22), .B(n672), .Z(n673) );
  NOR2_X1 U751 ( .A1(G218), .A2(n673), .ZN(n674) );
  NAND2_X1 U752 ( .A1(G96), .A2(n674), .ZN(n837) );
  NAND2_X1 U753 ( .A1(n837), .A2(G2106), .ZN(n675) );
  NAND2_X1 U754 ( .A1(n676), .A2(n675), .ZN(n856) );
  NAND2_X1 U755 ( .A1(G483), .A2(G661), .ZN(n677) );
  NOR2_X1 U756 ( .A1(n856), .A2(n677), .ZN(n834) );
  NAND2_X1 U757 ( .A1(n834), .A2(G36), .ZN(n678) );
  XOR2_X1 U758 ( .A(KEYINPUT91), .B(n678), .Z(G176) );
  NAND2_X1 U759 ( .A1(n882), .A2(G114), .ZN(n679) );
  XNOR2_X1 U760 ( .A(n679), .B(KEYINPUT92), .ZN(n681) );
  NAND2_X1 U761 ( .A1(G102), .A2(n886), .ZN(n680) );
  NAND2_X1 U762 ( .A1(n681), .A2(n680), .ZN(n685) );
  NAND2_X1 U763 ( .A1(G138), .A2(n887), .ZN(n683) );
  NAND2_X1 U764 ( .A1(G126), .A2(n883), .ZN(n682) );
  NAND2_X1 U765 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U766 ( .A1(n685), .A2(n684), .ZN(G164) );
  INV_X1 U767 ( .A(G166), .ZN(G303) );
  NAND2_X1 U768 ( .A1(G40), .A2(G160), .ZN(n801) );
  INV_X1 U769 ( .A(n801), .ZN(n690) );
  NOR2_X1 U770 ( .A1(G164), .A2(G1384), .ZN(n802) );
  NAND2_X1 U771 ( .A1(G8), .A2(n733), .ZN(n770) );
  NOR2_X1 U772 ( .A1(G1981), .A2(G305), .ZN(n686) );
  XOR2_X1 U773 ( .A(n686), .B(KEYINPUT24), .Z(n687) );
  NOR2_X1 U774 ( .A1(n770), .A2(n687), .ZN(n765) );
  XOR2_X1 U775 ( .A(G1981), .B(G305), .Z(n937) );
  AND2_X1 U776 ( .A1(G1341), .A2(KEYINPUT26), .ZN(n688) );
  NAND2_X1 U777 ( .A1(n733), .A2(n688), .ZN(n696) );
  AND2_X1 U778 ( .A1(n802), .A2(G1996), .ZN(n689) );
  NAND2_X1 U779 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U780 ( .A(n691), .B(KEYINPUT26), .ZN(n692) );
  NAND2_X1 U781 ( .A1(n696), .A2(n692), .ZN(n693) );
  NAND2_X1 U782 ( .A1(KEYINPUT100), .A2(n693), .ZN(n695) );
  NAND2_X1 U783 ( .A1(n695), .A2(n694), .ZN(n699) );
  INV_X1 U784 ( .A(n696), .ZN(n697) );
  NOR2_X1 U785 ( .A1(n697), .A2(KEYINPUT100), .ZN(n698) );
  NOR2_X2 U786 ( .A1(n699), .A2(n698), .ZN(n701) );
  NOR2_X1 U787 ( .A1(n701), .A2(n941), .ZN(n700) );
  XNOR2_X1 U788 ( .A(n700), .B(KEYINPUT101), .ZN(n707) );
  NAND2_X1 U789 ( .A1(n701), .A2(n941), .ZN(n705) );
  INV_X2 U790 ( .A(n733), .ZN(n719) );
  NOR2_X1 U791 ( .A1(n719), .A2(G1348), .ZN(n703) );
  NOR2_X1 U792 ( .A1(G2067), .A2(n733), .ZN(n702) );
  NOR2_X1 U793 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U794 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U795 ( .A1(n707), .A2(n706), .ZN(n712) );
  NAND2_X1 U796 ( .A1(n719), .A2(G2072), .ZN(n708) );
  XNOR2_X1 U797 ( .A(n708), .B(KEYINPUT27), .ZN(n710) );
  INV_X1 U798 ( .A(G1956), .ZN(n948) );
  NOR2_X1 U799 ( .A1(n948), .A2(n719), .ZN(n709) );
  NOR2_X1 U800 ( .A1(n710), .A2(n709), .ZN(n713) );
  NAND2_X1 U801 ( .A1(n922), .A2(n713), .ZN(n711) );
  NAND2_X1 U802 ( .A1(n712), .A2(n711), .ZN(n716) );
  NOR2_X1 U803 ( .A1(n922), .A2(n713), .ZN(n714) );
  XOR2_X1 U804 ( .A(n714), .B(KEYINPUT28), .Z(n715) );
  NAND2_X1 U805 ( .A1(n716), .A2(n715), .ZN(n718) );
  XNOR2_X1 U806 ( .A(n718), .B(n717), .ZN(n723) );
  OR2_X1 U807 ( .A1(n719), .A2(G1961), .ZN(n721) );
  XNOR2_X1 U808 ( .A(G2078), .B(KEYINPUT25), .ZN(n977) );
  NAND2_X1 U809 ( .A1(n719), .A2(n977), .ZN(n720) );
  NAND2_X1 U810 ( .A1(n721), .A2(n720), .ZN(n727) );
  NAND2_X1 U811 ( .A1(n727), .A2(G171), .ZN(n722) );
  NAND2_X1 U812 ( .A1(n723), .A2(n722), .ZN(n732) );
  NOR2_X1 U813 ( .A1(G1966), .A2(n770), .ZN(n745) );
  NOR2_X1 U814 ( .A1(G2084), .A2(n733), .ZN(n741) );
  NOR2_X1 U815 ( .A1(n745), .A2(n741), .ZN(n724) );
  NAND2_X1 U816 ( .A1(G8), .A2(n724), .ZN(n725) );
  XNOR2_X1 U817 ( .A(KEYINPUT30), .B(n725), .ZN(n726) );
  NOR2_X1 U818 ( .A1(G168), .A2(n726), .ZN(n729) );
  NOR2_X1 U819 ( .A1(G171), .A2(n727), .ZN(n728) );
  NOR2_X1 U820 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U821 ( .A(KEYINPUT31), .B(n730), .Z(n731) );
  NAND2_X1 U822 ( .A1(n732), .A2(n731), .ZN(n743) );
  NAND2_X1 U823 ( .A1(n743), .A2(G286), .ZN(n738) );
  NOR2_X1 U824 ( .A1(G1971), .A2(n770), .ZN(n735) );
  NOR2_X1 U825 ( .A1(G2090), .A2(n733), .ZN(n734) );
  NOR2_X1 U826 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U827 ( .A1(n736), .A2(G303), .ZN(n737) );
  NAND2_X1 U828 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U829 ( .A1(n739), .A2(G8), .ZN(n740) );
  XNOR2_X1 U830 ( .A(n740), .B(KEYINPUT32), .ZN(n749) );
  NAND2_X1 U831 ( .A1(G8), .A2(n741), .ZN(n742) );
  XOR2_X1 U832 ( .A(KEYINPUT99), .B(n742), .Z(n747) );
  INV_X1 U833 ( .A(n743), .ZN(n744) );
  NOR2_X1 U834 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U835 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U836 ( .A1(n749), .A2(n748), .ZN(n768) );
  NOR2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n928) );
  NOR2_X1 U838 ( .A1(G1971), .A2(G303), .ZN(n750) );
  NOR2_X1 U839 ( .A1(n928), .A2(n750), .ZN(n752) );
  INV_X1 U840 ( .A(KEYINPUT33), .ZN(n751) );
  AND2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U842 ( .A1(n768), .A2(n753), .ZN(n757) );
  INV_X1 U843 ( .A(n770), .ZN(n754) );
  NAND2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n923) );
  AND2_X1 U845 ( .A1(n754), .A2(n923), .ZN(n755) );
  OR2_X1 U846 ( .A1(KEYINPUT33), .A2(n755), .ZN(n756) );
  NAND2_X1 U847 ( .A1(n757), .A2(n756), .ZN(n760) );
  NAND2_X1 U848 ( .A1(n928), .A2(KEYINPUT33), .ZN(n758) );
  NOR2_X1 U849 ( .A1(n758), .A2(n770), .ZN(n759) );
  NAND2_X1 U850 ( .A1(n937), .A2(n761), .ZN(n762) );
  INV_X1 U851 ( .A(n763), .ZN(n764) );
  NOR2_X1 U852 ( .A1(n765), .A2(n764), .ZN(n816) );
  NAND2_X1 U853 ( .A1(G8), .A2(G166), .ZN(n766) );
  NOR2_X1 U854 ( .A1(G2090), .A2(n766), .ZN(n767) );
  XNOR2_X1 U855 ( .A(n767), .B(KEYINPUT103), .ZN(n769) );
  NAND2_X1 U856 ( .A1(n769), .A2(n768), .ZN(n771) );
  NAND2_X1 U857 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U858 ( .A(n772), .B(KEYINPUT104), .ZN(n814) );
  XNOR2_X1 U859 ( .A(KEYINPUT37), .B(G2067), .ZN(n809) );
  NAND2_X1 U860 ( .A1(n886), .A2(G104), .ZN(n773) );
  XNOR2_X1 U861 ( .A(n773), .B(KEYINPUT94), .ZN(n775) );
  NAND2_X1 U862 ( .A1(G140), .A2(n887), .ZN(n774) );
  NAND2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U864 ( .A(KEYINPUT34), .B(n776), .ZN(n783) );
  NAND2_X1 U865 ( .A1(n883), .A2(G128), .ZN(n777) );
  XNOR2_X1 U866 ( .A(KEYINPUT95), .B(n777), .ZN(n780) );
  NAND2_X1 U867 ( .A1(n882), .A2(G116), .ZN(n778) );
  XOR2_X1 U868 ( .A(KEYINPUT96), .B(n778), .Z(n779) );
  NOR2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U870 ( .A(n781), .B(KEYINPUT35), .ZN(n782) );
  NOR2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U872 ( .A(KEYINPUT36), .B(n784), .ZN(n879) );
  NAND2_X1 U873 ( .A1(n809), .A2(n879), .ZN(n1014) );
  NAND2_X1 U874 ( .A1(G117), .A2(n882), .ZN(n786) );
  NAND2_X1 U875 ( .A1(G141), .A2(n887), .ZN(n785) );
  NAND2_X1 U876 ( .A1(n786), .A2(n785), .ZN(n789) );
  NAND2_X1 U877 ( .A1(n886), .A2(G105), .ZN(n787) );
  XOR2_X1 U878 ( .A(KEYINPUT38), .B(n787), .Z(n788) );
  NOR2_X1 U879 ( .A1(n789), .A2(n788), .ZN(n791) );
  NAND2_X1 U880 ( .A1(n883), .A2(G129), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n791), .A2(n790), .ZN(n893) );
  NOR2_X1 U882 ( .A1(n893), .A2(G1996), .ZN(n792) );
  XNOR2_X1 U883 ( .A(n792), .B(KEYINPUT105), .ZN(n1008) );
  NAND2_X1 U884 ( .A1(G107), .A2(n882), .ZN(n794) );
  NAND2_X1 U885 ( .A1(G95), .A2(n886), .ZN(n793) );
  NAND2_X1 U886 ( .A1(n794), .A2(n793), .ZN(n798) );
  NAND2_X1 U887 ( .A1(G131), .A2(n887), .ZN(n796) );
  NAND2_X1 U888 ( .A1(G119), .A2(n883), .ZN(n795) );
  NAND2_X1 U889 ( .A1(n796), .A2(n795), .ZN(n797) );
  OR2_X1 U890 ( .A1(n798), .A2(n797), .ZN(n865) );
  NOR2_X1 U891 ( .A1(G1991), .A2(n865), .ZN(n997) );
  NOR2_X1 U892 ( .A1(G1986), .A2(G290), .ZN(n799) );
  NOR2_X1 U893 ( .A1(n997), .A2(n799), .ZN(n800) );
  XOR2_X1 U894 ( .A(KEYINPUT106), .B(n800), .Z(n806) );
  NOR2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n821) );
  XNOR2_X1 U896 ( .A(KEYINPUT98), .B(n821), .ZN(n805) );
  NAND2_X1 U897 ( .A1(G1996), .A2(n893), .ZN(n804) );
  NAND2_X1 U898 ( .A1(G1991), .A2(n865), .ZN(n803) );
  NAND2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n1005) );
  NAND2_X1 U900 ( .A1(n805), .A2(n1005), .ZN(n819) );
  NAND2_X1 U901 ( .A1(n806), .A2(n819), .ZN(n807) );
  NAND2_X1 U902 ( .A1(n1008), .A2(n807), .ZN(n808) );
  XOR2_X1 U903 ( .A(KEYINPUT39), .B(n808), .Z(n811) );
  NOR2_X1 U904 ( .A1(n809), .A2(n879), .ZN(n1017) );
  NAND2_X1 U905 ( .A1(n821), .A2(n1017), .ZN(n810) );
  XOR2_X1 U906 ( .A(KEYINPUT97), .B(n810), .Z(n818) );
  NAND2_X1 U907 ( .A1(n811), .A2(n818), .ZN(n812) );
  NAND2_X1 U908 ( .A1(n1014), .A2(n812), .ZN(n813) );
  NAND2_X1 U909 ( .A1(n813), .A2(n821), .ZN(n817) );
  AND2_X1 U910 ( .A1(n814), .A2(n817), .ZN(n815) );
  NAND2_X1 U911 ( .A1(n816), .A2(n815), .ZN(n827) );
  INV_X1 U912 ( .A(n817), .ZN(n825) );
  NAND2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n823) );
  XOR2_X1 U914 ( .A(G1986), .B(KEYINPUT93), .Z(n820) );
  XNOR2_X1 U915 ( .A(G290), .B(n820), .ZN(n932) );
  AND2_X1 U916 ( .A1(n932), .A2(n821), .ZN(n822) );
  NOR2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n824) );
  OR2_X1 U918 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U919 ( .A(n828), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n829), .ZN(G217) );
  NAND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n831) );
  INV_X1 U922 ( .A(G661), .ZN(n830) );
  NOR2_X1 U923 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U924 ( .A(n832), .B(KEYINPUT109), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n833) );
  XNOR2_X1 U926 ( .A(KEYINPUT110), .B(n833), .ZN(n835) );
  NAND2_X1 U927 ( .A1(n835), .A2(n834), .ZN(G188) );
  INV_X1 U929 ( .A(G120), .ZN(G236) );
  INV_X1 U930 ( .A(G108), .ZN(G238) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  INV_X1 U932 ( .A(G69), .ZN(G235) );
  NOR2_X1 U933 ( .A1(n837), .A2(n836), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  XOR2_X1 U935 ( .A(G2100), .B(G2096), .Z(n839) );
  XNOR2_X1 U936 ( .A(KEYINPUT42), .B(G2678), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U938 ( .A(KEYINPUT43), .B(G2090), .Z(n841) );
  XNOR2_X1 U939 ( .A(G2067), .B(G2072), .ZN(n840) );
  XNOR2_X1 U940 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U941 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U942 ( .A(G2078), .B(G2084), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(G227) );
  XOR2_X1 U944 ( .A(G1971), .B(G1961), .Z(n847) );
  XNOR2_X1 U945 ( .A(G1986), .B(G1966), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U947 ( .A(G1956), .B(G1981), .Z(n849) );
  XNOR2_X1 U948 ( .A(G1996), .B(G1991), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U950 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U951 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(n855) );
  XOR2_X1 U953 ( .A(G1976), .B(G2474), .Z(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(G229) );
  INV_X1 U955 ( .A(n856), .ZN(G319) );
  NAND2_X1 U956 ( .A1(G124), .A2(n883), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n857), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U958 ( .A1(G100), .A2(n886), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n858), .B(KEYINPUT112), .ZN(n859) );
  NAND2_X1 U960 ( .A1(n860), .A2(n859), .ZN(n864) );
  NAND2_X1 U961 ( .A1(G112), .A2(n882), .ZN(n862) );
  NAND2_X1 U962 ( .A1(G136), .A2(n887), .ZN(n861) );
  NAND2_X1 U963 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U964 ( .A1(n864), .A2(n863), .ZN(G162) );
  XNOR2_X1 U965 ( .A(KEYINPUT46), .B(KEYINPUT114), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n865), .B(KEYINPUT48), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n867), .B(n866), .ZN(n878) );
  NAND2_X1 U968 ( .A1(G103), .A2(n886), .ZN(n869) );
  NAND2_X1 U969 ( .A1(G139), .A2(n887), .ZN(n868) );
  NAND2_X1 U970 ( .A1(n869), .A2(n868), .ZN(n875) );
  NAND2_X1 U971 ( .A1(G115), .A2(n882), .ZN(n871) );
  NAND2_X1 U972 ( .A1(G127), .A2(n883), .ZN(n870) );
  NAND2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U974 ( .A(KEYINPUT113), .B(n872), .ZN(n873) );
  XNOR2_X1 U975 ( .A(KEYINPUT47), .B(n873), .ZN(n874) );
  NOR2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n998) );
  XOR2_X1 U977 ( .A(G164), .B(n998), .Z(n876) );
  XNOR2_X1 U978 ( .A(G160), .B(n876), .ZN(n877) );
  XNOR2_X1 U979 ( .A(n878), .B(n877), .ZN(n881) );
  XNOR2_X1 U980 ( .A(n879), .B(n996), .ZN(n880) );
  XNOR2_X1 U981 ( .A(n881), .B(n880), .ZN(n897) );
  NAND2_X1 U982 ( .A1(G118), .A2(n882), .ZN(n885) );
  NAND2_X1 U983 ( .A1(G130), .A2(n883), .ZN(n884) );
  NAND2_X1 U984 ( .A1(n885), .A2(n884), .ZN(n892) );
  NAND2_X1 U985 ( .A1(G106), .A2(n886), .ZN(n889) );
  NAND2_X1 U986 ( .A1(G142), .A2(n887), .ZN(n888) );
  NAND2_X1 U987 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U988 ( .A(n890), .B(KEYINPUT45), .Z(n891) );
  NOR2_X1 U989 ( .A1(n892), .A2(n891), .ZN(n894) );
  XNOR2_X1 U990 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U991 ( .A(G162), .B(n895), .Z(n896) );
  XNOR2_X1 U992 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U993 ( .A1(G37), .A2(n898), .ZN(n899) );
  XOR2_X1 U994 ( .A(KEYINPUT115), .B(n899), .Z(G395) );
  XOR2_X1 U995 ( .A(n900), .B(G286), .Z(n902) );
  XNOR2_X1 U996 ( .A(G171), .B(n941), .ZN(n901) );
  XNOR2_X1 U997 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U998 ( .A1(G37), .A2(n903), .ZN(G397) );
  NOR2_X1 U999 ( .A1(G227), .A2(G229), .ZN(n905) );
  XNOR2_X1 U1000 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n918) );
  XNOR2_X1 U1002 ( .A(G2451), .B(G2427), .ZN(n915) );
  XOR2_X1 U1003 ( .A(KEYINPUT107), .B(G2443), .Z(n907) );
  XNOR2_X1 U1004 ( .A(G2435), .B(G2438), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n911) );
  XOR2_X1 U1006 ( .A(G2454), .B(G2430), .Z(n909) );
  XNOR2_X1 U1007 ( .A(G1348), .B(G1341), .ZN(n908) );
  XNOR2_X1 U1008 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1009 ( .A(n911), .B(n910), .Z(n913) );
  XNOR2_X1 U1010 ( .A(G2446), .B(KEYINPUT108), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(n915), .B(n914), .ZN(n916) );
  NAND2_X1 U1013 ( .A1(n916), .A2(G14), .ZN(n921) );
  NAND2_X1 U1014 ( .A1(G319), .A2(n921), .ZN(n917) );
  NOR2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n919) );
  NAND2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(n921), .ZN(G401) );
  XNOR2_X1 U1020 ( .A(KEYINPUT56), .B(G16), .ZN(n947) );
  XNOR2_X1 U1021 ( .A(n922), .B(G1956), .ZN(n924) );
  NAND2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n927) );
  XOR2_X1 U1023 ( .A(G1971), .B(G166), .Z(n925) );
  XNOR2_X1 U1024 ( .A(KEYINPUT124), .B(n925), .ZN(n926) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n934) );
  XNOR2_X1 U1026 ( .A(n928), .B(KEYINPUT123), .ZN(n930) );
  XNOR2_X1 U1027 ( .A(G171), .B(G1961), .ZN(n929) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n940) );
  XNOR2_X1 U1031 ( .A(G1966), .B(G168), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(n935), .B(KEYINPUT122), .ZN(n936) );
  NAND2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1034 ( .A(KEYINPUT57), .B(n938), .Z(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n945) );
  XOR2_X1 U1036 ( .A(n694), .B(G1341), .Z(n943) );
  XOR2_X1 U1037 ( .A(G1348), .B(n941), .Z(n942) );
  NOR2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n1025) );
  XNOR2_X1 U1041 ( .A(n948), .B(G20), .ZN(n956) );
  XOR2_X1 U1042 ( .A(G1981), .B(G6), .Z(n951) );
  XOR2_X1 U1043 ( .A(G19), .B(KEYINPUT126), .Z(n949) );
  XNOR2_X1 U1044 ( .A(G1341), .B(n949), .ZN(n950) );
  NAND2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n954) );
  XOR2_X1 U1046 ( .A(KEYINPUT59), .B(G1348), .Z(n952) );
  XNOR2_X1 U1047 ( .A(G4), .B(n952), .ZN(n953) );
  NOR2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(n957), .B(KEYINPUT60), .ZN(n969) );
  XNOR2_X1 U1051 ( .A(G1986), .B(G24), .ZN(n962) );
  XNOR2_X1 U1052 ( .A(G1971), .B(G22), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(G1976), .B(G23), .ZN(n958) );
  NOR2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(KEYINPUT127), .B(n960), .ZN(n961) );
  NOR2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(KEYINPUT58), .B(n963), .ZN(n967) );
  XNOR2_X1 U1058 ( .A(G1966), .B(G21), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(G1961), .B(G5), .ZN(n964) );
  NOR2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(n970), .B(KEYINPUT61), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(G16), .B(KEYINPUT125), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(G11), .A2(n973), .ZN(n1023) );
  XOR2_X1 U1067 ( .A(G1991), .B(G25), .Z(n974) );
  NAND2_X1 U1068 ( .A1(n974), .A2(G28), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(G32), .B(G1996), .ZN(n975) );
  NOR2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n984) );
  XOR2_X1 U1071 ( .A(n977), .B(G27), .Z(n982) );
  XNOR2_X1 U1072 ( .A(G2067), .B(G26), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(G2072), .B(G33), .ZN(n978) );
  NOR2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(KEYINPUT119), .B(n980), .ZN(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(KEYINPUT53), .B(n985), .ZN(n989) );
  XOR2_X1 U1079 ( .A(KEYINPUT120), .B(G34), .Z(n987) );
  XNOR2_X1 U1080 ( .A(G2084), .B(KEYINPUT54), .ZN(n986) );
  XNOR2_X1 U1081 ( .A(n987), .B(n986), .ZN(n988) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(KEYINPUT118), .B(G2090), .ZN(n990) );
  XNOR2_X1 U1084 ( .A(G35), .B(n990), .ZN(n991) );
  NOR2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1086 ( .A(KEYINPUT121), .B(n993), .Z(n994) );
  NOR2_X1 U1087 ( .A1(G29), .A2(n994), .ZN(n995) );
  XNOR2_X1 U1088 ( .A(n995), .B(KEYINPUT55), .ZN(n1021) );
  NOR2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n1007) );
  XOR2_X1 U1090 ( .A(G2072), .B(n998), .Z(n1000) );
  XOR2_X1 U1091 ( .A(G164), .B(G2078), .Z(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1093 ( .A(KEYINPUT50), .B(n1001), .ZN(n1003) );
  XNOR2_X1 U1094 ( .A(G160), .B(G2084), .ZN(n1002) );
  NAND2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(G2090), .B(G162), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(n1010), .B(KEYINPUT51), .ZN(n1011) );
  XNOR2_X1 U1101 ( .A(n1011), .B(KEYINPUT117), .ZN(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1105 ( .A(KEYINPUT52), .B(n1018), .Z(n1019) );
  NAND2_X1 U1106 ( .A1(G29), .A2(n1019), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1026), .Z(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

