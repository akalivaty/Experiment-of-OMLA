//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975;
  INV_X1    g000(.A(KEYINPUT18), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT17), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT14), .ZN(new_n204));
  NOR3_X1   g003(.A1(new_n204), .A2(G29gat), .A3(G36gat), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  INV_X1    g005(.A(G36gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(new_n206), .B2(new_n207), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n205), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT15), .ZN(new_n211));
  XOR2_X1   g010(.A(G43gat), .B(G50gat), .Z(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n211), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n210), .A2(KEYINPUT15), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n203), .B(new_n213), .C1(new_n216), .C2(new_n212), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n209), .A2(new_n208), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(new_n204), .B2(new_n208), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT15), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n212), .B1(new_n221), .B2(new_n211), .ZN(new_n222));
  INV_X1    g021(.A(new_n213), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT17), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(G15gat), .B(G22gat), .Z(new_n225));
  INV_X1    g024(.A(G1gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT87), .ZN(new_n228));
  AOI21_X1  g027(.A(G8gat), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT16), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n230), .A2(G1gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n227), .B1(new_n231), .B2(new_n225), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n229), .B(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n224), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n233), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n222), .A2(new_n223), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(G229gat), .A2(G233gat), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n202), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n233), .B1(new_n222), .B2(new_n223), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n239), .B(KEYINPUT13), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n234), .A2(new_n237), .A3(KEYINPUT18), .A4(new_n239), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n241), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(G169gat), .B(G197gat), .Z(new_n249));
  XNOR2_X1  g048(.A(G113gat), .B(G141gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g050(.A(KEYINPUT86), .B(KEYINPUT11), .Z(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n253), .B(KEYINPUT12), .Z(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n248), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n248), .A2(new_n255), .ZN(new_n258));
  AND2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G227gat), .A2(G233gat), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT28), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT27), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n263), .A2(G183gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT66), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n265), .A2(new_n263), .A3(G183gat), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n264), .B1(new_n266), .B2(KEYINPUT65), .ZN(new_n267));
  INV_X1    g066(.A(G183gat), .ZN(new_n268));
  OAI211_X1 g067(.A(KEYINPUT65), .B(KEYINPUT27), .C1(new_n268), .C2(KEYINPUT66), .ZN(new_n269));
  INV_X1    g068(.A(G190gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n262), .B1(new_n267), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT67), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT27), .B(G183gat), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n274), .A2(KEYINPUT28), .A3(new_n270), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n276), .B(new_n262), .C1(new_n267), .C2(new_n271), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n273), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT26), .ZN(new_n280));
  NAND2_X1  g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n280), .A2(new_n281), .B1(G183gat), .B2(G190gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n270), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G190gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n281), .B(new_n284), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT23), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n279), .B(new_n290), .ZN(new_n291));
  OR2_X1    g090(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n292));
  NAND2_X1  g091(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n289), .A2(new_n291), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n279), .B(KEYINPUT23), .ZN(new_n295));
  OAI211_X1 g094(.A(KEYINPUT64), .B(KEYINPUT25), .C1(new_n295), .C2(new_n288), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G127gat), .ZN(new_n300));
  INV_X1    g099(.A(G134gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G127gat), .A2(G134gat), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT1), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G120gat), .ZN(new_n305));
  OR2_X1    g104(.A1(KEYINPUT70), .A2(G113gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(KEYINPUT70), .A2(G113gat), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G113gat), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT69), .B1(new_n309), .B2(G120gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT69), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n311), .A2(new_n305), .A3(G113gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n304), .B1(new_n308), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT71), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n301), .A2(KEYINPUT68), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT68), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G134gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n316), .A2(new_n318), .A3(G127gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(G113gat), .B(G120gat), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n319), .B(new_n302), .C1(KEYINPUT1), .C2(new_n320), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n314), .A2(new_n315), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n315), .B1(new_n314), .B2(new_n321), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n299), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n297), .B1(new_n278), .B2(new_n282), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(new_n324), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n261), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n326), .A2(new_n261), .A3(new_n328), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT34), .B1(new_n261), .B2(KEYINPUT73), .ZN(new_n331));
  AND3_X1   g130(.A1(new_n330), .A2(KEYINPUT32), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n331), .B1(new_n330), .B2(KEYINPUT32), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n329), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G15gat), .B(G43gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n335), .B(KEYINPUT72), .ZN(new_n336));
  XOR2_X1   g135(.A(G71gat), .B(G99gat), .Z(new_n337));
  XOR2_X1   g136(.A(new_n336), .B(new_n337), .Z(new_n338));
  AND3_X1   g137(.A1(new_n283), .A2(new_n324), .A3(new_n298), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n324), .B1(new_n283), .B2(new_n298), .ZN(new_n340));
  NOR3_X1   g139(.A1(new_n339), .A2(new_n340), .A3(new_n260), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n338), .B1(new_n341), .B2(KEYINPUT33), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n331), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT32), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n344), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n330), .A2(KEYINPUT32), .A3(new_n331), .ZN(new_n347));
  INV_X1    g146(.A(new_n329), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n334), .A2(new_n343), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n343), .B1(new_n334), .B2(new_n349), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G22gat), .B(G50gat), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  XOR2_X1   g153(.A(G78gat), .B(G106gat), .Z(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT31), .ZN(new_n357));
  NAND2_X1  g156(.A1(G228gat), .A2(G233gat), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G197gat), .B(G204gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT22), .ZN(new_n361));
  NAND2_X1  g160(.A1(G211gat), .A2(G218gat), .ZN(new_n362));
  INV_X1    g161(.A(G211gat), .ZN(new_n363));
  INV_X1    g162(.A(G218gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n361), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT22), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n362), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n360), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT74), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G155gat), .A2(G162gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT2), .ZN(new_n374));
  INV_X1    g173(.A(G148gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n375), .A2(G141gat), .ZN(new_n376));
  INV_X1    g175(.A(G141gat), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n377), .A2(G148gat), .ZN(new_n378));
  OAI211_X1 g177(.A(KEYINPUT79), .B(new_n374), .C1(new_n376), .C2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G155gat), .B(G162gat), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT3), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n377), .A2(G148gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n375), .A2(G141gat), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(new_n380), .A3(new_n374), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n382), .A2(new_n383), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT29), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n372), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n382), .A2(new_n388), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n370), .A2(new_n390), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n395), .B1(new_n396), .B2(new_n383), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n359), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n370), .B(KEYINPUT74), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n391), .ZN(new_n400));
  OR2_X1    g199(.A1(new_n366), .A2(KEYINPUT83), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n366), .A2(KEYINPUT83), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(new_n369), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT3), .B1(new_n403), .B2(new_n390), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n400), .B(new_n358), .C1(new_n404), .C2(new_n395), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n357), .B1(new_n398), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n398), .A2(new_n405), .A3(new_n357), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n356), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n408), .ZN(new_n410));
  NOR3_X1   g209(.A1(new_n410), .A2(new_n406), .A3(new_n355), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n354), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n407), .A2(new_n408), .A3(new_n356), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n355), .B1(new_n410), .B2(new_n406), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n413), .A2(new_n414), .A3(new_n353), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n352), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT5), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n314), .A2(new_n321), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n394), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n314), .A2(new_n382), .A3(new_n321), .A4(new_n388), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(KEYINPUT80), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT81), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT81), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n422), .A2(new_n428), .A3(new_n425), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n418), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  OAI211_X1 g229(.A(KEYINPUT4), .B(new_n395), .C1(new_n322), .C2(new_n323), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n394), .A2(KEYINPUT3), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n432), .A2(new_n419), .A3(new_n389), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n433), .A2(KEYINPUT4), .ZN(new_n434));
  INV_X1    g233(.A(new_n421), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n431), .B(new_n424), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(KEYINPUT4), .ZN(new_n437));
  INV_X1    g236(.A(new_n323), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n314), .A2(new_n321), .A3(new_n315), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n394), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n433), .B(new_n437), .C1(new_n440), .C2(KEYINPUT4), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n425), .A2(KEYINPUT5), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n430), .A2(new_n436), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n445));
  XNOR2_X1  g244(.A(G1gat), .B(G29gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(G57gat), .B(G85gat), .ZN(new_n448));
  XOR2_X1   g247(.A(new_n447), .B(new_n448), .Z(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT6), .B1(new_n444), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT4), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n452), .B1(new_n324), .B2(new_n394), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n453), .A2(new_n433), .A3(new_n437), .A4(new_n443), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n435), .B1(new_n433), .B2(KEYINPUT4), .ZN(new_n455));
  INV_X1    g254(.A(new_n431), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n455), .A2(new_n456), .A3(new_n425), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n428), .B1(new_n422), .B2(new_n425), .ZN(new_n458));
  AOI211_X1 g257(.A(KEYINPUT81), .B(new_n424), .C1(new_n420), .C2(new_n421), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT5), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n454), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n449), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n451), .B(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT78), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT76), .ZN(new_n465));
  NAND2_X1  g264(.A1(G226gat), .A2(G233gat), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n299), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n466), .B(KEYINPUT75), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n469), .B1(new_n327), .B2(KEYINPUT29), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n465), .B1(new_n471), .B2(new_n399), .ZN(new_n472));
  AOI211_X1 g271(.A(KEYINPUT76), .B(new_n372), .C1(new_n468), .C2(new_n470), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n469), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n299), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n466), .B1(new_n327), .B2(KEYINPUT29), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(new_n477), .A3(new_n372), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT77), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT77), .A4(new_n372), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT30), .ZN(new_n483));
  XOR2_X1   g282(.A(G8gat), .B(G36gat), .Z(new_n484));
  XNOR2_X1  g283(.A(new_n484), .B(G64gat), .ZN(new_n485));
  INV_X1    g284(.A(G92gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  NOR4_X1   g286(.A1(new_n474), .A2(new_n482), .A3(new_n483), .A4(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n487), .ZN(new_n489));
  INV_X1    g288(.A(new_n472), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n471), .A2(new_n465), .A3(new_n399), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n482), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n489), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n464), .B1(new_n488), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT30), .A4(new_n489), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n480), .B(new_n481), .C1(new_n472), .C2(new_n473), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(new_n487), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n496), .A2(new_n498), .A3(KEYINPUT78), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n483), .B1(new_n497), .B2(new_n487), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n417), .A2(new_n463), .A3(new_n495), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT35), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT35), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n461), .A2(KEYINPUT85), .A3(new_n449), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT85), .B1(new_n461), .B2(new_n449), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n451), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n462), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AND4_X1   g309(.A1(new_n504), .A2(new_n352), .A3(new_n416), .A4(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n500), .A2(new_n498), .A3(new_n496), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n503), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n487), .B1(new_n497), .B2(KEYINPUT37), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT37), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n517), .B1(new_n492), .B2(new_n493), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT38), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n492), .A2(new_n493), .A3(new_n489), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n507), .A2(new_n520), .A3(new_n509), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n476), .A2(new_n477), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n522), .A2(new_n372), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n523), .B1(new_n372), .B2(new_n471), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT38), .B1(new_n524), .B2(KEYINPUT37), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n525), .B(new_n487), .C1(KEYINPUT37), .C2(new_n497), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n519), .A2(new_n521), .A3(new_n526), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n505), .A2(new_n506), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n441), .A2(new_n425), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n529), .B(KEYINPUT39), .C1(new_n425), .C2(new_n422), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n530), .B(new_n450), .C1(KEYINPUT39), .C2(new_n529), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT40), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n512), .A2(new_n528), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n527), .A2(new_n416), .A3(new_n533), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n495), .A2(new_n463), .A3(new_n499), .A4(new_n500), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT84), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n413), .A2(new_n414), .A3(new_n353), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n353), .B1(new_n413), .B2(new_n414), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n412), .A2(KEYINPUT84), .A3(new_n415), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT36), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n543), .B1(new_n350), .B2(new_n351), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n332), .A2(new_n333), .A3(new_n329), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n348), .B1(new_n346), .B2(new_n347), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n342), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n334), .A2(new_n343), .A3(new_n349), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(KEYINPUT36), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n544), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n542), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n259), .B1(new_n515), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT95), .ZN(new_n553));
  NAND2_X1  g352(.A1(G85gat), .A2(G92gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n554), .B(new_n555), .Z(new_n556));
  XOR2_X1   g355(.A(G99gat), .B(G106gat), .Z(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G99gat), .A2(G106gat), .ZN(new_n559));
  INV_X1    g358(.A(G85gat), .ZN(new_n560));
  AOI22_X1  g359(.A1(KEYINPUT8), .A2(new_n559), .B1(new_n560), .B2(new_n486), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n556), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT94), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n556), .A2(KEYINPUT94), .A3(new_n558), .A4(new_n561), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n556), .A2(new_n561), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(new_n557), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n217), .A2(new_n224), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n236), .A2(new_n568), .A3(new_n566), .ZN(new_n571));
  NAND2_X1  g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT92), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT41), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n570), .A2(new_n571), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(G190gat), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n570), .A2(new_n571), .A3(new_n270), .A4(new_n575), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n577), .A2(G218gat), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(G218gat), .B1(new_n577), .B2(new_n578), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n553), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n577), .A2(new_n578), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(new_n364), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n577), .A2(G218gat), .A3(new_n578), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n583), .A2(KEYINPUT95), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n573), .A2(new_n574), .ZN(new_n586));
  XOR2_X1   g385(.A(G134gat), .B(G162gat), .Z(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n581), .A2(new_n585), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n588), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n553), .B(new_n590), .C1(new_n579), .C2(new_n580), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n552), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(KEYINPUT89), .A2(G57gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(G64gat), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT9), .ZN(new_n596));
  INV_X1    g395(.A(G71gat), .ZN(new_n597));
  INV_X1    g396(.A(G78gat), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT90), .ZN(new_n600));
  XNOR2_X1  g399(.A(G71gat), .B(G78gat), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT90), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n602), .B(new_n596), .C1(new_n597), .C2(new_n598), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n595), .A2(new_n600), .A3(new_n601), .A4(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT91), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT88), .B(G57gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(G64gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(new_n599), .ZN(new_n609));
  INV_X1    g408(.A(new_n601), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n613), .A2(KEYINPUT21), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(G127gat), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT21), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n233), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n614), .B(new_n300), .ZN(new_n619));
  INV_X1    g418(.A(new_n617), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n623));
  XNOR2_X1  g422(.A(G155gat), .B(G183gat), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n623), .B(new_n624), .Z(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G231gat), .A2(G233gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(new_n363), .ZN(new_n628));
  INV_X1    g427(.A(new_n625), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n618), .A2(new_n621), .A3(new_n629), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n626), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n628), .B1(new_n626), .B2(new_n630), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n612), .A2(new_n569), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n606), .A2(new_n611), .A3(new_n568), .A4(new_n562), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n613), .A2(KEYINPUT10), .A3(new_n568), .A4(new_n566), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G230gat), .A2(G233gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT98), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n634), .A2(new_n636), .ZN(new_n643));
  INV_X1    g442(.A(new_n640), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT98), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n639), .A2(new_n646), .A3(new_n640), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n642), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(G120gat), .B(G148gat), .ZN(new_n649));
  INV_X1    g448(.A(G176gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(G204gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n637), .A2(new_n638), .A3(KEYINPUT96), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT96), .B1(new_n637), .B2(new_n638), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n640), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n653), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n645), .A2(KEYINPUT97), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n645), .A2(KEYINPUT97), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n657), .A2(new_n658), .A3(new_n659), .A4(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n654), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n633), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n593), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(new_n463), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(new_n226), .ZN(G1324gat));
  AND2_X1   g465(.A1(new_n593), .A2(new_n663), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n512), .ZN(new_n668));
  INV_X1    g467(.A(G8gat), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n230), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n230), .A2(new_n669), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT42), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n671), .A2(new_n672), .B1(G8gat), .B2(new_n668), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n675), .B1(new_n676), .B2(new_n674), .ZN(G1325gat));
  INV_X1    g476(.A(new_n352), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n664), .A2(new_n678), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n544), .A2(KEYINPUT99), .A3(new_n549), .ZN(new_n680));
  AOI21_X1  g479(.A(KEYINPUT99), .B1(new_n544), .B2(new_n549), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(G15gat), .ZN(new_n683));
  OAI22_X1  g482(.A1(new_n679), .A2(G15gat), .B1(new_n664), .B2(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT100), .Z(G1326gat));
  INV_X1    g484(.A(new_n541), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n664), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT43), .B(G22gat), .Z(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1327gat));
  NOR2_X1   g488(.A1(new_n631), .A2(new_n632), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(new_n662), .ZN(new_n691));
  INV_X1    g490(.A(new_n592), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n694), .A2(KEYINPUT101), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(KEYINPUT101), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n552), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n451), .B(new_n508), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n697), .A2(new_n206), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT45), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701));
  AOI22_X1  g500(.A1(new_n502), .A2(KEYINPUT35), .B1(new_n513), .B2(new_n511), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n534), .A2(new_n542), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT102), .B1(new_n703), .B2(new_n682), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT99), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n550), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n544), .A2(KEYINPUT99), .A3(new_n549), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT102), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n708), .A2(new_n709), .A3(new_n542), .A4(new_n534), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n702), .B1(new_n704), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n701), .B1(new_n711), .B2(new_n592), .ZN(new_n712));
  INV_X1    g511(.A(new_n259), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n515), .A2(new_n551), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n714), .A2(KEYINPUT44), .A3(new_n692), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n712), .A2(new_n713), .A3(new_n691), .A4(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G29gat), .B1(new_n716), .B2(new_n463), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n700), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT103), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n700), .A2(KEYINPUT103), .A3(new_n717), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(G1328gat));
  NAND3_X1  g521(.A1(new_n697), .A2(new_n207), .A3(new_n512), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n723), .B1(KEYINPUT104), .B2(KEYINPUT46), .ZN(new_n724));
  OR2_X1    g523(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(G36gat), .B1(new_n716), .B2(new_n513), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(G1329gat));
  OR3_X1    g527(.A1(new_n716), .A2(KEYINPUT105), .A3(new_n708), .ZN(new_n729));
  OAI21_X1  g528(.A(KEYINPUT105), .B1(new_n716), .B2(new_n708), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n729), .A2(G43gat), .A3(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n697), .ZN(new_n732));
  OR3_X1    g531(.A1(new_n732), .A2(G43gat), .A3(new_n678), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT47), .ZN(new_n734));
  OAI21_X1  g533(.A(G43gat), .B1(new_n716), .B2(new_n708), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  OAI22_X1  g535(.A1(new_n731), .A2(new_n734), .B1(KEYINPUT47), .B2(new_n736), .ZN(G1330gat));
  NOR3_X1   g536(.A1(new_n732), .A2(G50gat), .A3(new_n686), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(G50gat), .B1(new_n716), .B2(new_n416), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n739), .A2(KEYINPUT48), .A3(new_n740), .ZN(new_n741));
  OR2_X1    g540(.A1(new_n716), .A2(new_n686), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n738), .B1(new_n742), .B2(G50gat), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n741), .B1(new_n743), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g543(.A1(new_n704), .A2(new_n710), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n515), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n592), .A2(new_n259), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n633), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n746), .A2(new_n662), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n749), .A2(new_n463), .ZN(new_n750));
  XNOR2_X1  g549(.A(KEYINPUT106), .B(G57gat), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1332gat));
  NOR2_X1   g551(.A1(new_n749), .A2(new_n513), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT49), .B(G64gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(new_n753), .B2(new_n756), .ZN(G1333gat));
  OAI21_X1  g556(.A(new_n597), .B1(new_n749), .B2(new_n678), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n746), .A2(G71gat), .A3(new_n662), .A4(new_n748), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n708), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT107), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n759), .A2(KEYINPUT107), .A3(new_n708), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n758), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g564(.A1(new_n749), .A2(new_n686), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(new_n598), .ZN(G1335gat));
  NOR2_X1   g566(.A1(new_n690), .A2(new_n713), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n662), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n712), .A2(new_n715), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(G85gat), .B1(new_n772), .B2(new_n463), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n592), .B1(new_n745), .B2(new_n515), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT51), .B1(new_n774), .B2(new_n768), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT51), .ZN(new_n776));
  NOR4_X1   g575(.A1(new_n711), .A2(new_n776), .A3(new_n592), .A4(new_n769), .ZN(new_n777));
  OR3_X1    g576(.A1(new_n775), .A2(new_n777), .A3(KEYINPUT108), .ZN(new_n778));
  OAI21_X1  g577(.A(KEYINPUT108), .B1(new_n775), .B2(new_n777), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n780), .A2(new_n560), .A3(new_n662), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n773), .B1(new_n781), .B2(new_n463), .ZN(G1336gat));
  OAI21_X1  g581(.A(G92gat), .B1(new_n772), .B2(new_n513), .ZN(new_n783));
  NAND2_X1  g582(.A1(KEYINPUT110), .A2(KEYINPUT52), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n512), .A2(new_n486), .A3(new_n662), .ZN(new_n785));
  XOR2_X1   g584(.A(new_n785), .B(KEYINPUT109), .Z(new_n786));
  OAI21_X1  g585(.A(new_n786), .B1(new_n775), .B2(new_n777), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n783), .A2(new_n784), .A3(new_n787), .ZN(new_n788));
  OR2_X1    g587(.A1(KEYINPUT110), .A2(KEYINPUT52), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(G1337gat));
  OAI21_X1  g589(.A(G99gat), .B1(new_n772), .B2(new_n708), .ZN(new_n791));
  INV_X1    g590(.A(G99gat), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n780), .A2(new_n792), .A3(new_n662), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n793), .B2(new_n678), .ZN(G1338gat));
  NOR3_X1   g593(.A1(new_n770), .A2(new_n416), .A3(G106gat), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(new_n775), .B2(new_n777), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT112), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n712), .A2(new_n541), .A3(new_n715), .A4(new_n771), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(G106gat), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(KEYINPUT111), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT111), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n799), .A2(new_n802), .A3(G106gat), .ZN(new_n803));
  OAI211_X1 g602(.A(KEYINPUT112), .B(new_n795), .C1(new_n775), .C2(new_n777), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n798), .A2(new_n801), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(KEYINPUT53), .ZN(new_n806));
  OAI21_X1  g605(.A(G106gat), .B1(new_n772), .B2(new_n416), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(new_n808), .A3(new_n796), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n806), .A2(new_n809), .ZN(G1339gat));
  NOR3_X1   g609(.A1(new_n633), .A2(new_n662), .A3(new_n747), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n812), .B1(new_n238), .B2(new_n240), .ZN(new_n813));
  AOI211_X1 g612(.A(KEYINPUT114), .B(new_n239), .C1(new_n234), .C2(new_n237), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n243), .A2(new_n245), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(new_n253), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n817), .A2(new_n256), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n592), .A2(new_n662), .A3(new_n818), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n589), .B(new_n591), .C1(new_n256), .C2(new_n817), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n637), .A2(new_n638), .A3(new_n644), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n657), .A2(KEYINPUT54), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT54), .B1(new_n642), .B2(new_n647), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT113), .B1(new_n824), .B2(new_n658), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n646), .B1(new_n639), .B2(new_n640), .ZN(new_n827));
  AOI211_X1 g626(.A(KEYINPUT98), .B(new_n644), .C1(new_n637), .C2(new_n638), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(new_n830), .A3(new_n653), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n823), .B1(new_n825), .B2(new_n831), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n820), .B(new_n661), .C1(new_n832), .C2(KEYINPUT55), .ZN(new_n833));
  INV_X1    g632(.A(new_n831), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n830), .B1(new_n829), .B2(new_n653), .ZN(new_n835));
  OAI211_X1 g634(.A(KEYINPUT55), .B(new_n822), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n747), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n819), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n811), .B1(new_n838), .B2(new_n633), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n839), .A2(new_n463), .A3(new_n512), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n840), .A2(new_n417), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n259), .B1(new_n306), .B2(new_n307), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n839), .A2(new_n541), .A3(new_n678), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n512), .A2(new_n463), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(G113gat), .B1(new_n846), .B2(new_n259), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n843), .A2(new_n847), .ZN(G1340gat));
  OAI21_X1  g647(.A(G120gat), .B1(new_n846), .B2(new_n770), .ZN(new_n849));
  INV_X1    g648(.A(new_n841), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n662), .A2(new_n305), .ZN(new_n851));
  XOR2_X1   g650(.A(new_n851), .B(KEYINPUT115), .Z(new_n852));
  OAI21_X1  g651(.A(new_n849), .B1(new_n850), .B2(new_n852), .ZN(G1341gat));
  AOI21_X1  g652(.A(G127gat), .B1(new_n841), .B2(new_n690), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n846), .A2(new_n300), .A3(new_n633), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n854), .A2(new_n855), .ZN(G1342gat));
  NAND2_X1  g655(.A1(new_n316), .A2(new_n318), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n841), .A2(new_n857), .A3(new_n692), .ZN(new_n858));
  XOR2_X1   g657(.A(new_n858), .B(KEYINPUT56), .Z(new_n859));
  OAI21_X1  g658(.A(G134gat), .B1(new_n846), .B2(new_n592), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(G1343gat));
  NOR2_X1   g660(.A1(new_n682), .A2(new_n416), .ZN(new_n862));
  AND4_X1   g661(.A1(new_n377), .A2(new_n840), .A3(new_n713), .A4(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n864), .B1(new_n839), .B2(new_n416), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT116), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n839), .A2(new_n686), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT57), .ZN(new_n869));
  OAI211_X1 g668(.A(KEYINPUT116), .B(new_n864), .C1(new_n839), .C2(new_n416), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n867), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n708), .A2(new_n845), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(new_n713), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n863), .B1(new_n873), .B2(G141gat), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n875), .B1(new_n873), .B2(G141gat), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n874), .A2(new_n876), .A3(KEYINPUT58), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n878));
  AOI221_X4 g677(.A(new_n863), .B1(new_n875), .B2(new_n878), .C1(new_n873), .C2(G141gat), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n877), .A2(new_n879), .ZN(G1344gat));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n840), .A2(new_n375), .A3(new_n662), .A4(new_n862), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n868), .A2(KEYINPUT57), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n839), .A2(new_n864), .A3(new_n416), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n662), .B(new_n872), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(G148gat), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n886), .A2(KEYINPUT59), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n662), .A3(new_n872), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n375), .A2(KEYINPUT59), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n881), .B(new_n882), .C1(new_n887), .C2(new_n890), .ZN(new_n891));
  AOI22_X1  g690(.A1(KEYINPUT59), .A2(new_n886), .B1(new_n888), .B2(new_n889), .ZN(new_n892));
  INV_X1    g691(.A(new_n882), .ZN(new_n893));
  OAI21_X1  g692(.A(KEYINPUT118), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n891), .A2(new_n894), .ZN(G1345gat));
  NAND2_X1  g694(.A1(new_n871), .A2(new_n872), .ZN(new_n896));
  INV_X1    g695(.A(G155gat), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n896), .A2(new_n897), .A3(new_n633), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n840), .A2(new_n690), .A3(new_n862), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n897), .B2(new_n899), .ZN(G1346gat));
  INV_X1    g699(.A(G162gat), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n896), .A2(new_n901), .A3(new_n592), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n840), .A2(new_n692), .A3(new_n862), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n901), .B2(new_n903), .ZN(G1347gat));
  NOR2_X1   g703(.A1(new_n513), .A2(new_n698), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n844), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(G169gat), .B1(new_n906), .B2(new_n259), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n838), .A2(new_n633), .ZN(new_n908));
  OAI211_X1 g707(.A(KEYINPUT119), .B(new_n463), .C1(new_n908), .C2(new_n811), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT119), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n910), .B1(new_n839), .B2(new_n698), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n513), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT120), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n912), .A2(new_n913), .A3(new_n417), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n912), .B2(new_n417), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n259), .A2(G169gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n907), .B1(new_n916), .B2(new_n917), .ZN(G1348gat));
  NAND2_X1  g717(.A1(new_n662), .A2(new_n650), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n912), .A2(new_n417), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT120), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n912), .A2(new_n913), .A3(new_n417), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n919), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(G176gat), .B1(new_n906), .B2(new_n770), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT121), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT121), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n927), .B(new_n924), .C1(new_n916), .C2(new_n919), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n926), .A2(new_n928), .ZN(G1349gat));
  INV_X1    g728(.A(KEYINPUT122), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n930), .B1(new_n906), .B2(new_n633), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n844), .A2(KEYINPUT122), .A3(new_n690), .A4(new_n905), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n931), .A2(G183gat), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n690), .A2(new_n274), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n933), .B(new_n934), .C1(new_n920), .C2(new_n935), .ZN(new_n936));
  OR2_X1    g735(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n936), .B(new_n937), .ZN(G1350gat));
  OAI21_X1  g737(.A(G190gat), .B1(new_n906), .B2(new_n592), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT61), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n692), .A2(new_n270), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n916), .B2(new_n941), .ZN(G1351gat));
  NOR2_X1   g741(.A1(new_n259), .A2(G197gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n912), .A2(KEYINPUT124), .A3(new_n862), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT124), .B1(new_n912), .B2(new_n862), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n883), .A2(new_n884), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n708), .A2(new_n905), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n949), .A2(new_n713), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(G197gat), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT125), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n947), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n954), .B1(new_n947), .B2(new_n953), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n955), .A2(new_n956), .ZN(G1352gat));
  NAND4_X1  g756(.A1(new_n912), .A2(new_n652), .A3(new_n662), .A4(new_n862), .ZN(new_n958));
  XOR2_X1   g757(.A(new_n958), .B(KEYINPUT62), .Z(new_n959));
  NOR3_X1   g758(.A1(new_n948), .A2(new_n770), .A3(new_n950), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n652), .B2(new_n960), .ZN(G1353gat));
  OAI211_X1 g760(.A(new_n363), .B(new_n690), .C1(new_n945), .C2(new_n946), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n948), .A2(new_n633), .A3(new_n950), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n963), .A2(new_n363), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n964), .A2(KEYINPUT63), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n964), .A2(KEYINPUT63), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n962), .B1(new_n965), .B2(new_n966), .ZN(G1354gat));
  NOR2_X1   g766(.A1(new_n948), .A2(new_n950), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n592), .A2(new_n364), .ZN(new_n970));
  OAI22_X1  g769(.A1(new_n968), .A2(KEYINPUT126), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n968), .A2(KEYINPUT126), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n970), .A2(new_n969), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n692), .B1(new_n945), .B2(new_n946), .ZN(new_n975));
  AOI22_X1  g774(.A1(new_n973), .A2(new_n974), .B1(new_n364), .B2(new_n975), .ZN(G1355gat));
endmodule


