//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1273, new_n1274;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(KEYINPUT64), .ZN(new_n203));
  NAND2_X1  g0003(.A1(G1), .A2(G20), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n203), .B1(new_n204), .B2(G13), .ZN(new_n205));
  INV_X1    g0005(.A(G13), .ZN(new_n206));
  NAND4_X1  g0006(.A1(new_n206), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  NAND2_X1  g0010(.A1(G107), .A2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(G116), .ZN(new_n212));
  INV_X1    g0012(.A(G270), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI22_X1  g0018(.A1(new_n215), .A2(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  XOR2_X1   g0019(.A(KEYINPUT65), .B(G244), .Z(new_n220));
  AOI211_X1 g0020(.A(new_n214), .B(new_n219), .C1(new_n220), .C2(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  INV_X1    g0023(.A(G97), .ZN(new_n224));
  INV_X1    g0024(.A(G257), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(G50), .ZN(new_n227));
  INV_X1    g0027(.A(G226), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n204), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT66), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT1), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  INV_X1    g0033(.A(G20), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NOR2_X1   g0035(.A1(G58), .A2(G68), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n237), .A2(G50), .ZN(new_n238));
  INV_X1    g0038(.A(new_n238), .ZN(new_n239));
  AOI211_X1 g0039(.A(new_n210), .B(new_n232), .C1(new_n235), .C2(new_n239), .ZN(G361));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n223), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G264), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n213), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G358));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G107), .B(G116), .Z(new_n252));
  XNOR2_X1  g0052(.A(G87), .B(G97), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G77), .ZN(new_n259));
  OAI22_X1  g0059(.A1(new_n256), .A2(new_n258), .B1(new_n234), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT69), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n234), .A2(G33), .ZN(new_n262));
  XOR2_X1   g0062(.A(KEYINPUT15), .B(G87), .Z(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n261), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n233), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G20), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n265), .A2(new_n267), .B1(G77), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n269), .A2(G13), .A3(G20), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n259), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n276), .B(KEYINPUT70), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G238), .A2(G1698), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n279), .B(new_n280), .C1(new_n223), .C2(G1698), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n281), .B(new_n282), .C1(G107), .C2(new_n279), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n269), .B1(G41), .B2(G45), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G274), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n282), .A2(new_n285), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n220), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n283), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(G179), .ZN(new_n290));
  INV_X1    g0090(.A(G169), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n290), .B1(new_n291), .B2(new_n289), .ZN(new_n292));
  AND2_X1   g0092(.A1(new_n278), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT13), .ZN(new_n294));
  INV_X1    g0094(.A(G33), .ZN(new_n295));
  INV_X1    g0095(.A(G41), .ZN(new_n296));
  OAI211_X1 g0096(.A(G1), .B(G13), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G1698), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n228), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n279), .B(new_n299), .C1(G232), .C2(new_n298), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G97), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n297), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G274), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n284), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n297), .A2(new_n284), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n306), .A2(new_n216), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n294), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  NOR4_X1   g0109(.A1(new_n302), .A2(KEYINPUT13), .A3(new_n307), .A4(new_n304), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G200), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT73), .B(KEYINPUT12), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n269), .A2(new_n215), .A3(G13), .A4(G20), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  XOR2_X1   g0116(.A(new_n316), .B(KEYINPUT74), .Z(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(KEYINPUT12), .B2(new_n315), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT68), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(new_n295), .B2(G20), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n234), .A2(KEYINPUT68), .A3(G33), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n322), .A2(G77), .B1(G50), .B2(new_n257), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(new_n234), .B2(G68), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT11), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n324), .A2(new_n325), .A3(new_n267), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n325), .B1(new_n324), .B2(new_n267), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n318), .B1(new_n215), .B2(new_n271), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G190), .ZN(new_n329));
  NOR3_X1   g0129(.A1(new_n309), .A2(new_n329), .A3(new_n310), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT14), .B1(new_n311), .B2(new_n291), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT14), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n333), .B(G169), .C1(new_n309), .C2(new_n310), .ZN(new_n334));
  INV_X1    g0134(.A(G179), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n332), .B(new_n334), .C1(new_n312), .C2(new_n335), .ZN(new_n336));
  AOI221_X4 g0136(.A(new_n293), .B1(new_n313), .B2(new_n331), .C1(new_n336), .C2(new_n328), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT16), .ZN(new_n338));
  OR2_X1    g0138(.A1(KEYINPUT3), .A2(G33), .ZN(new_n339));
  NAND2_X1  g0139(.A1(KEYINPUT3), .A2(G33), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n339), .A2(new_n234), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT7), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n339), .A2(KEYINPUT7), .A3(new_n234), .A4(new_n340), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n215), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n222), .A2(new_n215), .ZN(new_n346));
  OAI21_X1  g0146(.A(G20), .B1(new_n346), .B2(new_n236), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n257), .A2(G159), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n338), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  AND2_X1   g0150(.A1(KEYINPUT3), .A2(G33), .ZN(new_n351));
  NOR2_X1   g0151(.A1(KEYINPUT3), .A2(G33), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT7), .B1(new_n353), .B2(new_n234), .ZN(new_n354));
  NOR4_X1   g0154(.A1(new_n351), .A2(new_n352), .A3(new_n342), .A4(G20), .ZN(new_n355));
  OAI21_X1  g0155(.A(G68), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n349), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(KEYINPUT16), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n350), .A2(new_n358), .A3(new_n267), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT76), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n222), .A2(KEYINPUT8), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT8), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G58), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT67), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n361), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n222), .A2(KEYINPUT67), .A3(KEYINPUT8), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n274), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n272), .B2(new_n367), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n304), .B1(new_n287), .B2(G232), .ZN(new_n370));
  OR2_X1    g0170(.A1(G223), .A2(G1698), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n228), .A2(G1698), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n371), .B(new_n372), .C1(new_n351), .C2(new_n352), .ZN(new_n373));
  NAND2_X1  g0173(.A1(G33), .A2(G87), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n282), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n370), .A2(new_n376), .A3(new_n329), .ZN(new_n377));
  INV_X1    g0177(.A(G200), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n286), .B1(new_n306), .B2(new_n223), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n297), .B1(new_n373), .B2(new_n374), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n359), .A2(new_n360), .A3(new_n369), .A4(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT75), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n359), .A2(new_n384), .A3(new_n369), .A4(new_n382), .ZN(new_n385));
  AOI22_X1  g0185(.A1(KEYINPUT75), .A2(new_n383), .B1(new_n385), .B2(KEYINPUT17), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n383), .A2(KEYINPUT75), .A3(KEYINPUT17), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n370), .A2(new_n376), .A3(new_n335), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n379), .A2(new_n380), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n388), .B1(G169), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n359), .B2(new_n369), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n391), .A2(KEYINPUT18), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n391), .A2(KEYINPUT18), .ZN(new_n393));
  OAI22_X1  g0193(.A1(new_n386), .A2(new_n387), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n394), .A2(KEYINPUT77), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n298), .A2(G222), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G223), .A2(G1698), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n279), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n398), .B(new_n282), .C1(G77), .C2(new_n279), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n287), .A2(G226), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(new_n286), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n291), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(G179), .B2(new_n401), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n271), .A2(new_n227), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n274), .A2(G50), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n322), .A2(new_n365), .A3(new_n366), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n236), .A2(new_n227), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n409), .A2(G20), .B1(G150), .B2(new_n257), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n405), .B(new_n407), .C1(new_n411), .C2(new_n268), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n403), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT71), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT9), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n268), .B1(new_n408), .B2(new_n410), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n417), .A2(new_n406), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n416), .B1(new_n418), .B2(new_n405), .ZN(new_n419));
  NOR4_X1   g0219(.A1(new_n417), .A2(new_n404), .A3(KEYINPUT9), .A4(new_n406), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n415), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n412), .A2(KEYINPUT9), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n418), .A2(new_n416), .A3(new_n405), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(KEYINPUT71), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n401), .A2(G200), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n399), .A2(G190), .A3(new_n286), .A4(new_n400), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT10), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n421), .A2(new_n424), .A3(new_n428), .A4(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT72), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n419), .A2(new_n420), .ZN(new_n433));
  AOI21_X1  g0233(.A(KEYINPUT10), .B1(new_n433), .B2(KEYINPUT71), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n422), .A2(new_n423), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n427), .B1(new_n435), .B2(new_n415), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n436), .A3(KEYINPUT72), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT10), .B1(new_n433), .B2(new_n427), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n414), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n289), .A2(G200), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n289), .A2(new_n329), .ZN(new_n442));
  AND4_X1   g0242(.A1(new_n273), .A2(new_n277), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n443), .B1(new_n394), .B2(KEYINPUT77), .ZN(new_n444));
  AND4_X1   g0244(.A1(new_n337), .A2(new_n395), .A3(new_n440), .A4(new_n444), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n295), .A2(new_n212), .A3(G20), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT23), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(new_n234), .B2(G107), .ZN(new_n448));
  INV_X1    g0248(.A(G107), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(KEYINPUT23), .A3(G20), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n446), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT22), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n217), .A2(KEYINPUT84), .ZN(new_n453));
  AND4_X1   g0253(.A1(new_n452), .A2(new_n279), .A3(new_n234), .A4(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(G20), .B1(new_n339), .B2(new_n340), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n452), .B1(new_n455), .B2(new_n453), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n451), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT24), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(KEYINPUT24), .B(new_n451), .C1(new_n454), .C2(new_n456), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(new_n267), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT85), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n462), .B(KEYINPUT25), .C1(new_n274), .C2(G107), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n269), .A2(G33), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n268), .A2(new_n274), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G107), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n461), .A2(new_n463), .A3(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n279), .B1(G257), .B2(new_n298), .ZN(new_n469));
  NOR2_X1   g0269(.A1(G250), .A2(G1698), .ZN(new_n470));
  INV_X1    g0270(.A(G294), .ZN(new_n471));
  OAI22_X1  g0271(.A1(new_n469), .A2(new_n470), .B1(new_n295), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G45), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(G1), .ZN(new_n474));
  AND2_X1   g0274(.A1(KEYINPUT5), .A2(G41), .ZN(new_n475));
  NOR2_X1   g0275(.A1(KEYINPUT5), .A2(G41), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AND2_X1   g0277(.A1(new_n477), .A2(new_n297), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n472), .A2(new_n282), .B1(G264), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n474), .B(G274), .C1(new_n476), .C2(new_n475), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G200), .ZN(new_n482));
  INV_X1    g0282(.A(new_n481), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G190), .ZN(new_n484));
  OR2_X1    g0284(.A1(new_n462), .A2(KEYINPUT25), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n462), .A2(KEYINPUT25), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n275), .A2(new_n485), .A3(new_n449), .A4(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n468), .A2(new_n482), .A3(new_n484), .A4(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n449), .A2(KEYINPUT6), .A3(G97), .ZN(new_n489));
  XOR2_X1   g0289(.A(G97), .B(G107), .Z(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(new_n490), .B2(KEYINPUT6), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n491), .A2(G20), .B1(G77), .B2(new_n257), .ZN(new_n492));
  OAI21_X1  g0292(.A(G107), .B1(new_n354), .B2(new_n355), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n268), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n465), .A2(new_n224), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n274), .A2(G97), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT78), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n279), .A2(KEYINPUT4), .A3(G244), .A4(new_n298), .ZN(new_n500));
  OAI21_X1  g0300(.A(G244), .B1(new_n351), .B2(new_n352), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT4), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G283), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n500), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n279), .A2(G250), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n298), .B1(new_n506), .B2(KEYINPUT4), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n499), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(KEYINPUT4), .B1(new_n353), .B2(new_n218), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G1698), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n501), .A2(new_n502), .B1(G33), .B2(G283), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n510), .A2(KEYINPUT78), .A3(new_n511), .A4(new_n500), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n508), .A2(new_n282), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n480), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n514), .B1(new_n478), .B2(G257), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n291), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n498), .B(new_n517), .C1(G179), .C2(new_n516), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n513), .A2(G190), .A3(new_n515), .ZN(new_n519));
  INV_X1    g0319(.A(new_n516), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n497), .B(new_n519), .C1(new_n520), .C2(new_n378), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n488), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n263), .A2(new_n274), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT19), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n234), .B1(new_n301), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(G97), .A2(G107), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n217), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT81), .ZN(new_n529));
  XNOR2_X1  g0329(.A(new_n528), .B(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n455), .A2(G68), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n524), .B1(new_n262), .B2(new_n224), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n523), .B1(new_n534), .B2(new_n267), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n264), .B2(new_n465), .ZN(new_n536));
  OAI211_X1 g0336(.A(G244), .B(G1698), .C1(new_n351), .C2(new_n352), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT79), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT79), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n279), .A2(new_n539), .A3(G244), .A4(G1698), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(G1698), .B1(new_n339), .B2(new_n340), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n542), .A2(G238), .B1(G33), .B2(G116), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n541), .A2(KEYINPUT80), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT80), .B1(new_n541), .B2(new_n543), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n282), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n474), .A2(new_n303), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n547), .B(new_n297), .C1(G250), .C2(new_n474), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n335), .A3(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n548), .ZN(new_n550));
  INV_X1    g0350(.A(G244), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n339), .B2(new_n340), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n539), .B1(new_n552), .B2(G1698), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n537), .A2(KEYINPUT79), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n543), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT80), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n541), .A2(KEYINPUT80), .A3(new_n543), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n550), .B1(new_n559), .B2(new_n282), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n536), .B(new_n549), .C1(new_n560), .C2(G169), .ZN(new_n561));
  INV_X1    g0361(.A(G303), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n339), .A2(new_n562), .A3(new_n340), .ZN(new_n563));
  NAND2_X1  g0363(.A1(G264), .A2(G1698), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n225), .B2(G1698), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n563), .B(new_n282), .C1(new_n353), .C2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n477), .A2(G270), .A3(new_n297), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n566), .A2(new_n480), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(KEYINPUT21), .A3(G169), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n566), .A2(new_n567), .A3(G179), .A4(new_n480), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n269), .A2(new_n212), .A3(G13), .A4(G20), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n268), .A2(G116), .A3(new_n274), .A4(new_n464), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n266), .A2(new_n233), .B1(G20), .B2(new_n212), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n504), .B(new_n234), .C1(G33), .C2(new_n224), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n574), .A2(KEYINPUT20), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT20), .B1(new_n574), .B2(new_n575), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n572), .B(new_n573), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n571), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT82), .ZN(new_n580));
  INV_X1    g0380(.A(new_n578), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n570), .B2(new_n569), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT82), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n578), .A2(G169), .A3(new_n568), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT21), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT83), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n585), .A2(KEYINPUT83), .A3(new_n586), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n580), .A2(new_n584), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n546), .A2(G190), .A3(new_n548), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n465), .A2(new_n217), .ZN(new_n593));
  AOI211_X1 g0393(.A(new_n523), .B(new_n593), .C1(new_n534), .C2(new_n267), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n592), .B(new_n594), .C1(new_n560), .C2(new_n378), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n568), .A2(G200), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n581), .B(new_n596), .C1(new_n329), .C2(new_n568), .ZN(new_n597));
  AND4_X1   g0397(.A1(new_n561), .A2(new_n591), .A3(new_n595), .A4(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n461), .A2(new_n487), .A3(new_n463), .A4(new_n467), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n481), .A2(new_n291), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n483), .A2(new_n335), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  AND4_X1   g0402(.A1(new_n445), .A2(new_n522), .A3(new_n598), .A4(new_n602), .ZN(G372));
  XNOR2_X1  g0403(.A(new_n391), .B(KEYINPUT18), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n336), .A2(new_n328), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n331), .A2(new_n313), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n606), .B1(new_n607), .B2(new_n293), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n385), .A2(KEYINPUT17), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n383), .A2(KEYINPUT75), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n383), .A2(KEYINPUT75), .A3(KEYINPUT17), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n604), .B1(new_n608), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n438), .A2(new_n439), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n414), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n445), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n513), .A2(new_n335), .A3(new_n515), .ZN(new_n619));
  AOI21_X1  g0419(.A(G169), .B1(new_n513), .B2(new_n515), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n619), .A2(new_n620), .A3(new_n497), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n582), .B1(new_n589), .B2(new_n590), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n602), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n621), .B1(new_n623), .B2(new_n488), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n534), .A2(new_n267), .ZN(new_n625));
  INV_X1    g0425(.A(new_n523), .ZN(new_n626));
  INV_X1    g0426(.A(new_n593), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(new_n560), .B2(G190), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n546), .A2(KEYINPUT86), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT86), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n631), .B(new_n282), .C1(new_n544), .C2(new_n545), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n550), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n629), .B1(new_n633), .B2(new_n378), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT26), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(new_n635), .A3(new_n521), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n624), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n621), .A2(new_n561), .A3(new_n595), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT26), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n536), .A2(new_n549), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n631), .B1(new_n559), .B2(new_n282), .ZN(new_n641));
  INV_X1    g0441(.A(new_n632), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n548), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n640), .B1(new_n643), .B2(new_n291), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n637), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n617), .B1(new_n618), .B2(new_n647), .ZN(new_n648));
  XOR2_X1   g0448(.A(new_n648), .B(KEYINPUT87), .Z(G369));
  INV_X1    g0449(.A(new_n622), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n269), .A2(new_n234), .A3(G13), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(G213), .A3(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(G343), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n581), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n650), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n591), .A2(new_n597), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n658), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(G330), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n599), .A2(new_n656), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n488), .A2(new_n602), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n602), .B2(new_n657), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n665), .A2(new_n591), .A3(new_n656), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n669));
  XOR2_X1   g0469(.A(new_n656), .B(KEYINPUT88), .Z(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n668), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n667), .A2(new_n672), .ZN(G399));
  NOR2_X1   g0473(.A1(new_n527), .A2(G116), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT89), .ZN(new_n675));
  INV_X1    g0475(.A(new_n208), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(G41), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n675), .A2(new_n677), .A3(new_n269), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n678), .B1(new_n239), .B2(new_n677), .ZN(new_n679));
  XOR2_X1   g0479(.A(new_n679), .B(KEYINPUT28), .Z(new_n680));
  INV_X1    g0480(.A(KEYINPUT29), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n634), .A2(new_n621), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n644), .B1(new_n682), .B2(KEYINPUT26), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n638), .A2(KEYINPUT26), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT92), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n571), .A2(new_n583), .A3(new_n578), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n583), .B1(new_n571), .B2(new_n578), .ZN(new_n687));
  INV_X1    g0487(.A(new_n590), .ZN(new_n688));
  AOI21_X1  g0488(.A(KEYINPUT83), .B1(new_n585), .B2(new_n586), .ZN(new_n689));
  OAI22_X1  g0489(.A1(new_n686), .A2(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n685), .B1(new_n669), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n645), .A2(new_n691), .A3(new_n634), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n591), .A2(KEYINPUT92), .A3(new_n602), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n693), .A2(new_n518), .A3(new_n521), .A4(new_n488), .ZN(new_n694));
  OAI211_X1 g0494(.A(new_n683), .B(new_n684), .C1(new_n692), .C2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n681), .B1(new_n695), .B2(new_n657), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n647), .A2(KEYINPUT29), .A3(new_n670), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n479), .B1(KEYINPUT90), .B2(new_n570), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n570), .A2(KEYINPUT90), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n520), .A2(new_n560), .A3(new_n700), .A4(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT30), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n546), .A2(new_n548), .A3(new_n701), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n516), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT30), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(new_n706), .A3(new_n700), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n481), .A2(new_n568), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n643), .A2(new_n335), .A3(new_n516), .A4(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n657), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(KEYINPUT91), .B1(new_n711), .B2(KEYINPUT31), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n706), .B1(new_n705), .B2(new_n700), .ZN(new_n713));
  NOR4_X1   g0513(.A1(new_n704), .A2(new_n516), .A3(KEYINPUT30), .A4(new_n699), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n710), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n656), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT91), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT31), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n715), .A2(KEYINPUT31), .A3(new_n670), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n598), .A2(new_n522), .A3(new_n602), .A4(new_n671), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n712), .A2(new_n719), .A3(new_n720), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G330), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n698), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n680), .B1(new_n725), .B2(G1), .ZN(G364));
  OR2_X1    g0526(.A1(new_n661), .A2(G330), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n206), .A2(G20), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n269), .B1(new_n728), .B2(G45), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n677), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n727), .A2(new_n662), .A3(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n676), .A2(new_n353), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G355), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n251), .A2(new_n473), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n676), .A2(new_n279), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(G45), .B2(new_n238), .ZN(new_n738));
  OAI221_X1 g0538(.A(new_n735), .B1(G116), .B2(new_n208), .C1(new_n736), .C2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G13), .A2(G33), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n234), .ZN(new_n741));
  XOR2_X1   g0541(.A(new_n741), .B(KEYINPUT93), .Z(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n233), .B1(G20), .B2(new_n291), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n739), .A2(new_n745), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n731), .B(new_n746), .C1(new_n661), .C2(new_n742), .ZN(new_n747));
  INV_X1    g0547(.A(new_n744), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n335), .A2(new_n378), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n234), .A2(G190), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  XNOR2_X1  g0552(.A(KEYINPUT33), .B(G317), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n378), .A2(G179), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n750), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n752), .A2(new_n753), .B1(new_n756), .B2(G283), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n234), .A2(new_n329), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(new_n749), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G326), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G179), .A2(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n750), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G329), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n757), .A2(new_n761), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n335), .A2(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n758), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n769), .A2(G322), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n758), .A2(new_n754), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n562), .ZN(new_n772));
  NOR4_X1   g0572(.A1(new_n766), .A2(new_n279), .A3(new_n770), .A4(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n234), .B1(new_n762), .B2(G190), .ZN(new_n774));
  INV_X1    g0574(.A(G311), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n750), .A2(new_n767), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n773), .B1(new_n471), .B2(new_n774), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT94), .Z(new_n778));
  NAND2_X1  g0578(.A1(new_n764), .A2(G159), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT32), .ZN(new_n780));
  INV_X1    g0580(.A(new_n776), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n353), .B(new_n780), .C1(G77), .C2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n756), .A2(G107), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n774), .A2(new_n224), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n222), .A2(new_n768), .B1(new_n751), .B2(new_n215), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n784), .B(new_n785), .C1(G50), .C2(new_n760), .ZN(new_n786));
  INV_X1    g0586(.A(new_n771), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G87), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n782), .A2(new_n783), .A3(new_n786), .A4(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n748), .B1(new_n778), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n733), .B1(new_n747), .B2(new_n790), .ZN(G396));
  NAND2_X1  g0591(.A1(new_n293), .A2(new_n657), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n278), .A2(new_n292), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n657), .B1(new_n273), .B2(new_n277), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n793), .B1(new_n443), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(new_n647), .B2(new_n670), .ZN(new_n797));
  INV_X1    g0597(.A(new_n796), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n671), .B(new_n798), .C1(new_n637), .C2(new_n646), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(new_n723), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(new_n732), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G143), .A2(new_n769), .B1(new_n781), .B2(G159), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n760), .A2(G137), .ZN(new_n804));
  INV_X1    g0604(.A(G150), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n803), .B(new_n804), .C1(new_n805), .C2(new_n751), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT34), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n279), .B1(new_n774), .B2(new_n222), .ZN(new_n808));
  INV_X1    g0608(.A(G132), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n755), .A2(new_n215), .B1(new_n763), .B2(new_n809), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n808), .B(new_n810), .C1(G50), .C2(new_n787), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n784), .B1(G294), .B2(new_n769), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT95), .Z(new_n814));
  AOI211_X1 g0614(.A(new_n279), .B(new_n814), .C1(G303), .C2(new_n760), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n787), .A2(G107), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n752), .A2(G283), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G116), .A2(new_n781), .B1(new_n764), .B2(G311), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n815), .A2(new_n816), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n755), .A2(new_n217), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n812), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n732), .B1(new_n821), .B2(new_n744), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n744), .A2(new_n740), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n740), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n822), .B1(G77), .B2(new_n824), .C1(new_n825), .C2(new_n798), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n802), .A2(new_n826), .ZN(G384));
  NAND3_X1  g0627(.A1(new_n715), .A2(KEYINPUT31), .A3(new_n656), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n721), .B(new_n828), .C1(KEYINPUT31), .C2(new_n711), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n606), .A2(new_n656), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n328), .A2(new_n656), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n605), .A2(new_n607), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n796), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  AND3_X1   g0633(.A1(new_n829), .A2(new_n833), .A3(KEYINPUT40), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n654), .B1(new_n359), .B2(new_n369), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n394), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT37), .ZN(new_n837));
  AND3_X1   g0637(.A1(new_n359), .A2(new_n369), .A3(new_n382), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n838), .A2(new_n391), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n359), .A2(new_n369), .ZN(new_n840));
  INV_X1    g0640(.A(new_n654), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n837), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n390), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n654), .B(KEYINPUT98), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n840), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n359), .A2(new_n369), .A3(new_n382), .ZN(new_n848));
  AND4_X1   g0648(.A1(new_n837), .A2(new_n845), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(KEYINPUT99), .B1(new_n843), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT99), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n845), .A2(new_n847), .A3(new_n837), .A4(new_n848), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n838), .A2(new_n391), .A3(new_n835), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n851), .B(new_n852), .C1(new_n853), .C2(new_n837), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n836), .A2(new_n850), .A3(KEYINPUT38), .A4(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT38), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n847), .B1(new_n613), .B2(new_n604), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n837), .B1(new_n839), .B2(new_n847), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n858), .A2(new_n849), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n856), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n855), .A2(new_n860), .A3(KEYINPUT100), .ZN(new_n861));
  INV_X1    g0661(.A(new_n854), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n845), .A2(new_n842), .A3(new_n848), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT37), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n851), .B1(new_n864), .B2(new_n852), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT100), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n866), .A2(new_n867), .A3(KEYINPUT38), .A4(new_n836), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n861), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n834), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT40), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n836), .A2(new_n850), .A3(new_n854), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n856), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n873), .A2(new_n855), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n829), .A2(new_n833), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n871), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n870), .A2(new_n876), .A3(G330), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n445), .A2(G330), .A3(new_n829), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n873), .A2(new_n855), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n880), .A2(new_n833), .A3(new_n829), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n869), .A2(new_n834), .B1(new_n881), .B2(new_n871), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n882), .A2(new_n445), .A3(new_n829), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n604), .A2(new_n846), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n336), .A2(new_n328), .B1(new_n313), .B2(new_n331), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n606), .A2(new_n656), .B1(new_n886), .B2(new_n831), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n799), .B2(new_n792), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n885), .B1(new_n888), .B2(new_n880), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT39), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n861), .A2(new_n868), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n606), .A2(new_n657), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n873), .A2(KEYINPUT39), .A3(new_n855), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n889), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n884), .B(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n617), .B1(new_n698), .B2(new_n618), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n897), .B(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n269), .B2(new_n728), .ZN(new_n900));
  OAI21_X1  g0700(.A(G77), .B1(new_n222), .B2(new_n215), .ZN(new_n901));
  OAI22_X1  g0701(.A1(new_n238), .A2(new_n901), .B1(G50), .B2(new_n215), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n902), .A2(G1), .A3(new_n206), .ZN(new_n903));
  OAI211_X1 g0703(.A(G116), .B(new_n235), .C1(new_n491), .C2(KEYINPUT35), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT96), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n491), .A2(KEYINPUT35), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XOR2_X1   g0707(.A(KEYINPUT97), .B(KEYINPUT36), .Z(new_n908));
  XNOR2_X1  g0708(.A(new_n907), .B(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n900), .A2(new_n903), .A3(new_n909), .ZN(G367));
  INV_X1    g0710(.A(new_n667), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n518), .B(new_n521), .C1(new_n497), .C2(new_n671), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT103), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n518), .B2(new_n671), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n668), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT42), .Z(new_n916));
  OAI21_X1  g0716(.A(new_n518), .B1(new_n913), .B2(new_n602), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n671), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n645), .B(new_n634), .C1(new_n594), .C2(new_n657), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n594), .A2(new_n657), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n920), .A2(KEYINPUT101), .B1(new_n644), .B2(new_n921), .ZN(new_n922));
  AND3_X1   g0722(.A1(new_n644), .A2(KEYINPUT101), .A3(new_n921), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n924), .B(KEYINPUT102), .Z(new_n925));
  INV_X1    g0725(.A(KEYINPUT43), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n919), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n919), .B(new_n927), .C1(new_n926), .C2(new_n924), .ZN(new_n929));
  AND4_X1   g0729(.A1(new_n911), .A2(new_n928), .A3(new_n929), .A4(new_n914), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n928), .A2(new_n929), .B1(new_n911), .B2(new_n914), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n914), .A2(new_n672), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n933), .B(KEYINPUT44), .Z(new_n934));
  NAND2_X1  g0734(.A1(new_n914), .A2(new_n672), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT45), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n666), .B1(new_n690), .B2(new_n657), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n662), .B1(new_n938), .B2(new_n668), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n667), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n725), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n937), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n725), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n677), .B(KEYINPUT41), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n729), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n932), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(KEYINPUT104), .B(G137), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n279), .B1(new_n763), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(G143), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n759), .A2(new_n952), .B1(new_n768), .B2(new_n805), .ZN(new_n953));
  INV_X1    g0753(.A(new_n774), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n953), .B1(G68), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n756), .A2(G77), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n787), .A2(G58), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n781), .A2(G50), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n955), .A2(new_n956), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n951), .B(new_n959), .C1(G159), .C2(new_n752), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT105), .Z(new_n961));
  NAND2_X1  g0761(.A1(new_n756), .A2(G97), .ZN(new_n962));
  INV_X1    g0762(.A(G283), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n962), .B1(new_n963), .B2(new_n776), .C1(new_n471), .C2(new_n751), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(G317), .B2(new_n764), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n353), .B1(new_n774), .B2(new_n449), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(G303), .B2(new_n769), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n965), .B(new_n967), .C1(new_n775), .C2(new_n759), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n771), .A2(new_n212), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT46), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n961), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT47), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n744), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n924), .A2(new_n743), .ZN(new_n974));
  INV_X1    g0774(.A(new_n737), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n745), .B1(new_n208), .B2(new_n264), .C1(new_n247), .C2(new_n975), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n973), .A2(new_n974), .A3(new_n731), .A4(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT106), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n949), .A2(new_n979), .ZN(G387));
  AOI22_X1  g0780(.A1(G322), .A2(new_n760), .B1(new_n752), .B2(G311), .ZN(new_n981));
  INV_X1    g0781(.A(G317), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n981), .B1(new_n562), .B2(new_n776), .C1(new_n982), .C2(new_n768), .ZN(new_n983));
  XOR2_X1   g0783(.A(KEYINPUT108), .B(KEYINPUT48), .Z(new_n984));
  XNOR2_X1  g0784(.A(new_n983), .B(new_n984), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n963), .B2(new_n774), .C1(new_n471), .C2(new_n771), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT49), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n756), .A2(G116), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n764), .A2(G326), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n988), .A2(new_n353), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n986), .A2(new_n987), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n367), .A2(new_n751), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n264), .A2(new_n774), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n279), .B1(new_n776), .B2(new_n215), .C1(new_n227), .C2(new_n768), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(G159), .C2(new_n760), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n771), .A2(new_n259), .B1(new_n763), .B2(new_n805), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT107), .Z(new_n998));
  NAND3_X1  g0798(.A1(new_n996), .A2(new_n962), .A3(new_n998), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n991), .A2(new_n992), .B1(new_n993), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n744), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n975), .B1(new_n244), .B2(G45), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n675), .B2(new_n734), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n256), .A2(G50), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT50), .Z(new_n1005));
  NOR2_X1   g0805(.A1(new_n215), .A2(new_n259), .ZN(new_n1006));
  NOR4_X1   g0806(.A1(new_n1005), .A2(G45), .A3(new_n675), .A4(new_n1006), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n1003), .A2(new_n1007), .B1(G107), .B2(new_n208), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n732), .B1(new_n1008), .B2(new_n745), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1001), .B(new_n1009), .C1(new_n666), .C2(new_n742), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n677), .B1(new_n725), .B2(new_n941), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1010), .B1(new_n729), .B2(new_n940), .C1(new_n943), .C2(new_n1011), .ZN(G393));
  OR4_X1    g0812(.A1(KEYINPUT109), .A2(new_n934), .A3(new_n667), .A4(new_n936), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n667), .A2(KEYINPUT109), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n667), .A2(KEYINPUT109), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n937), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n677), .B(new_n944), .C1(new_n1017), .C2(new_n943), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n914), .A2(new_n742), .ZN(new_n1019));
  INV_X1    g0819(.A(G159), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n759), .A2(new_n805), .B1(new_n768), .B2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT51), .Z(new_n1022));
  OAI21_X1  g0822(.A(new_n279), .B1(new_n755), .B2(new_n217), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n771), .A2(new_n215), .B1(new_n776), .B2(new_n256), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n751), .A2(new_n227), .ZN(new_n1025));
  NOR4_X1   g0825(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n259), .B2(new_n774), .C1(new_n952), .C2(new_n763), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n783), .B1(new_n963), .B2(new_n771), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n759), .A2(new_n982), .B1(new_n768), .B2(new_n775), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1029), .B(new_n1030), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n1028), .B(new_n1031), .C1(G294), .C2(new_n781), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n764), .A2(G322), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n954), .A2(G116), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n279), .B1(new_n752), .B2(G303), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n748), .B1(new_n1027), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n745), .B1(new_n254), .B2(new_n975), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(G97), .B2(new_n676), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n1037), .A2(new_n732), .A3(new_n1039), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n1017), .A2(new_n730), .B1(new_n1019), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1018), .A2(new_n1041), .ZN(G390));
  AND3_X1   g0842(.A1(new_n861), .A2(new_n868), .A3(new_n890), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n894), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n740), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n788), .A2(new_n353), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT116), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n755), .A2(new_n215), .B1(new_n774), .B2(new_n259), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n751), .A2(new_n449), .B1(new_n776), .B2(new_n224), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n759), .A2(new_n963), .ZN(new_n1050));
  NOR4_X1   g0850(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n212), .B2(new_n768), .C1(new_n471), .C2(new_n763), .ZN(new_n1052));
  OAI21_X1  g0852(.A(KEYINPUT53), .B1(new_n771), .B2(new_n805), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n1020), .B2(new_n774), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n279), .B1(new_n755), .B2(new_n227), .C1(new_n751), .C2(new_n950), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n771), .A2(KEYINPUT53), .A3(new_n805), .ZN(new_n1056));
  NOR3_X1   g0856(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n760), .A2(G128), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n764), .A2(G125), .ZN(new_n1059));
  XOR2_X1   g0859(.A(KEYINPUT54), .B(G143), .Z(new_n1060));
  AOI22_X1  g0860(.A1(G132), .A2(new_n769), .B1(new_n781), .B2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .A4(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n748), .B1(new_n1052), .B2(new_n1062), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n732), .B(new_n1063), .C1(new_n367), .C2(new_n823), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n1045), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n861), .A2(new_n868), .A3(new_n892), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n695), .A2(new_n657), .A3(new_n795), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1068), .A2(new_n792), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1067), .B1(new_n1069), .B2(new_n887), .ZN(new_n1070));
  INV_X1    g0870(.A(G330), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n717), .B1(new_n716), .B2(new_n718), .ZN(new_n1072));
  AOI211_X1 g0872(.A(KEYINPUT91), .B(KEYINPUT31), .C1(new_n715), .C2(new_n656), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n721), .A2(new_n720), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1071), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n887), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT111), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n829), .A2(new_n833), .A3(new_n1078), .A4(G330), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1076), .A2(new_n798), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n1043), .A2(new_n1044), .B1(new_n893), .B2(new_n888), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1070), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n829), .A2(new_n833), .A3(G330), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1083), .A2(KEYINPUT111), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n799), .A2(new_n792), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n1077), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1086), .A2(new_n892), .B1(new_n891), .B2(new_n894), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1068), .A2(new_n792), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1066), .B1(new_n1088), .B2(new_n1077), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1084), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1082), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(KEYINPUT115), .B1(new_n1091), .B2(new_n729), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT115), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1082), .A2(new_n1090), .A3(new_n1093), .A4(new_n730), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1091), .A2(KEYINPUT113), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT113), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1082), .A2(new_n1090), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT112), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n878), .B(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1099), .A2(new_n898), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT114), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n722), .A2(G330), .A3(new_n798), .A4(new_n1077), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n829), .A2(G330), .A3(new_n798), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n887), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1102), .A2(new_n1069), .A3(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n722), .A2(G330), .A3(new_n798), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1083), .B1(new_n1106), .B2(new_n887), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1085), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1105), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n1100), .A2(new_n1101), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1101), .B1(new_n1100), .B2(new_n1109), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1095), .B(new_n1097), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1100), .A2(new_n1109), .A3(new_n1082), .A4(new_n1090), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1113), .A2(new_n677), .ZN(new_n1114));
  AOI221_X4 g0914(.A(new_n1065), .B1(new_n1092), .B2(new_n1094), .C1(new_n1112), .C2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(G378));
  INV_X1    g0916(.A(KEYINPUT120), .ZN(new_n1117));
  XOR2_X1   g0917(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1118));
  XNOR2_X1  g0918(.A(new_n440), .B(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n412), .A2(new_n841), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT118), .Z(new_n1121));
  AND2_X1   g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT119), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1124), .B1(new_n877), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n889), .A2(new_n895), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n882), .A2(new_n1127), .A3(KEYINPUT119), .A4(G330), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n870), .A2(new_n876), .A3(KEYINPUT119), .A4(G330), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n896), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n1126), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n877), .A2(new_n1125), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1124), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1128), .A2(new_n1130), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1117), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1126), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1126), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1138), .A2(KEYINPUT120), .A3(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1135), .A2(new_n1140), .A3(new_n730), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n731), .B1(G50), .B2(new_n824), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n227), .B1(new_n351), .B2(G41), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n259), .A2(new_n771), .B1(new_n768), .B2(new_n449), .ZN(new_n1144));
  AOI211_X1 g0944(.A(G41), .B(new_n1144), .C1(G68), .C2(new_n954), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n279), .B1(new_n756), .B2(G58), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n781), .A2(new_n263), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(G97), .A2(new_n752), .B1(new_n764), .B2(G283), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G116), .B2(new_n760), .ZN(new_n1150));
  XOR2_X1   g0950(.A(new_n1150), .B(KEYINPUT58), .Z(new_n1151));
  OAI22_X1  g0951(.A1(new_n751), .A2(new_n809), .B1(new_n774), .B2(new_n805), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n787), .A2(new_n1060), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT117), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1153), .A2(new_n1154), .B1(new_n760), .B2(G125), .ZN(new_n1155));
  INV_X1    g0955(.A(G128), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1155), .B1(new_n1156), .B2(new_n768), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1152), .B(new_n1157), .C1(G137), .C2(new_n781), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n1154), .B2(new_n1153), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1159), .A2(KEYINPUT59), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(KEYINPUT59), .ZN(new_n1161));
  AOI21_X1  g0961(.A(G33), .B1(new_n764), .B2(G124), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1160), .A2(new_n296), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n755), .A2(new_n1020), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1143), .B(new_n1151), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1142), .B1(new_n1165), .B2(new_n744), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n1133), .B2(new_n825), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1141), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1131), .A2(new_n1134), .A3(new_n1117), .ZN(new_n1170));
  AOI21_X1  g0970(.A(KEYINPUT120), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1113), .A2(new_n1100), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT121), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1109), .ZN(new_n1176));
  OAI211_X1 g0976(.A(KEYINPUT121), .B(new_n1100), .C1(new_n1091), .C2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT57), .B1(new_n1172), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1177), .ZN(new_n1180));
  AOI21_X1  g0980(.A(KEYINPUT121), .B1(new_n1113), .B2(new_n1100), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1138), .A2(KEYINPUT57), .A3(new_n1139), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n677), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1169), .B1(new_n1179), .B2(new_n1184), .ZN(G375));
  OR2_X1    g0985(.A1(new_n1100), .A2(new_n1109), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n946), .B(new_n1186), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT122), .Z(new_n1188));
  NAND2_X1  g0988(.A1(new_n887), .A2(new_n740), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(G116), .A2(new_n752), .B1(new_n781), .B2(G107), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n279), .B(new_n994), .C1(new_n1190), .C2(KEYINPUT123), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1190), .A2(KEYINPUT123), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n760), .A2(G294), .B1(new_n764), .B2(G303), .ZN(new_n1193));
  AND4_X1   g0993(.A1(new_n956), .A2(new_n1191), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1194), .B1(new_n224), .B2(new_n771), .C1(new_n963), .C2(new_n768), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G159), .A2(new_n787), .B1(new_n756), .B2(G58), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1196), .B1(new_n227), .B2(new_n774), .C1(new_n768), .C2(new_n950), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n279), .B1(new_n776), .B2(new_n805), .C1(new_n809), .C2(new_n759), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n752), .A2(new_n1060), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(new_n1156), .C2(new_n763), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n748), .B1(new_n1195), .B2(new_n1201), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n732), .B(new_n1202), .C1(new_n215), .C2(new_n823), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1109), .A2(new_n730), .B1(new_n1189), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1188), .A2(new_n1204), .ZN(G381));
  INV_X1    g1005(.A(KEYINPUT57), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1135), .A2(new_n1140), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1206), .B1(new_n1207), .B2(new_n1182), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n677), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1183), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1209), .B1(new_n1178), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1168), .B1(new_n1208), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n1115), .ZN(new_n1213));
  NOR4_X1   g1013(.A1(new_n1213), .A2(G384), .A3(G381), .A4(G387), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(G390), .A2(G396), .A3(G393), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(G407));
  OAI211_X1 g1016(.A(G407), .B(G213), .C1(G343), .C2(new_n1213), .ZN(G409));
  NAND2_X1  g1017(.A1(new_n655), .A2(G213), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1178), .A2(new_n946), .A3(new_n1140), .A4(new_n1135), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1138), .A2(new_n730), .A3(new_n1139), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1115), .A2(new_n1219), .A3(new_n1167), .A4(new_n1220), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1218), .B(new_n1221), .C1(new_n1212), .C2(new_n1115), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT62), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT60), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1186), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1100), .A2(new_n1109), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1186), .A2(new_n1225), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1226), .A2(new_n677), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n1204), .ZN(new_n1230));
  INV_X1    g1030(.A(G384), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1229), .A2(G384), .A3(new_n1204), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1223), .A2(new_n1224), .A3(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(G390), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(G387), .A2(new_n1237), .ZN(new_n1238));
  XOR2_X1   g1038(.A(G393), .B(G396), .Z(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(KEYINPUT127), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1240), .B1(G387), .B2(new_n1237), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n949), .A2(new_n1239), .A3(G390), .A4(new_n979), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1241), .B1(new_n1244), .B2(new_n1238), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT61), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n655), .A2(G213), .A3(G2897), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1234), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1247), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1232), .A2(new_n1233), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1222), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1236), .A2(new_n1245), .A3(new_n1246), .A4(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1224), .B1(new_n1223), .B2(new_n1235), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT124), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n1222), .B2(new_n1234), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT63), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1256), .B(KEYINPUT63), .C1(new_n1222), .C2(new_n1234), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G375), .A2(G378), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT125), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1262), .A2(new_n1263), .A3(new_n1218), .A4(new_n1221), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1222), .A2(KEYINPUT125), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1264), .A2(new_n1265), .A3(new_n1251), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(KEYINPUT126), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT126), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1264), .A2(new_n1265), .A3(new_n1268), .A4(new_n1251), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1261), .A2(new_n1267), .A3(new_n1246), .A4(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1245), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1255), .B1(new_n1270), .B2(new_n1271), .ZN(G405));
  NAND2_X1  g1072(.A1(new_n1262), .A2(new_n1213), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1273), .B(new_n1235), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1274), .B(new_n1271), .ZN(G402));
endmodule


