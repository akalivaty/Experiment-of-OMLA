//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 0 0 0 0 0 1 0 1 1 0 1 1 0 1 1 0 1 0 0 1 1 1 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 1 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n805, new_n806, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G43gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G71gat), .B(G99gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  NAND2_X1  g004(.A1(G227gat), .A2(G233gat), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n206), .B(KEYINPUT64), .Z(new_n207));
  INV_X1    g006(.A(G183gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT27), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT68), .ZN(new_n210));
  AOI21_X1  g009(.A(G190gat), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT27), .B(G183gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n211), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT69), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n211), .B(KEYINPUT69), .C1(new_n210), .C2(new_n212), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT28), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G190gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n212), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT28), .ZN(new_n220));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n223), .A2(KEYINPUT26), .ZN(new_n224));
  NAND2_X1  g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT26), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n225), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n220), .B(new_n221), .C1(new_n224), .C2(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n217), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n222), .A2(KEYINPUT23), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(new_n225), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT67), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT25), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT67), .B1(new_n230), .B2(new_n225), .ZN(new_n235));
  NOR3_X1   g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  XOR2_X1   g035(.A(KEYINPUT66), .B(KEYINPUT23), .Z(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(new_n223), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT24), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n221), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n240), .B(new_n241), .C1(G183gat), .C2(G190gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n238), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT65), .B(G176gat), .ZN(new_n245));
  INV_X1    g044(.A(G169gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT23), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n248), .A2(new_n238), .A3(new_n242), .A4(new_n225), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n236), .A2(new_n244), .B1(new_n249), .B2(new_n234), .ZN(new_n250));
  INV_X1    g049(.A(G113gat), .ZN(new_n251));
  INV_X1    g050(.A(G120gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT1), .ZN(new_n254));
  NAND2_X1  g053(.A1(G113gat), .A2(G120gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G134gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G127gat), .ZN(new_n258));
  INV_X1    g057(.A(G127gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G134gat), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT70), .B1(new_n257), .B2(G127gat), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n256), .A2(new_n258), .A3(new_n260), .A4(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n254), .B1(G113gat), .B2(G120gat), .ZN(new_n263));
  INV_X1    g062(.A(new_n255), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n258), .A2(new_n260), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n262), .A2(new_n267), .A3(KEYINPUT71), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT71), .B1(new_n262), .B2(new_n267), .ZN(new_n270));
  OAI22_X1  g069(.A1(new_n229), .A2(new_n250), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n225), .B1(new_n245), .B2(new_n247), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n234), .B1(new_n243), .B2(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n235), .A2(new_n234), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n274), .B1(new_n232), .B2(new_n231), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n275), .B2(new_n243), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n269), .A2(new_n270), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n276), .B(new_n277), .C1(new_n217), .C2(new_n228), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n207), .B1(new_n271), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n205), .B1(new_n279), .B2(KEYINPUT33), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT32), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n280), .B(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n271), .A2(new_n278), .ZN(new_n284));
  INV_X1    g083(.A(new_n206), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT34), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT34), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n271), .A2(new_n278), .A3(new_n287), .A4(new_n207), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n283), .B(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT86), .ZN(new_n291));
  NAND2_X1  g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT75), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT75), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n294), .A2(G155gat), .A3(G162gat), .ZN(new_n295));
  INV_X1    g094(.A(G155gat), .ZN(new_n296));
  INV_X1    g095(.A(G162gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n293), .A2(new_n295), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n294), .A2(KEYINPUT2), .ZN(new_n300));
  INV_X1    g099(.A(G148gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(G141gat), .ZN(new_n302));
  INV_X1    g101(.A(G141gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n303), .A2(G148gat), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n300), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT76), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(new_n301), .B2(G141gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n303), .A2(KEYINPUT76), .A3(G148gat), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n307), .B(new_n308), .C1(new_n303), .C2(G148gat), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n292), .B1(new_n298), .B2(KEYINPUT2), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n299), .A2(new_n305), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT79), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT79), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n311), .A2(new_n315), .A3(new_n312), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT29), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G197gat), .B(G204gat), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n319), .A2(KEYINPUT73), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(KEYINPUT73), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n318), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  XOR2_X1   g121(.A(G211gat), .B(G218gat), .Z(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n323), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n325), .B(new_n318), .C1(new_n320), .C2(new_n321), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n291), .B1(new_n317), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT29), .ZN(new_n329));
  INV_X1    g128(.A(new_n316), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n315), .B1(new_n311), .B2(new_n312), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n327), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(KEYINPUT86), .A3(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n327), .A2(KEYINPUT85), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT85), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n329), .B1(new_n326), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n312), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n299), .A2(new_n305), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n309), .A2(new_n310), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n328), .A2(new_n334), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(G228gat), .ZN(new_n344));
  INV_X1    g143(.A(G233gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(G22gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n332), .A2(KEYINPUT87), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT87), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n317), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n350), .A2(new_n352), .A3(new_n333), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(new_n333), .B2(KEYINPUT29), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n347), .B1(new_n355), .B2(new_n341), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n348), .A2(new_n349), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT89), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n343), .A2(new_n347), .B1(new_n353), .B2(new_n356), .ZN(new_n360));
  OAI21_X1  g159(.A(G22gat), .B1(new_n360), .B2(KEYINPUT88), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n348), .A2(KEYINPUT88), .A3(new_n357), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n359), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT88), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n343), .A2(new_n347), .ZN(new_n365));
  INV_X1    g164(.A(new_n357), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n360), .A2(KEYINPUT88), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n367), .A2(KEYINPUT89), .A3(new_n368), .A4(G22gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(G78gat), .B(G106gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT31), .B(G50gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n363), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(G22gat), .B1(new_n365), .B2(new_n366), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n372), .B1(new_n374), .B2(new_n358), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n290), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT93), .ZN(new_n378));
  XNOR2_X1  g177(.A(G8gat), .B(G36gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(G64gat), .B(G92gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(G226gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n382), .A2(new_n345), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n383), .A2(KEYINPUT29), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT74), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n276), .B(new_n386), .C1(new_n217), .C2(new_n228), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT74), .B1(new_n229), .B2(new_n250), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n385), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NOR4_X1   g188(.A1(new_n229), .A2(new_n250), .A3(new_n382), .A4(new_n345), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n389), .A2(new_n327), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n387), .A2(new_n388), .A3(new_n383), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n384), .B1(new_n229), .B2(new_n250), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n333), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n381), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n392), .A2(new_n393), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n327), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n387), .A2(new_n388), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(new_n384), .ZN(new_n399));
  INV_X1    g198(.A(new_n390), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(new_n333), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n381), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n397), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n395), .A2(new_n403), .A3(KEYINPUT30), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n391), .A2(new_n394), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT30), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(new_n406), .A3(new_n402), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n262), .A2(new_n267), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n311), .A2(new_n409), .ZN(new_n410));
  OR3_X1    g209(.A1(new_n410), .A2(KEYINPUT80), .A3(KEYINPUT4), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT80), .B1(new_n410), .B2(KEYINPUT4), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT4), .ZN(new_n413));
  NOR3_X1   g212(.A1(new_n269), .A2(new_n341), .A3(new_n270), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n411), .B(new_n412), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(G225gat), .A2(G233gat), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n314), .A2(new_n316), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n341), .A2(KEYINPUT3), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT77), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n409), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n262), .A2(new_n267), .A3(KEYINPUT77), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n419), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n417), .B1(new_n418), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n415), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n421), .A2(new_n341), .A3(new_n422), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n416), .B1(new_n426), .B2(new_n410), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT5), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT81), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n427), .A2(KEYINPUT81), .A3(new_n428), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n425), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n410), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT82), .B1(new_n433), .B2(new_n413), .ZN(new_n434));
  INV_X1    g233(.A(new_n270), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n435), .A2(new_n413), .A3(new_n311), .A4(new_n268), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT82), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n410), .A2(new_n437), .A3(KEYINPUT4), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n434), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n418), .A2(new_n423), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n417), .A2(KEYINPUT5), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(G1gat), .B(G29gat), .ZN(new_n444));
  INV_X1    g243(.A(G85gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(KEYINPUT0), .B(G57gat), .ZN(new_n447));
  XOR2_X1   g246(.A(new_n446), .B(new_n447), .Z(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n432), .A2(new_n443), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n432), .A2(new_n443), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n449), .B1(new_n453), .B2(KEYINPUT90), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT90), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n432), .A2(new_n443), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n452), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n427), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT81), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(new_n459), .A3(KEYINPUT5), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n460), .A2(new_n429), .B1(new_n415), .B2(new_n424), .ZN(new_n461));
  OAI211_X1 g260(.A(KEYINPUT6), .B(new_n448), .C1(new_n461), .C2(new_n442), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT84), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT84), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n453), .A2(new_n464), .A3(KEYINPUT6), .A4(new_n448), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n378), .B(new_n408), .C1(new_n457), .C2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT90), .B1(new_n461), .B2(new_n442), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(new_n456), .A3(new_n448), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n461), .A2(new_n442), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT6), .B1(new_n471), .B2(new_n449), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n473), .A2(new_n465), .A3(new_n463), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n378), .B1(new_n474), .B2(new_n408), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n202), .B(new_n377), .C1(new_n468), .C2(new_n475), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n404), .A2(new_n407), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT83), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n452), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n453), .A2(new_n448), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n450), .A2(KEYINPUT83), .A3(new_n451), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n466), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n477), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n373), .A2(new_n376), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT72), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n283), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(new_n289), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n484), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT35), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n482), .A2(new_n483), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n408), .ZN(new_n492));
  INV_X1    g291(.A(new_n372), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n367), .A2(G22gat), .A3(new_n368), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n493), .B1(new_n494), .B2(new_n359), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n375), .B1(new_n495), .B2(new_n369), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT36), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n290), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n487), .A2(new_n286), .A3(new_n288), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n283), .A2(new_n486), .A3(new_n289), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(KEYINPUT36), .A3(new_n500), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n492), .A2(new_n496), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n439), .A2(new_n440), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n503), .A2(new_n416), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT39), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n448), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n426), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n507), .A2(new_n433), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n505), .B1(new_n508), .B2(new_n416), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n509), .B1(new_n503), .B2(new_n416), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT40), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n506), .A2(KEYINPUT40), .A3(new_n510), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n477), .A2(new_n470), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT92), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT37), .ZN(new_n517));
  OAI211_X1 g316(.A(KEYINPUT91), .B(new_n327), .C1(new_n389), .C2(new_n390), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n392), .A2(new_n333), .A3(new_n393), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT91), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n389), .A2(new_n390), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n521), .B1(new_n522), .B2(new_n333), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n517), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n397), .A2(new_n401), .A3(new_n517), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT38), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(new_n526), .A3(new_n381), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n516), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n399), .A2(new_n400), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT91), .B1(new_n529), .B2(new_n327), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n518), .A2(new_n519), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT37), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n402), .B1(new_n405), .B2(new_n517), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n532), .A2(new_n533), .A3(KEYINPUT92), .A4(new_n526), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n525), .A2(new_n381), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n405), .A2(new_n517), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT38), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n528), .A2(new_n534), .A3(new_n403), .A4(new_n537), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n485), .B(new_n515), .C1(new_n538), .C2(new_n474), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n476), .A2(new_n490), .B1(new_n502), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G231gat), .A2(G233gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(new_n208), .ZN(new_n542));
  INV_X1    g341(.A(G211gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(G71gat), .A2(G78gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT97), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(G71gat), .ZN(new_n551));
  INV_X1    g350(.A(G78gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(KEYINPUT97), .A2(G71gat), .A3(G78gat), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n550), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT98), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(G57gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(G64gat), .ZN(new_n559));
  INV_X1    g358(.A(G64gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(G57gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT9), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n550), .A2(new_n553), .A3(KEYINPUT98), .A4(new_n554), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n557), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n553), .A2(new_n548), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n562), .A2(new_n568), .A3(new_n564), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT99), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT99), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n562), .A2(new_n568), .A3(new_n571), .A4(new_n564), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n567), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(KEYINPUT100), .B(KEYINPUT21), .Z(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(new_n259), .ZN(new_n576));
  XNOR2_X1  g375(.A(G15gat), .B(G22gat), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT16), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n577), .B1(new_n578), .B2(G1gat), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n579), .B1(G1gat), .B2(new_n577), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(G8gat), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT21), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n582), .B1(new_n583), .B2(new_n573), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n576), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT103), .B(G155gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n576), .A2(new_n584), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n586), .B1(new_n585), .B2(new_n587), .ZN(new_n589));
  XNOR2_X1  g388(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n590));
  NOR3_X1   g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n590), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n576), .B(new_n584), .ZN(new_n593));
  INV_X1    g392(.A(new_n586), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n592), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n547), .B1(new_n591), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n590), .B1(new_n588), .B2(new_n589), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n595), .A2(new_n592), .A3(new_n596), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(new_n600), .A3(new_n546), .ZN(new_n601));
  XNOR2_X1  g400(.A(G190gat), .B(G218gat), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n602), .A2(KEYINPUT106), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT104), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n604), .A2(G92gat), .ZN(new_n605));
  INV_X1    g404(.A(G92gat), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n606), .A2(KEYINPUT104), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n445), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  AND2_X1   g407(.A1(G99gat), .A2(G106gat), .ZN(new_n609));
  NOR2_X1   g408(.A1(G99gat), .A2(G106gat), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT7), .ZN(new_n613));
  NAND2_X1  g412(.A1(G85gat), .A2(G92gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(G99gat), .A2(G106gat), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n613), .A2(new_n614), .B1(new_n615), .B2(KEYINPUT8), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n608), .A2(new_n611), .A3(new_n612), .A4(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n609), .A2(new_n610), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(KEYINPUT8), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n614), .A2(new_n613), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n619), .A2(new_n620), .A3(new_n612), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n606), .A2(KEYINPUT104), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n604), .A2(G92gat), .ZN(new_n623));
  AOI21_X1  g422(.A(G85gat), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n618), .B1(new_n621), .B2(new_n624), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n617), .A2(new_n625), .A3(KEYINPUT105), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT105), .B1(new_n617), .B2(new_n625), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(G29gat), .A2(G36gat), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT14), .ZN(new_n631));
  INV_X1    g430(.A(G29gat), .ZN(new_n632));
  INV_X1    g431(.A(G36gat), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n630), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AND2_X1   g435(.A1(G43gat), .A2(G50gat), .ZN(new_n637));
  NOR2_X1   g436(.A1(G43gat), .A2(G50gat), .ZN(new_n638));
  OAI21_X1  g437(.A(KEYINPUT15), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(G43gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(KEYINPUT94), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT94), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(G43gat), .ZN(new_n643));
  AOI21_X1  g442(.A(G50gat), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT15), .ZN(new_n645));
  INV_X1    g444(.A(G50gat), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n645), .B1(new_n640), .B2(new_n646), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n636), .B(new_n639), .C1(new_n644), .C2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n634), .A2(new_n635), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n629), .ZN(new_n650));
  INV_X1    g449(.A(new_n639), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(KEYINPUT95), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT17), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT95), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n648), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n654), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n656), .B1(new_n648), .B2(new_n652), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n649), .A2(new_n639), .A3(new_n629), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n641), .A2(new_n643), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n646), .ZN(new_n662));
  INV_X1    g461(.A(new_n647), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(KEYINPUT95), .B1(new_n660), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(KEYINPUT17), .B1(new_n659), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n628), .B1(new_n658), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT105), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n619), .A2(new_n620), .A3(new_n612), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n611), .B1(new_n670), .B2(new_n608), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n621), .A2(new_n624), .A3(new_n618), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n669), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n617), .A2(new_n625), .A3(KEYINPUT105), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n659), .A2(new_n665), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n668), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n603), .B1(new_n667), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n602), .A2(KEYINPUT106), .ZN(new_n679));
  AOI21_X1  g478(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(G134gat), .B(G162gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n678), .A2(new_n684), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n603), .B(new_n683), .C1(new_n667), .C2(new_n677), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n598), .A2(new_n601), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(G120gat), .B(G148gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(G176gat), .B(G204gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(G230gat), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n345), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n567), .A2(KEYINPUT10), .A3(new_n570), .A4(new_n572), .ZN(new_n694));
  OAI21_X1  g493(.A(KEYINPUT108), .B1(new_n675), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n694), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT108), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n696), .A2(new_n697), .A3(new_n674), .A4(new_n673), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n617), .A2(new_n625), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n573), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n573), .A2(new_n700), .ZN(new_n702));
  XOR2_X1   g501(.A(KEYINPUT107), .B(KEYINPUT10), .Z(new_n703));
  NAND3_X1  g502(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n693), .B1(new_n699), .B2(new_n704), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n573), .B(new_n700), .Z(new_n706));
  INV_X1    g505(.A(new_n693), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n691), .B1(new_n705), .B2(new_n708), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n706), .A2(new_n707), .ZN(new_n710));
  INV_X1    g509(.A(new_n691), .ZN(new_n711));
  AOI22_X1  g510(.A1(new_n706), .A2(new_n703), .B1(new_n695), .B2(new_n698), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n710), .B(new_n711), .C1(new_n712), .C2(new_n693), .ZN(new_n713));
  AOI21_X1  g512(.A(KEYINPUT109), .B1(new_n709), .B2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n709), .A2(new_n713), .A3(KEYINPUT109), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT96), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n655), .B1(new_n654), .B2(new_n657), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n659), .A2(new_n665), .A3(KEYINPUT17), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n719), .B(new_n582), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(G229gat), .A2(G233gat), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n581), .B1(new_n658), .B2(new_n666), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n654), .A2(new_n657), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT96), .B1(new_n725), .B2(new_n581), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n722), .B(new_n723), .C1(new_n724), .C2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT18), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n725), .A2(new_n581), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n719), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n582), .B1(new_n720), .B2(new_n721), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n733), .A2(KEYINPUT18), .A3(new_n723), .A4(new_n722), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n723), .B(KEYINPUT13), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n582), .A2(new_n676), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n735), .B1(new_n736), .B2(new_n730), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n729), .A2(new_n734), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(G113gat), .B(G141gat), .ZN(new_n740));
  INV_X1    g539(.A(G197gat), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(KEYINPUT11), .B(G169gat), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT12), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n739), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n737), .B1(new_n727), .B2(new_n728), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n748), .A2(new_n734), .A3(new_n745), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n718), .A2(new_n750), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n540), .A2(new_n688), .A3(new_n751), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n491), .A2(KEYINPUT110), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n491), .A2(KEYINPUT110), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G1gat), .ZN(G1324gat));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n752), .A2(new_n477), .ZN(new_n759));
  XNOR2_X1  g558(.A(KEYINPUT16), .B(G8gat), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n758), .B1(new_n761), .B2(KEYINPUT42), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT42), .ZN(new_n763));
  NOR4_X1   g562(.A1(new_n759), .A2(KEYINPUT111), .A3(new_n763), .A4(new_n760), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n759), .B2(G8gat), .ZN(new_n765));
  OAI22_X1  g564(.A1(new_n762), .A2(new_n764), .B1(new_n765), .B2(new_n761), .ZN(G1325gat));
  NAND2_X1  g565(.A1(new_n498), .A2(new_n501), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n752), .A2(G15gat), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n290), .ZN(new_n770));
  AOI21_X1  g569(.A(G15gat), .B1(new_n752), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n769), .A2(new_n771), .ZN(G1326gat));
  NAND2_X1  g571(.A1(new_n752), .A2(new_n496), .ZN(new_n773));
  XNOR2_X1  g572(.A(KEYINPUT43), .B(G22gat), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(G1327gat));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n598), .A2(new_n601), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(new_n751), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n540), .A2(new_n687), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n755), .A2(new_n632), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n776), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n781), .A2(KEYINPUT113), .A3(new_n632), .A4(new_n755), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XOR2_X1   g585(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n784), .A2(new_n785), .A3(new_n787), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT44), .B1(new_n540), .B2(new_n687), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n687), .B(KEYINPUT114), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n793), .A2(KEYINPUT44), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n408), .B1(new_n457), .B2(new_n466), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT93), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT35), .B1(new_n796), .B2(new_n467), .ZN(new_n797));
  AOI22_X1  g596(.A1(new_n797), .A2(new_n377), .B1(KEYINPUT35), .B2(new_n489), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n492), .A2(new_n496), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n539), .A2(new_n799), .A3(new_n767), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n794), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n780), .B1(new_n791), .B2(new_n801), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n802), .A2(new_n755), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n789), .B(new_n790), .C1(new_n632), .C2(new_n803), .ZN(G1328gat));
  NAND2_X1  g603(.A1(new_n477), .A2(new_n633), .ZN(new_n805));
  OR3_X1    g604(.A1(new_n782), .A2(KEYINPUT46), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT46), .B1(new_n782), .B2(new_n805), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n802), .A2(new_n477), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n806), .B(new_n807), .C1(new_n808), .C2(new_n633), .ZN(G1329gat));
  AOI21_X1  g608(.A(new_n661), .B1(new_n802), .B2(new_n768), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT47), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n781), .A2(new_n770), .A3(new_n661), .ZN(new_n812));
  OR3_X1    g611(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n811), .B1(new_n810), .B2(new_n812), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(G1330gat));
  AOI211_X1 g614(.A(new_n485), .B(new_n780), .C1(new_n791), .C2(new_n801), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT115), .B1(new_n816), .B2(new_n646), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n781), .A2(new_n646), .A3(new_n496), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(new_n816), .B2(new_n646), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT48), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n817), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  OAI221_X1 g620(.A(new_n818), .B1(KEYINPUT115), .B2(KEYINPUT48), .C1(new_n816), .C2(new_n646), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(G1331gat));
  NAND2_X1  g622(.A1(new_n476), .A2(new_n490), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n502), .A2(new_n539), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n688), .A2(new_n750), .A3(new_n718), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n755), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(new_n558), .ZN(G1332gat));
  NOR2_X1   g630(.A1(new_n828), .A2(new_n408), .ZN(new_n832));
  NOR2_X1   g631(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n833));
  AND2_X1   g632(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n835), .B1(new_n832), .B2(new_n833), .ZN(G1333gat));
  OAI21_X1  g635(.A(G71gat), .B1(new_n828), .B2(new_n767), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n770), .A2(new_n551), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n837), .B1(new_n828), .B2(new_n838), .ZN(new_n839));
  XOR2_X1   g638(.A(new_n839), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g639(.A1(new_n828), .A2(new_n485), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(new_n552), .ZN(G1335gat));
  INV_X1    g641(.A(new_n687), .ZN(new_n843));
  AND4_X1   g642(.A1(new_n734), .A2(new_n729), .A3(new_n738), .A4(new_n745), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n745), .B1(new_n748), .B2(new_n734), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n777), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT116), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n843), .B(new_n848), .C1(new_n798), .C2(new_n800), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT51), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n826), .A2(new_n851), .A3(new_n843), .A4(new_n848), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n850), .A2(new_n755), .A3(new_n717), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n848), .A2(new_n717), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n854), .B1(new_n791), .B2(new_n801), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n829), .A2(new_n445), .ZN(new_n856));
  AOI22_X1  g655(.A1(new_n853), .A2(new_n445), .B1(new_n855), .B2(new_n856), .ZN(G1336gat));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n408), .A2(G92gat), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n850), .A2(new_n717), .A3(new_n852), .A4(new_n859), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n855), .A2(new_n477), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n622), .A2(new_n623), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n858), .B(new_n860), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n860), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n862), .B1(new_n855), .B2(new_n477), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT52), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n863), .A2(new_n866), .ZN(G1337gat));
  NAND4_X1  g666(.A1(new_n850), .A2(new_n770), .A3(new_n717), .A4(new_n852), .ZN(new_n868));
  INV_X1    g667(.A(G99gat), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n767), .A2(new_n869), .ZN(new_n870));
  AOI22_X1  g669(.A1(new_n868), .A2(new_n869), .B1(new_n855), .B2(new_n870), .ZN(G1338gat));
  XNOR2_X1  g670(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(G106gat), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n485), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n850), .A2(new_n496), .A3(new_n717), .A4(new_n852), .ZN(new_n876));
  AOI221_X4 g675(.A(new_n873), .B1(new_n855), .B2(new_n875), .C1(new_n876), .C2(new_n874), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n874), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n855), .A2(new_n875), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n872), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n877), .A2(new_n880), .ZN(G1339gat));
  NOR3_X1   g680(.A1(new_n688), .A2(new_n750), .A3(new_n717), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n675), .A2(KEYINPUT108), .A3(new_n694), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n697), .B1(new_n628), .B2(new_n696), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n704), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n707), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n699), .A2(new_n693), .A3(new_n704), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(KEYINPUT54), .A3(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n711), .B1(new_n705), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n888), .A2(new_n890), .A3(KEYINPUT55), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n713), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT55), .B1(new_n888), .B2(new_n890), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n723), .B1(new_n733), .B2(new_n722), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n730), .A2(new_n736), .A3(new_n735), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n744), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n749), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n894), .A2(new_n792), .A3(new_n898), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n894), .A2(new_n750), .B1(new_n717), .B2(new_n898), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(new_n792), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n882), .B1(new_n901), .B2(new_n777), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n755), .A3(new_n408), .ZN(new_n904));
  INV_X1    g703(.A(new_n377), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(G113gat), .B1(new_n906), .B2(new_n846), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n485), .A2(new_n488), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n750), .A2(new_n251), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(G1340gat));
  OAI21_X1  g710(.A(G120gat), .B1(new_n906), .B2(new_n718), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n717), .A2(new_n252), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n912), .B1(new_n909), .B2(new_n913), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT118), .ZN(G1341gat));
  NOR3_X1   g714(.A1(new_n906), .A2(new_n259), .A3(new_n777), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n909), .A2(new_n777), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n259), .B2(new_n917), .ZN(G1342gat));
  NOR3_X1   g717(.A1(new_n909), .A2(G134gat), .A3(new_n687), .ZN(new_n919));
  XOR2_X1   g718(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n920));
  OR2_X1    g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(G134gat), .B1(new_n906), .B2(new_n687), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n919), .A2(new_n920), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(G1343gat));
  INV_X1    g723(.A(KEYINPUT120), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n891), .A2(new_n713), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n888), .A2(new_n890), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT55), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n926), .A2(new_n750), .A3(new_n929), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n709), .A2(KEYINPUT109), .A3(new_n713), .ZN(new_n931));
  OAI211_X1 g730(.A(new_n749), .B(new_n897), .C1(new_n931), .C2(new_n714), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n792), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n894), .A2(new_n792), .A3(new_n898), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n777), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n778), .A2(new_n687), .A3(new_n846), .A4(new_n718), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n485), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n925), .B1(new_n937), .B2(KEYINPUT57), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT57), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n485), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n929), .A2(new_n713), .A3(new_n891), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n932), .B1(new_n941), .B2(new_n846), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT121), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n930), .A2(KEYINPUT121), .A3(new_n932), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n944), .A2(new_n687), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n778), .B1(new_n946), .B2(new_n899), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n940), .B1(new_n947), .B2(new_n882), .ZN(new_n948));
  OAI211_X1 g747(.A(KEYINPUT120), .B(new_n939), .C1(new_n902), .C2(new_n485), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n938), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n755), .A2(new_n408), .A3(new_n767), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n950), .A2(new_n750), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(KEYINPUT122), .B1(new_n953), .B2(G141gat), .ZN(new_n954));
  INV_X1    g753(.A(new_n937), .ZN(new_n955));
  NOR4_X1   g754(.A1(new_n955), .A2(new_n951), .A3(G141gat), .A4(new_n846), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n956), .B1(new_n953), .B2(G141gat), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n954), .A2(new_n957), .A3(KEYINPUT58), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT58), .ZN(new_n959));
  AOI221_X4 g758(.A(new_n956), .B1(KEYINPUT122), .B2(new_n959), .C1(new_n953), .C2(G141gat), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n958), .A2(new_n960), .ZN(G1344gat));
  NOR2_X1   g760(.A1(new_n955), .A2(new_n951), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n962), .A2(new_n301), .A3(new_n717), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n950), .A2(new_n952), .ZN(new_n964));
  AOI211_X1 g763(.A(KEYINPUT59), .B(new_n301), .C1(new_n964), .C2(new_n717), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT59), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n894), .A2(new_n843), .A3(new_n898), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n778), .B1(new_n946), .B2(new_n967), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n939), .B(new_n496), .C1(new_n968), .C2(new_n882), .ZN(new_n969));
  OAI21_X1  g768(.A(KEYINPUT57), .B1(new_n902), .B2(new_n485), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n971), .A2(new_n717), .A3(new_n952), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n966), .B1(new_n972), .B2(G148gat), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n963), .B1(new_n965), .B2(new_n973), .ZN(G1345gat));
  AOI21_X1  g773(.A(G155gat), .B1(new_n962), .B2(new_n778), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n777), .A2(new_n296), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n975), .B1(new_n964), .B2(new_n976), .ZN(G1346gat));
  NAND3_X1  g776(.A1(new_n962), .A2(new_n297), .A3(new_n843), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n978), .B(KEYINPUT123), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n964), .A2(new_n792), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n979), .B1(new_n980), .B2(new_n297), .ZN(G1347gat));
  NAND2_X1  g780(.A1(new_n829), .A2(new_n477), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(KEYINPUT124), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n755), .A2(new_n408), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT124), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n903), .A2(new_n377), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n246), .B1(new_n989), .B2(new_n750), .ZN(new_n990));
  NOR3_X1   g789(.A1(new_n982), .A2(new_n908), .A3(new_n902), .ZN(new_n991));
  AND3_X1   g790(.A1(new_n991), .A2(new_n246), .A3(new_n750), .ZN(new_n992));
  OR2_X1    g791(.A1(new_n990), .A2(new_n992), .ZN(G1348gat));
  AOI21_X1  g792(.A(G176gat), .B1(new_n991), .B2(new_n717), .ZN(new_n994));
  AND2_X1   g793(.A1(new_n717), .A2(new_n245), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n994), .B1(new_n989), .B2(new_n995), .ZN(G1349gat));
  NAND3_X1  g795(.A1(new_n991), .A2(new_n212), .A3(new_n778), .ZN(new_n997));
  NOR3_X1   g796(.A1(new_n987), .A2(new_n988), .A3(new_n777), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n997), .B1(new_n998), .B2(new_n208), .ZN(new_n999));
  XNOR2_X1  g798(.A(new_n999), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g799(.A(new_n218), .B1(new_n989), .B2(new_n843), .ZN(new_n1001));
  XOR2_X1   g800(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n1002));
  OR2_X1    g801(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n991), .A2(new_n218), .A3(new_n792), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(G1351gat));
  NOR2_X1   g805(.A1(new_n987), .A2(new_n768), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1007), .A2(new_n971), .ZN(new_n1008));
  OAI21_X1  g807(.A(G197gat), .B1(new_n1008), .B2(new_n846), .ZN(new_n1009));
  NOR3_X1   g808(.A1(new_n982), .A2(new_n955), .A3(new_n768), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n1010), .A2(new_n741), .A3(new_n750), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1009), .A2(new_n1011), .ZN(G1352gat));
  NAND3_X1  g811(.A1(new_n1007), .A2(new_n717), .A3(new_n971), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1013), .A2(G204gat), .ZN(new_n1014));
  INV_X1    g813(.A(new_n1010), .ZN(new_n1015));
  NOR2_X1   g814(.A1(new_n718), .A2(G204gat), .ZN(new_n1016));
  INV_X1    g815(.A(new_n1016), .ZN(new_n1017));
  OAI21_X1  g816(.A(KEYINPUT62), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  OR3_X1    g817(.A1(new_n1015), .A2(KEYINPUT62), .A3(new_n1017), .ZN(new_n1019));
  NAND3_X1  g818(.A1(new_n1014), .A2(new_n1018), .A3(new_n1019), .ZN(G1353gat));
  NAND3_X1  g819(.A1(new_n1010), .A2(new_n543), .A3(new_n778), .ZN(new_n1021));
  NAND3_X1  g820(.A1(new_n1007), .A2(new_n778), .A3(new_n971), .ZN(new_n1022));
  AND3_X1   g821(.A1(new_n1022), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1023));
  AOI21_X1  g822(.A(KEYINPUT63), .B1(new_n1022), .B2(G211gat), .ZN(new_n1024));
  OAI21_X1  g823(.A(new_n1021), .B1(new_n1023), .B2(new_n1024), .ZN(G1354gat));
  INV_X1    g824(.A(G218gat), .ZN(new_n1026));
  NOR3_X1   g825(.A1(new_n1008), .A2(new_n1026), .A3(new_n687), .ZN(new_n1027));
  OAI21_X1  g826(.A(new_n1026), .B1(new_n1015), .B2(new_n793), .ZN(new_n1028));
  AND2_X1   g827(.A1(new_n1028), .A2(KEYINPUT126), .ZN(new_n1029));
  NOR2_X1   g828(.A1(new_n1028), .A2(KEYINPUT126), .ZN(new_n1030));
  NOR3_X1   g829(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .ZN(G1355gat));
endmodule


