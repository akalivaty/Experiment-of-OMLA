

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722;

  INV_X1 U369 ( .A(G953), .ZN(n708) );
  XOR2_X1 U370 ( .A(n655), .B(KEYINPUT62), .Z(n347) );
  XNOR2_X2 U371 ( .A(n440), .B(n439), .ZN(n377) );
  XNOR2_X2 U372 ( .A(n473), .B(n472), .ZN(n619) );
  NOR2_X1 U373 ( .A1(n719), .A2(n550), .ZN(n551) );
  XNOR2_X1 U374 ( .A(n529), .B(KEYINPUT117), .ZN(n719) );
  INV_X1 U375 ( .A(n619), .ZN(n592) );
  INV_X1 U376 ( .A(KEYINPUT39), .ZN(n389) );
  NOR2_X1 U377 ( .A1(n715), .A2(n717), .ZN(n537) );
  NOR2_X1 U378 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U379 ( .A(n388), .B(n358), .ZN(n715) );
  NOR2_X1 U380 ( .A1(n530), .A2(n670), .ZN(n388) );
  XNOR2_X1 U381 ( .A(n390), .B(n389), .ZN(n530) );
  XNOR2_X1 U382 ( .A(n563), .B(KEYINPUT0), .ZN(n590) );
  AND2_X1 U383 ( .A1(n427), .A2(n522), .ZN(n426) );
  NOR2_X1 U384 ( .A1(n589), .A2(n521), .ZN(n522) );
  XNOR2_X1 U385 ( .A(n592), .B(n474), .ZN(n575) );
  XNOR2_X1 U386 ( .A(n370), .B(n442), .ZN(n704) );
  XNOR2_X1 U387 ( .A(n419), .B(G131), .ZN(n449) );
  XNOR2_X1 U388 ( .A(G125), .B(G146), .ZN(n441) );
  NOR2_X1 U389 ( .A1(G953), .A2(G237), .ZN(n468) );
  XNOR2_X1 U390 ( .A(n378), .B(n462), .ZN(n705) );
  XNOR2_X1 U391 ( .A(n433), .B(KEYINPUT4), .ZN(n378) );
  XNOR2_X1 U392 ( .A(G469), .B(KEYINPUT69), .ZN(n439) );
  XNOR2_X1 U393 ( .A(KEYINPUT71), .B(G472), .ZN(n472) );
  XNOR2_X1 U394 ( .A(n506), .B(G134), .ZN(n462) );
  XNOR2_X1 U395 ( .A(n435), .B(G107), .ZN(n503) );
  XNOR2_X1 U396 ( .A(G104), .B(G110), .ZN(n435) );
  NAND2_X2 U397 ( .A1(n398), .A2(n359), .ZN(n397) );
  NAND2_X1 U398 ( .A1(n399), .A2(n696), .ZN(n398) );
  NOR2_X1 U399 ( .A1(n606), .A2(n605), .ZN(n396) );
  NAND2_X1 U400 ( .A1(n364), .A2(n608), .ZN(n407) );
  INV_X1 U401 ( .A(n610), .ZN(n364) );
  XNOR2_X1 U402 ( .A(G113), .B(G101), .ZN(n465) );
  OR2_X1 U403 ( .A1(n716), .A2(KEYINPUT44), .ZN(n385) );
  NOR2_X1 U404 ( .A1(n575), .A2(n584), .ZN(n576) );
  XNOR2_X1 U405 ( .A(n467), .B(n428), .ZN(n655) );
  XNOR2_X1 U406 ( .A(n484), .B(n429), .ZN(n485) );
  XNOR2_X1 U407 ( .A(n704), .B(n351), .ZN(n486) );
  XNOR2_X1 U408 ( .A(G116), .B(G107), .ZN(n455) );
  XNOR2_X1 U409 ( .A(n458), .B(n457), .ZN(n481) );
  XNOR2_X1 U410 ( .A(KEYINPUT81), .B(KEYINPUT8), .ZN(n457) );
  XNOR2_X1 U411 ( .A(n453), .B(n704), .ZN(n649) );
  XNOR2_X1 U412 ( .A(n420), .B(n418), .ZN(n451) );
  XNOR2_X1 U413 ( .A(n705), .B(n434), .ZN(n467) );
  INV_X1 U414 ( .A(G146), .ZN(n434) );
  XNOR2_X1 U415 ( .A(KEYINPUT75), .B(G140), .ZN(n395) );
  XNOR2_X1 U416 ( .A(n425), .B(n424), .ZN(n506) );
  INV_X1 U417 ( .A(G143), .ZN(n424) );
  XNOR2_X1 U418 ( .A(KEYINPUT77), .B(G128), .ZN(n425) );
  NOR2_X1 U419 ( .A1(n590), .A2(n566), .ZN(n567) );
  XNOR2_X1 U420 ( .A(G478), .B(n463), .ZN(n539) );
  NAND2_X1 U421 ( .A1(n400), .A2(n352), .ZN(n409) );
  XNOR2_X1 U422 ( .A(n534), .B(KEYINPUT28), .ZN(n400) );
  NAND2_X1 U423 ( .A1(n397), .A2(n350), .ZN(n393) );
  XNOR2_X1 U424 ( .A(n412), .B(n505), .ZN(n695) );
  XNOR2_X1 U425 ( .A(n413), .B(n503), .ZN(n412) );
  XNOR2_X1 U426 ( .A(n504), .B(KEYINPUT72), .ZN(n413) );
  XNOR2_X1 U427 ( .A(n414), .B(n695), .ZN(n678) );
  XNOR2_X1 U428 ( .A(n415), .B(n368), .ZN(n414) );
  XNOR2_X1 U429 ( .A(n509), .B(KEYINPUT4), .ZN(n415) );
  XNOR2_X1 U430 ( .A(n506), .B(n369), .ZN(n368) );
  INV_X1 U431 ( .A(KEYINPUT67), .ZN(n419) );
  OR2_X1 U432 ( .A1(G902), .A2(G237), .ZN(n511) );
  XOR2_X1 U433 ( .A(G137), .B(G128), .Z(n483) );
  XNOR2_X1 U434 ( .A(G119), .B(G110), .ZN(n482) );
  XNOR2_X1 U435 ( .A(G113), .B(G104), .ZN(n443) );
  XOR2_X1 U436 ( .A(G143), .B(G122), .Z(n444) );
  XNOR2_X1 U437 ( .A(KEYINPUT11), .B(KEYINPUT101), .ZN(n445) );
  XOR2_X1 U438 ( .A(KEYINPUT12), .B(KEYINPUT99), .Z(n446) );
  XNOR2_X1 U439 ( .A(n450), .B(KEYINPUT100), .ZN(n420) );
  INV_X1 U440 ( .A(n449), .ZN(n418) );
  INV_X1 U441 ( .A(G140), .ZN(n371) );
  AND2_X1 U442 ( .A1(n706), .A2(n646), .ZN(n399) );
  NAND2_X1 U443 ( .A1(G234), .A2(G237), .ZN(n491) );
  INV_X1 U444 ( .A(n407), .ZN(n363) );
  INV_X1 U445 ( .A(KEYINPUT38), .ZN(n365) );
  NAND2_X1 U446 ( .A1(n407), .A2(n406), .ZN(n404) );
  NOR2_X1 U447 ( .A1(n519), .A2(n564), .ZN(n616) );
  XNOR2_X1 U448 ( .A(n410), .B(n466), .ZN(n505) );
  XNOR2_X1 U449 ( .A(n465), .B(n411), .ZN(n410) );
  INV_X1 U450 ( .A(KEYINPUT3), .ZN(n411) );
  XNOR2_X1 U451 ( .A(n441), .B(KEYINPUT18), .ZN(n369) );
  XNOR2_X1 U452 ( .A(n508), .B(n507), .ZN(n509) );
  INV_X1 U453 ( .A(KEYINPUT17), .ZN(n507) );
  NAND2_X1 U454 ( .A1(n403), .A2(n401), .ZN(n636) );
  AND2_X1 U455 ( .A1(n405), .A2(n404), .ZN(n403) );
  OR2_X1 U456 ( .A1(n408), .A2(n402), .ZN(n401) );
  NAND2_X1 U457 ( .A1(n408), .A2(n406), .ZN(n405) );
  XNOR2_X1 U458 ( .A(n377), .B(KEYINPUT1), .ZN(n617) );
  XNOR2_X1 U459 ( .A(n423), .B(n421), .ZN(n531) );
  XNOR2_X1 U460 ( .A(n454), .B(n422), .ZN(n421) );
  OR2_X1 U461 ( .A1(n649), .A2(G902), .ZN(n423) );
  INV_X1 U462 ( .A(G475), .ZN(n422) );
  XNOR2_X1 U463 ( .A(n519), .B(n372), .ZN(n621) );
  INV_X1 U464 ( .A(KEYINPUT107), .ZN(n372) );
  XNOR2_X1 U465 ( .A(n367), .B(n366), .ZN(n461) );
  NAND2_X1 U466 ( .A1(n481), .A2(G217), .ZN(n366) );
  XNOR2_X1 U467 ( .A(n460), .B(n459), .ZN(n367) );
  XNOR2_X1 U468 ( .A(n503), .B(n394), .ZN(n437) );
  XNOR2_X1 U469 ( .A(n436), .B(n395), .ZN(n394) );
  XNOR2_X1 U470 ( .A(n381), .B(n380), .ZN(n379) );
  INV_X1 U471 ( .A(KEYINPUT80), .ZN(n380) );
  XNOR2_X1 U472 ( .A(n582), .B(n387), .ZN(n716) );
  XNOR2_X1 U473 ( .A(n588), .B(n587), .ZN(n675) );
  XNOR2_X1 U474 ( .A(n586), .B(KEYINPUT98), .ZN(n587) );
  INV_X1 U475 ( .A(n409), .ZN(n544) );
  XNOR2_X1 U476 ( .A(n595), .B(n417), .ZN(n416) );
  INV_X1 U477 ( .A(KEYINPUT108), .ZN(n417) );
  NAND2_X1 U478 ( .A1(n392), .A2(n680), .ZN(n391) );
  XNOR2_X1 U479 ( .A(n393), .B(n347), .ZN(n392) );
  INV_X1 U480 ( .A(KEYINPUT126), .ZN(n373) );
  NAND2_X1 U481 ( .A1(n375), .A2(n680), .ZN(n374) );
  XNOR2_X1 U482 ( .A(n376), .B(n360), .ZN(n375) );
  NOR2_X1 U483 ( .A1(n653), .A2(n693), .ZN(n654) );
  AND2_X1 U484 ( .A1(n681), .A2(n680), .ZN(n682) );
  AND2_X1 U485 ( .A1(n523), .A2(n522), .ZN(n348) );
  AND2_X1 U486 ( .A1(n592), .A2(n519), .ZN(n349) );
  AND2_X1 U487 ( .A1(n648), .A2(G472), .ZN(n350) );
  XOR2_X1 U488 ( .A(n480), .B(n479), .Z(n351) );
  XOR2_X1 U489 ( .A(n377), .B(KEYINPUT113), .Z(n352) );
  XOR2_X1 U490 ( .A(KEYINPUT68), .B(n498), .Z(n353) );
  AND2_X1 U491 ( .A1(n648), .A2(G210), .ZN(n354) );
  AND2_X1 U492 ( .A1(n648), .A2(G475), .ZN(n355) );
  XOR2_X1 U493 ( .A(n554), .B(n553), .Z(n356) );
  AND2_X1 U494 ( .A1(n348), .A2(n542), .ZN(n357) );
  XNOR2_X1 U495 ( .A(n524), .B(n365), .ZN(n408) );
  INV_X1 U496 ( .A(n532), .ZN(n406) );
  XNOR2_X1 U497 ( .A(KEYINPUT114), .B(KEYINPUT40), .ZN(n358) );
  XOR2_X1 U498 ( .A(n647), .B(KEYINPUT65), .Z(n359) );
  XNOR2_X1 U499 ( .A(n692), .B(KEYINPUT125), .ZN(n360) );
  XOR2_X1 U500 ( .A(n678), .B(n677), .Z(n361) );
  NOR2_X1 U501 ( .A1(G952), .A2(n708), .ZN(n693) );
  XNOR2_X1 U502 ( .A(KEYINPUT63), .B(KEYINPUT86), .ZN(n362) );
  NAND2_X1 U503 ( .A1(n363), .A2(n532), .ZN(n402) );
  AND2_X2 U504 ( .A1(n397), .A2(n648), .ZN(n688) );
  NAND2_X1 U505 ( .A1(n397), .A2(n354), .ZN(n679) );
  NAND2_X1 U506 ( .A1(n397), .A2(n355), .ZN(n652) );
  NAND2_X1 U507 ( .A1(n688), .A2(G217), .ZN(n376) );
  XNOR2_X1 U508 ( .A(n441), .B(n371), .ZN(n370) );
  AND2_X1 U509 ( .A1(n519), .A2(n353), .ZN(n533) );
  XNOR2_X1 U510 ( .A(n374), .B(n373), .ZN(G66) );
  NAND2_X1 U511 ( .A1(n377), .A2(n616), .ZN(n589) );
  NAND2_X1 U512 ( .A1(n379), .A2(n648), .ZN(n642) );
  NAND2_X1 U513 ( .A1(n382), .A2(n356), .ZN(n381) );
  XNOR2_X1 U514 ( .A(n602), .B(n383), .ZN(n382) );
  INV_X1 U515 ( .A(KEYINPUT82), .ZN(n383) );
  NAND2_X1 U516 ( .A1(n384), .A2(n600), .ZN(n601) );
  NAND2_X1 U517 ( .A1(n386), .A2(n385), .ZN(n384) );
  NAND2_X1 U518 ( .A1(n583), .A2(n716), .ZN(n386) );
  INV_X1 U519 ( .A(KEYINPUT35), .ZN(n387) );
  NAND2_X1 U520 ( .A1(n426), .A2(n523), .ZN(n390) );
  XNOR2_X1 U521 ( .A(n391), .B(n362), .ZN(G57) );
  NAND2_X1 U522 ( .A1(n396), .A2(n696), .ZN(n648) );
  XNOR2_X2 U523 ( .A(n601), .B(KEYINPUT45), .ZN(n696) );
  NOR2_X1 U524 ( .A1(n636), .A2(n409), .ZN(n536) );
  NAND2_X1 U525 ( .A1(n427), .A2(n608), .ZN(n611) );
  NAND2_X1 U526 ( .A1(n416), .A2(n349), .ZN(n663) );
  NAND2_X1 U527 ( .A1(n568), .A2(n569), .ZN(n595) );
  INV_X1 U528 ( .A(n408), .ZN(n427) );
  XNOR2_X1 U529 ( .A(n505), .B(n471), .ZN(n428) );
  XNOR2_X1 U530 ( .A(n652), .B(n432), .ZN(n653) );
  XNOR2_X1 U531 ( .A(n515), .B(n514), .ZN(n524) );
  XNOR2_X1 U532 ( .A(n467), .B(n438), .ZN(n684) );
  XOR2_X1 U533 ( .A(n483), .B(n482), .Z(n429) );
  XNOR2_X1 U534 ( .A(KEYINPUT111), .B(KEYINPUT30), .ZN(n430) );
  OR2_X1 U535 ( .A1(n530), .A2(n664), .ZN(n431) );
  XOR2_X1 U536 ( .A(n651), .B(n650), .Z(n432) );
  XNOR2_X1 U537 ( .A(n486), .B(n485), .ZN(n692) );
  XNOR2_X1 U538 ( .A(n437), .B(G101), .ZN(n438) );
  INV_X1 U539 ( .A(KEYINPUT31), .ZN(n586) );
  XOR2_X1 U540 ( .A(G137), .B(n449), .Z(n433) );
  NAND2_X1 U541 ( .A1(G227), .A2(n708), .ZN(n436) );
  NOR2_X1 U542 ( .A1(n684), .A2(G902), .ZN(n440) );
  INV_X1 U543 ( .A(n617), .ZN(n569) );
  XOR2_X1 U544 ( .A(KEYINPUT66), .B(KEYINPUT10), .Z(n442) );
  XNOR2_X1 U545 ( .A(n444), .B(n443), .ZN(n448) );
  XNOR2_X1 U546 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U547 ( .A(n448), .B(n447), .ZN(n452) );
  NAND2_X1 U548 ( .A1(n468), .A2(G214), .ZN(n450) );
  XNOR2_X1 U549 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U550 ( .A(KEYINPUT13), .B(KEYINPUT102), .ZN(n454) );
  XOR2_X1 U551 ( .A(KEYINPUT103), .B(G122), .Z(n456) );
  XNOR2_X1 U552 ( .A(n456), .B(n455), .ZN(n460) );
  XOR2_X1 U553 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n459) );
  NAND2_X1 U554 ( .A1(n708), .A2(G234), .ZN(n458) );
  XOR2_X1 U555 ( .A(n462), .B(n461), .Z(n690) );
  NOR2_X1 U556 ( .A1(G902), .A2(n690), .ZN(n463) );
  NAND2_X1 U557 ( .A1(n531), .A2(n539), .ZN(n464) );
  XNOR2_X1 U558 ( .A(n464), .B(KEYINPUT104), .ZN(n670) );
  XOR2_X1 U559 ( .A(G116), .B(G119), .Z(n466) );
  XOR2_X1 U560 ( .A(KEYINPUT95), .B(KEYINPUT5), .Z(n470) );
  NAND2_X1 U561 ( .A1(n468), .A2(G210), .ZN(n469) );
  XNOR2_X1 U562 ( .A(n470), .B(n469), .ZN(n471) );
  NOR2_X1 U563 ( .A1(n655), .A2(G902), .ZN(n473) );
  INV_X1 U564 ( .A(KEYINPUT6), .ZN(n474) );
  INV_X1 U565 ( .A(n575), .ZN(n596) );
  XOR2_X1 U566 ( .A(KEYINPUT93), .B(KEYINPUT25), .Z(n478) );
  XOR2_X1 U567 ( .A(G902), .B(KEYINPUT15), .Z(n475) );
  XNOR2_X1 U568 ( .A(KEYINPUT87), .B(n475), .ZN(n510) );
  NAND2_X1 U569 ( .A1(n510), .A2(G234), .ZN(n476) );
  XNOR2_X1 U570 ( .A(n476), .B(KEYINPUT20), .ZN(n489) );
  NAND2_X1 U571 ( .A1(n489), .A2(G217), .ZN(n477) );
  XNOR2_X1 U572 ( .A(n478), .B(n477), .ZN(n488) );
  XOR2_X1 U573 ( .A(KEYINPUT92), .B(KEYINPUT24), .Z(n480) );
  XNOR2_X1 U574 ( .A(KEYINPUT23), .B(KEYINPUT74), .ZN(n479) );
  NAND2_X1 U575 ( .A1(G221), .A2(n481), .ZN(n484) );
  NOR2_X1 U576 ( .A1(G902), .A2(n692), .ZN(n487) );
  XOR2_X1 U577 ( .A(n488), .B(n487), .Z(n519) );
  NAND2_X1 U578 ( .A1(n489), .A2(G221), .ZN(n490) );
  XNOR2_X1 U579 ( .A(n490), .B(KEYINPUT21), .ZN(n620) );
  INV_X1 U580 ( .A(n620), .ZN(n497) );
  XOR2_X1 U581 ( .A(KEYINPUT73), .B(KEYINPUT14), .Z(n492) );
  XNOR2_X1 U582 ( .A(n492), .B(n491), .ZN(n494) );
  NAND2_X1 U583 ( .A1(n494), .A2(G952), .ZN(n635) );
  NOR2_X1 U584 ( .A1(G953), .A2(n635), .ZN(n493) );
  XNOR2_X1 U585 ( .A(KEYINPUT89), .B(n493), .ZN(n555) );
  NAND2_X1 U586 ( .A1(G902), .A2(n494), .ZN(n557) );
  NOR2_X1 U587 ( .A1(G900), .A2(n557), .ZN(n495) );
  NAND2_X1 U588 ( .A1(G953), .A2(n495), .ZN(n496) );
  NAND2_X1 U589 ( .A1(n555), .A2(n496), .ZN(n520) );
  NAND2_X1 U590 ( .A1(n497), .A2(n520), .ZN(n498) );
  NAND2_X1 U591 ( .A1(n596), .A2(n533), .ZN(n499) );
  XNOR2_X1 U592 ( .A(n499), .B(KEYINPUT109), .ZN(n500) );
  NAND2_X1 U593 ( .A1(G214), .A2(n511), .ZN(n608) );
  NAND2_X1 U594 ( .A1(n500), .A2(n608), .ZN(n526) );
  NOR2_X1 U595 ( .A1(n670), .A2(n526), .ZN(n501) );
  NAND2_X1 U596 ( .A1(n569), .A2(n501), .ZN(n502) );
  XNOR2_X1 U597 ( .A(n502), .B(KEYINPUT43), .ZN(n516) );
  XOR2_X1 U598 ( .A(KEYINPUT16), .B(G122), .Z(n504) );
  NAND2_X1 U599 ( .A1(G224), .A2(n708), .ZN(n508) );
  INV_X1 U600 ( .A(n510), .ZN(n646) );
  NOR2_X1 U601 ( .A1(n678), .A2(n646), .ZN(n515) );
  XOR2_X1 U602 ( .A(KEYINPUT78), .B(KEYINPUT88), .Z(n513) );
  NAND2_X1 U603 ( .A1(G210), .A2(n511), .ZN(n512) );
  XNOR2_X1 U604 ( .A(n513), .B(n512), .ZN(n514) );
  NAND2_X1 U605 ( .A1(n516), .A2(n524), .ZN(n517) );
  XNOR2_X1 U606 ( .A(KEYINPUT110), .B(n517), .ZN(n718) );
  NAND2_X1 U607 ( .A1(n619), .A2(n608), .ZN(n518) );
  XNOR2_X1 U608 ( .A(n518), .B(n430), .ZN(n523) );
  XNOR2_X1 U609 ( .A(n620), .B(KEYINPUT94), .ZN(n564) );
  INV_X1 U610 ( .A(n520), .ZN(n521) );
  NOR2_X1 U611 ( .A1(n539), .A2(n531), .ZN(n674) );
  INV_X1 U612 ( .A(n674), .ZN(n664) );
  AND2_X1 U613 ( .A1(n718), .A2(n431), .ZN(n552) );
  INV_X1 U614 ( .A(n670), .ZN(n672) );
  INV_X1 U615 ( .A(n524), .ZN(n542) );
  NAND2_X1 U616 ( .A1(n672), .A2(n542), .ZN(n525) );
  XNOR2_X1 U617 ( .A(n527), .B(KEYINPUT36), .ZN(n528) );
  NAND2_X1 U618 ( .A1(n528), .A2(n617), .ZN(n529) );
  INV_X1 U619 ( .A(n531), .ZN(n538) );
  NAND2_X1 U620 ( .A1(n538), .A2(n539), .ZN(n610) );
  XOR2_X1 U621 ( .A(KEYINPUT41), .B(KEYINPUT115), .Z(n532) );
  AND2_X1 U622 ( .A1(n619), .A2(n533), .ZN(n534) );
  XNOR2_X1 U623 ( .A(KEYINPUT116), .B(KEYINPUT42), .ZN(n535) );
  XNOR2_X1 U624 ( .A(n536), .B(n535), .ZN(n717) );
  XNOR2_X1 U625 ( .A(n537), .B(KEYINPUT46), .ZN(n549) );
  NOR2_X1 U626 ( .A1(n539), .A2(n538), .ZN(n580) );
  INV_X1 U627 ( .A(n580), .ZN(n541) );
  XOR2_X1 U628 ( .A(KEYINPUT112), .B(n357), .Z(n540) );
  NOR2_X1 U629 ( .A1(n541), .A2(n540), .ZN(n668) );
  NAND2_X1 U630 ( .A1(n542), .A2(n608), .ZN(n543) );
  XNOR2_X1 U631 ( .A(n543), .B(KEYINPUT19), .ZN(n562) );
  NAND2_X1 U632 ( .A1(n544), .A2(n562), .ZN(n669) );
  NAND2_X1 U633 ( .A1(n664), .A2(n670), .ZN(n545) );
  XNOR2_X1 U634 ( .A(n545), .B(KEYINPUT105), .ZN(n612) );
  NOR2_X1 U635 ( .A1(n669), .A2(n612), .ZN(n546) );
  XOR2_X1 U636 ( .A(KEYINPUT47), .B(n546), .Z(n547) );
  NOR2_X1 U637 ( .A1(n668), .A2(n547), .ZN(n548) );
  NAND2_X1 U638 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U639 ( .A(n551), .B(KEYINPUT48), .ZN(n603) );
  AND2_X2 U640 ( .A1(n552), .A2(n603), .ZN(n706) );
  NOR2_X1 U641 ( .A1(KEYINPUT2), .A2(n706), .ZN(n554) );
  INV_X1 U642 ( .A(KEYINPUT83), .ZN(n553) );
  NOR2_X1 U643 ( .A1(KEYINPUT44), .A2(KEYINPUT85), .ZN(n574) );
  INV_X1 U644 ( .A(n555), .ZN(n559) );
  NOR2_X1 U645 ( .A1(G898), .A2(n708), .ZN(n556) );
  XOR2_X1 U646 ( .A(KEYINPUT90), .B(n556), .Z(n694) );
  NOR2_X1 U647 ( .A1(n694), .A2(n557), .ZN(n558) );
  NOR2_X1 U648 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U649 ( .A(KEYINPUT91), .B(n560), .ZN(n561) );
  NAND2_X1 U650 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U651 ( .A1(n610), .A2(n564), .ZN(n565) );
  XOR2_X1 U652 ( .A(KEYINPUT106), .B(n565), .Z(n566) );
  XNOR2_X1 U653 ( .A(KEYINPUT22), .B(n567), .ZN(n568) );
  AND2_X1 U654 ( .A1(n568), .A2(n621), .ZN(n571) );
  NOR2_X1 U655 ( .A1(n569), .A2(n596), .ZN(n570) );
  NAND2_X1 U656 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U657 ( .A(KEYINPUT32), .B(n572), .ZN(n722) );
  NAND2_X1 U658 ( .A1(n663), .A2(n722), .ZN(n573) );
  XNOR2_X1 U659 ( .A(n574), .B(n573), .ZN(n583) );
  NAND2_X1 U660 ( .A1(n616), .A2(n617), .ZN(n584) );
  XNOR2_X1 U661 ( .A(n576), .B(KEYINPUT33), .ZN(n607) );
  NOR2_X1 U662 ( .A1(n590), .A2(n607), .ZN(n579) );
  XNOR2_X1 U663 ( .A(KEYINPUT70), .B(KEYINPUT34), .ZN(n577) );
  XNOR2_X1 U664 ( .A(n577), .B(KEYINPUT76), .ZN(n578) );
  XNOR2_X1 U665 ( .A(n579), .B(n578), .ZN(n581) );
  NAND2_X1 U666 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U667 ( .A1(n584), .A2(n592), .ZN(n585) );
  XNOR2_X1 U668 ( .A(KEYINPUT97), .B(n585), .ZN(n627) );
  NOR2_X1 U669 ( .A1(n590), .A2(n627), .ZN(n588) );
  NOR2_X1 U670 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U671 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U672 ( .A(KEYINPUT96), .B(n593), .Z(n658) );
  NOR2_X1 U673 ( .A1(n675), .A2(n658), .ZN(n594) );
  NOR2_X1 U674 ( .A1(n612), .A2(n594), .ZN(n599) );
  NOR2_X1 U675 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U676 ( .A(KEYINPUT84), .B(n597), .Z(n598) );
  NOR2_X1 U677 ( .A1(n621), .A2(n598), .ZN(n656) );
  NOR2_X1 U678 ( .A1(n599), .A2(n656), .ZN(n600) );
  NOR2_X1 U679 ( .A1(n696), .A2(KEYINPUT2), .ZN(n602) );
  NAND2_X1 U680 ( .A1(n603), .A2(n718), .ZN(n606) );
  NAND2_X1 U681 ( .A1(KEYINPUT2), .A2(n431), .ZN(n604) );
  XOR2_X1 U682 ( .A(KEYINPUT79), .B(n604), .Z(n605) );
  NOR2_X1 U683 ( .A1(n427), .A2(n608), .ZN(n609) );
  NOR2_X1 U684 ( .A1(n610), .A2(n609), .ZN(n614) );
  NOR2_X1 U685 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U686 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U687 ( .A1(n607), .A2(n615), .ZN(n632) );
  OR2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U689 ( .A(n618), .B(KEYINPUT50), .ZN(n626) );
  XNOR2_X1 U690 ( .A(KEYINPUT49), .B(KEYINPUT121), .ZN(n623) );
  NAND2_X1 U691 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U692 ( .A(n623), .B(n622), .Z(n624) );
  NOR2_X1 U693 ( .A1(n619), .A2(n624), .ZN(n625) );
  NAND2_X1 U694 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U695 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U696 ( .A(KEYINPUT51), .B(n629), .ZN(n630) );
  NOR2_X1 U697 ( .A1(n636), .A2(n630), .ZN(n631) );
  NOR2_X1 U698 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U699 ( .A(n633), .B(KEYINPUT52), .ZN(n634) );
  NOR2_X1 U700 ( .A1(n635), .A2(n634), .ZN(n639) );
  OR2_X1 U701 ( .A1(n636), .A2(n607), .ZN(n637) );
  XOR2_X1 U702 ( .A(KEYINPUT122), .B(n637), .Z(n638) );
  OR2_X1 U703 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U704 ( .A1(n640), .A2(G953), .ZN(n641) );
  AND2_X1 U705 ( .A1(n642), .A2(n641), .ZN(n645) );
  INV_X1 U706 ( .A(KEYINPUT123), .ZN(n643) );
  XNOR2_X1 U707 ( .A(n643), .B(KEYINPUT53), .ZN(n644) );
  XNOR2_X1 U708 ( .A(n645), .B(n644), .ZN(G75) );
  NAND2_X1 U709 ( .A1(n646), .A2(KEYINPUT2), .ZN(n647) );
  XNOR2_X1 U710 ( .A(KEYINPUT124), .B(KEYINPUT64), .ZN(n651) );
  XNOR2_X1 U711 ( .A(n649), .B(KEYINPUT59), .ZN(n650) );
  XNOR2_X1 U712 ( .A(n654), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U713 ( .A(G101), .B(n656), .Z(G3) );
  NAND2_X1 U714 ( .A1(n658), .A2(n672), .ZN(n657) );
  XNOR2_X1 U715 ( .A(n657), .B(G104), .ZN(G6) );
  XNOR2_X1 U716 ( .A(G107), .B(KEYINPUT118), .ZN(n662) );
  XOR2_X1 U717 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n660) );
  NAND2_X1 U718 ( .A1(n674), .A2(n658), .ZN(n659) );
  XNOR2_X1 U719 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U720 ( .A(n662), .B(n661), .ZN(G9) );
  XNOR2_X1 U721 ( .A(n663), .B(G110), .ZN(G12) );
  NOR2_X1 U722 ( .A1(n664), .A2(n669), .ZN(n666) );
  XNOR2_X1 U723 ( .A(KEYINPUT119), .B(KEYINPUT29), .ZN(n665) );
  XNOR2_X1 U724 ( .A(n666), .B(n665), .ZN(n667) );
  XOR2_X1 U725 ( .A(G128), .B(n667), .Z(G30) );
  XOR2_X1 U726 ( .A(G143), .B(n668), .Z(G45) );
  NOR2_X1 U727 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U728 ( .A(G146), .B(n671), .Z(G48) );
  NAND2_X1 U729 ( .A1(n672), .A2(n675), .ZN(n673) );
  XNOR2_X1 U730 ( .A(G113), .B(n673), .ZN(G15) );
  NAND2_X1 U731 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U732 ( .A(n676), .B(G116), .ZN(G18) );
  XNOR2_X1 U733 ( .A(G134), .B(n431), .ZN(G36) );
  XOR2_X1 U734 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n677) );
  XNOR2_X1 U735 ( .A(n679), .B(n361), .ZN(n681) );
  INV_X1 U736 ( .A(n693), .ZN(n680) );
  XNOR2_X1 U737 ( .A(n682), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U738 ( .A1(n688), .A2(G469), .ZN(n686) );
  XOR2_X1 U739 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n683) );
  XNOR2_X1 U740 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U741 ( .A(n686), .B(n685), .ZN(n687) );
  NOR2_X1 U742 ( .A1(n693), .A2(n687), .ZN(G54) );
  NAND2_X1 U743 ( .A1(G478), .A2(n688), .ZN(n689) );
  XNOR2_X1 U744 ( .A(n690), .B(n689), .ZN(n691) );
  NOR2_X1 U745 ( .A1(n693), .A2(n691), .ZN(G63) );
  NAND2_X1 U746 ( .A1(n695), .A2(n694), .ZN(n703) );
  NAND2_X1 U747 ( .A1(n708), .A2(n696), .ZN(n700) );
  NAND2_X1 U748 ( .A1(G953), .A2(G224), .ZN(n697) );
  XNOR2_X1 U749 ( .A(KEYINPUT61), .B(n697), .ZN(n698) );
  NAND2_X1 U750 ( .A1(n698), .A2(G898), .ZN(n699) );
  NAND2_X1 U751 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U752 ( .A(n701), .B(KEYINPUT127), .ZN(n702) );
  XNOR2_X1 U753 ( .A(n703), .B(n702), .ZN(G69) );
  XNOR2_X1 U754 ( .A(n705), .B(n704), .ZN(n710) );
  INV_X1 U755 ( .A(n710), .ZN(n707) );
  XNOR2_X1 U756 ( .A(n707), .B(n706), .ZN(n709) );
  NAND2_X1 U757 ( .A1(n709), .A2(n708), .ZN(n714) );
  XNOR2_X1 U758 ( .A(G227), .B(n710), .ZN(n711) );
  NAND2_X1 U759 ( .A1(n711), .A2(G900), .ZN(n712) );
  NAND2_X1 U760 ( .A1(n712), .A2(G953), .ZN(n713) );
  NAND2_X1 U761 ( .A1(n714), .A2(n713), .ZN(G72) );
  XOR2_X1 U762 ( .A(n715), .B(G131), .Z(G33) );
  XNOR2_X1 U763 ( .A(n716), .B(G122), .ZN(G24) );
  XOR2_X1 U764 ( .A(G137), .B(n717), .Z(G39) );
  XNOR2_X1 U765 ( .A(G140), .B(n718), .ZN(G42) );
  XNOR2_X1 U766 ( .A(n719), .B(KEYINPUT37), .ZN(n720) );
  XNOR2_X1 U767 ( .A(n720), .B(KEYINPUT120), .ZN(n721) );
  XNOR2_X1 U768 ( .A(G125), .B(n721), .ZN(G27) );
  XNOR2_X1 U769 ( .A(G119), .B(n722), .ZN(G21) );
endmodule

