//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 1 1 1 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  OAI21_X1  g001(.A(G210), .B1(G237), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  OR3_X1    g003(.A1(new_n189), .A2(KEYINPUT65), .A3(G146), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT65), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n189), .A2(G146), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  AND2_X1   g009(.A1(KEYINPUT0), .A2(G128), .ZN(new_n196));
  NOR2_X1   g010(.A1(KEYINPUT0), .A2(G128), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n194), .A2(new_n192), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(new_n196), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G125), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT88), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n192), .A2(KEYINPUT1), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n195), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT68), .B1(new_n201), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT68), .ZN(new_n213));
  NOR4_X1   g027(.A1(new_n200), .A2(new_n213), .A3(KEYINPUT1), .A4(new_n210), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n209), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(G125), .ZN(new_n216));
  MUX2_X1   g030(.A(new_n206), .B(KEYINPUT88), .S(new_n216), .Z(new_n217));
  INV_X1    g031(.A(G953), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G224), .ZN(new_n219));
  XOR2_X1   g033(.A(new_n217), .B(new_n219), .Z(new_n220));
  XOR2_X1   g034(.A(G110), .B(G122), .Z(new_n221));
  XOR2_X1   g035(.A(new_n221), .B(KEYINPUT85), .Z(new_n222));
  INV_X1    g036(.A(KEYINPUT71), .ZN(new_n223));
  AND2_X1   g037(.A1(KEYINPUT70), .A2(G116), .ZN(new_n224));
  NOR2_X1   g038(.A1(KEYINPUT70), .A2(G116), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n223), .B(G119), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G119), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n228));
  INV_X1    g042(.A(G116), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(KEYINPUT70), .A2(G116), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n227), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT71), .B1(new_n229), .B2(G119), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n226), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT5), .ZN(new_n235));
  NOR3_X1   g049(.A1(new_n229), .A2(KEYINPUT5), .A3(G119), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n235), .A2(G113), .A3(new_n237), .ZN(new_n238));
  XOR2_X1   g052(.A(KEYINPUT2), .B(G113), .Z(new_n239));
  NAND2_X1  g053(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G104), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G107), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n241), .A2(G107), .ZN(new_n244));
  OAI21_X1  g058(.A(G101), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT3), .B1(new_n241), .B2(G107), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT3), .ZN(new_n247));
  INV_X1    g061(.A(G107), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n248), .A3(G104), .ZN(new_n249));
  INV_X1    g063(.A(G101), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n246), .A2(new_n249), .A3(new_n250), .A4(new_n242), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n245), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n238), .A2(new_n240), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT83), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n238), .A2(KEYINPUT83), .A3(new_n240), .A4(new_n253), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n234), .B(new_n239), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n251), .A2(KEYINPUT4), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n246), .A2(new_n249), .A3(new_n242), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G101), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n259), .B(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n256), .A2(new_n257), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT84), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n254), .A2(new_n255), .B1(new_n258), .B2(new_n262), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT84), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n267), .A3(new_n257), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n222), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  XOR2_X1   g083(.A(KEYINPUT87), .B(KEYINPUT6), .Z(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT6), .B1(new_n269), .B2(KEYINPUT86), .ZN(new_n272));
  INV_X1    g086(.A(new_n222), .ZN(new_n273));
  AND4_X1   g087(.A1(new_n267), .A2(new_n256), .A3(new_n257), .A4(new_n263), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n267), .B1(new_n266), .B2(new_n257), .ZN(new_n275));
  OAI211_X1 g089(.A(KEYINPUT86), .B(new_n273), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n264), .A2(new_n221), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n220), .B(new_n271), .C1(new_n272), .C2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT89), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT86), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n277), .B1(new_n269), .B2(KEYINPUT86), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n288), .A2(KEYINPUT89), .A3(new_n220), .A4(new_n271), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n282), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n219), .A2(KEYINPUT7), .ZN(new_n291));
  XOR2_X1   g105(.A(new_n217), .B(new_n291), .Z(new_n292));
  NAND2_X1  g106(.A1(new_n238), .A2(new_n240), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n252), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(KEYINPUT90), .A3(new_n254), .ZN(new_n295));
  XOR2_X1   g109(.A(new_n221), .B(KEYINPUT8), .Z(new_n296));
  OAI211_X1 g110(.A(new_n295), .B(new_n296), .C1(KEYINPUT90), .C2(new_n294), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n292), .A2(new_n297), .A3(new_n278), .ZN(new_n298));
  INV_X1    g112(.A(G902), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n188), .B1(new_n290), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n188), .ZN(new_n303));
  AOI211_X1 g117(.A(new_n303), .B(new_n300), .C1(new_n282), .C2(new_n289), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n187), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT91), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI211_X1 g121(.A(KEYINPUT91), .B(new_n187), .C1(new_n302), .C2(new_n304), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NOR3_X1   g123(.A1(new_n205), .A2(KEYINPUT16), .A3(G140), .ZN(new_n310));
  XNOR2_X1  g124(.A(G125), .B(G140), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n310), .B1(new_n311), .B2(KEYINPUT16), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(new_n191), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n227), .A2(G128), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n227), .A2(G128), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XOR2_X1   g131(.A(KEYINPUT24), .B(G110), .Z(new_n318));
  AOI21_X1  g132(.A(new_n313), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G110), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT23), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  NOR3_X1   g136(.A1(new_n227), .A2(KEYINPUT23), .A3(G128), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n314), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  XOR2_X1   g138(.A(new_n324), .B(KEYINPUT76), .Z(new_n325));
  OAI21_X1  g139(.A(new_n319), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n312), .A2(G146), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  XOR2_X1   g142(.A(KEYINPUT77), .B(G110), .Z(new_n329));
  OAI22_X1  g143(.A1(new_n324), .A2(new_n329), .B1(new_n317), .B2(new_n318), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n311), .A2(new_n191), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT22), .B(G137), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(KEYINPUT78), .ZN(new_n335));
  INV_X1    g149(.A(G221), .ZN(new_n336));
  INV_X1    g150(.A(G234), .ZN(new_n337));
  NOR3_X1   g151(.A1(new_n336), .A2(new_n337), .A3(G953), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n335), .B(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n333), .B(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  OAI211_X1 g155(.A(KEYINPUT79), .B(KEYINPUT25), .C1(new_n341), .C2(G902), .ZN(new_n342));
  OAI21_X1  g156(.A(G217), .B1(new_n337), .B2(G902), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n343), .B(KEYINPUT75), .ZN(new_n344));
  NAND2_X1  g158(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n345));
  OR2_X1    g159(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n340), .A2(new_n299), .A3(new_n345), .A4(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n342), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT80), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT80), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n342), .A2(new_n347), .A3(new_n350), .A4(new_n344), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n344), .A2(G902), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n340), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n349), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT11), .ZN(new_n355));
  INV_X1    g169(.A(G134), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n355), .B1(new_n356), .B2(G137), .ZN(new_n357));
  INV_X1    g171(.A(G137), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(KEYINPUT11), .A3(G134), .ZN(new_n359));
  INV_X1    g173(.A(G131), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n356), .A2(G137), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n357), .A2(new_n359), .A3(new_n360), .A4(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n362), .B(KEYINPUT66), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n357), .A2(new_n361), .A3(new_n359), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT67), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT67), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n357), .A2(new_n359), .A3(new_n366), .A4(new_n361), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n365), .A2(G131), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT72), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT72), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n363), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n203), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n361), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n356), .A2(G137), .ZN(new_n375));
  OAI21_X1  g189(.A(G131), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n215), .A2(new_n363), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT30), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT69), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n369), .A2(new_n204), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n215), .A2(KEYINPUT69), .A3(new_n363), .A4(new_n376), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  XOR2_X1   g199(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n380), .A2(new_n387), .A3(new_n258), .ZN(new_n388));
  INV_X1    g202(.A(new_n258), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n379), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(G101), .ZN(new_n392));
  INV_X1    g206(.A(G237), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT73), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT73), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G237), .ZN(new_n396));
  AOI21_X1  g210(.A(G953), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G210), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n392), .B(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n388), .A2(new_n390), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT31), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n385), .A2(new_n258), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT28), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n403), .B1(new_n379), .B2(new_n389), .ZN(new_n404));
  NOR4_X1   g218(.A1(new_n373), .A2(KEYINPUT28), .A3(new_n258), .A4(new_n378), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n402), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n399), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT31), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n388), .A2(new_n409), .A3(new_n390), .A4(new_n399), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n401), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(G472), .A2(G902), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n411), .A2(KEYINPUT32), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(KEYINPUT32), .B1(new_n411), .B2(new_n412), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT74), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n379), .A2(new_n389), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n399), .A2(KEYINPUT29), .ZN(new_n418));
  INV_X1    g232(.A(new_n404), .ZN(new_n419));
  INV_X1    g233(.A(new_n405), .ZN(new_n420));
  AOI211_X1 g234(.A(new_n417), .B(new_n418), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n416), .B1(new_n421), .B2(G902), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n417), .B1(new_n419), .B2(new_n420), .ZN(new_n423));
  INV_X1    g237(.A(new_n418), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(KEYINPUT74), .A3(new_n299), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n406), .A2(new_n399), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n388), .A2(new_n390), .A3(new_n407), .ZN(new_n429));
  AOI21_X1  g243(.A(KEYINPUT29), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(G472), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n354), .B1(new_n415), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G475), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT94), .ZN(new_n434));
  AOI21_X1  g248(.A(G143), .B1(new_n397), .B2(G214), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n397), .A2(G143), .A3(G214), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(KEYINPUT17), .A3(G131), .ZN(new_n439));
  INV_X1    g253(.A(new_n437), .ZN(new_n440));
  OAI21_X1  g254(.A(G131), .B1(new_n440), .B2(new_n435), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n436), .A2(new_n360), .A3(new_n437), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n313), .B(new_n439), .C1(new_n443), .C2(KEYINPUT17), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n311), .A2(new_n191), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT93), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n445), .B(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n331), .A2(KEYINPUT92), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n438), .A2(KEYINPUT18), .A3(G131), .ZN(new_n450));
  OR2_X1    g264(.A1(new_n445), .A2(new_n446), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n445), .A2(new_n446), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n451), .A2(KEYINPUT92), .A3(new_n331), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(KEYINPUT18), .A2(G131), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n436), .A2(new_n437), .A3(new_n454), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n449), .A2(new_n450), .A3(new_n453), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n444), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G113), .B(G122), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(new_n241), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n434), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n444), .A2(new_n456), .A3(KEYINPUT94), .A4(new_n459), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n457), .A2(new_n460), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n433), .B1(new_n465), .B2(new_n299), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n311), .B(KEYINPUT19), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n443), .B(new_n328), .C1(G146), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n456), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n460), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n463), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(new_n433), .A3(new_n299), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT20), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT95), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT20), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n472), .A2(new_n477), .A3(new_n433), .A4(new_n299), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  OR3_X1    g293(.A1(new_n473), .A2(KEYINPUT95), .A3(KEYINPUT20), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n466), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(G234), .A2(G237), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(G952), .A3(new_n218), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  XOR2_X1   g298(.A(KEYINPUT21), .B(G898), .Z(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n482), .A2(G902), .A3(G953), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n484), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(G128), .B(G143), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n356), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n491), .A2(KEYINPUT13), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n189), .A2(G128), .ZN(new_n494));
  OAI21_X1  g308(.A(G134), .B1(new_n494), .B2(KEYINPUT13), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT96), .B(G122), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(new_n229), .ZN(new_n497));
  INV_X1    g311(.A(G122), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n498), .B1(new_n230), .B2(new_n231), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  XOR2_X1   g314(.A(new_n500), .B(KEYINPUT97), .Z(new_n501));
  AND2_X1   g315(.A1(new_n501), .A2(new_n248), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n501), .A2(new_n248), .ZN(new_n503));
  OAI221_X1 g317(.A(new_n492), .B1(new_n493), .B2(new_n495), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n491), .B(G134), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n499), .B(KEYINPUT14), .ZN(new_n506));
  INV_X1    g320(.A(new_n497), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n248), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OR3_X1    g322(.A1(new_n502), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  XOR2_X1   g324(.A(KEYINPUT9), .B(G234), .Z(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(G217), .A3(new_n218), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n512), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n504), .A2(new_n509), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n299), .ZN(new_n517));
  INV_X1    g331(.A(G478), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(KEYINPUT15), .ZN(new_n519));
  XOR2_X1   g333(.A(new_n517), .B(new_n519), .Z(new_n520));
  NAND3_X1  g334(.A1(new_n481), .A2(new_n490), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(G469), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n262), .A2(new_n204), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n215), .A2(KEYINPUT10), .A3(new_n253), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n201), .A2(new_n211), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n213), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n201), .A2(KEYINPUT68), .A3(new_n211), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n208), .A2(new_n200), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n529), .A2(KEYINPUT81), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(KEYINPUT81), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n528), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n532), .A2(new_n253), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n523), .B(new_n524), .C1(new_n533), .C2(KEYINPUT10), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n370), .A2(new_n372), .ZN(new_n535));
  OR2_X1    g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XOR2_X1   g350(.A(G110), .B(G140), .Z(new_n537));
  INV_X1    g351(.A(G227), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(G953), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n537), .B(new_n539), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n215), .A2(new_n253), .ZN(new_n542));
  OR2_X1    g356(.A1(new_n542), .A2(KEYINPUT82), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(KEYINPUT82), .ZN(new_n544));
  AND2_X1   g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(KEYINPUT12), .B(new_n369), .C1(new_n545), .C2(new_n533), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n533), .B1(new_n543), .B2(new_n544), .ZN(new_n547));
  INV_X1    g361(.A(new_n535), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n546), .B1(KEYINPUT12), .B2(new_n549), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n541), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n534), .A2(new_n535), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n540), .B1(new_n536), .B2(new_n552), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n522), .B(new_n299), .C1(new_n551), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n541), .A2(new_n552), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n550), .A2(new_n536), .ZN(new_n556));
  OAI211_X1 g370(.A(G469), .B(new_n555), .C1(new_n556), .C2(new_n540), .ZN(new_n557));
  NAND2_X1  g371(.A1(G469), .A2(G902), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n554), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n336), .B1(new_n511), .B2(new_n299), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n521), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n309), .A2(new_n432), .A3(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(G101), .ZN(G3));
  NAND2_X1  g379(.A1(new_n411), .A2(new_n299), .ZN(new_n566));
  NAND2_X1  g380(.A1(KEYINPUT98), .A2(G472), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NOR3_X1   g383(.A1(new_n569), .A2(new_n354), .A3(new_n562), .ZN(new_n570));
  INV_X1    g384(.A(new_n187), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n290), .A2(new_n301), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n303), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n290), .A2(new_n188), .A3(new_n301), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n571), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n517), .A2(G478), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n518), .A2(new_n299), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  AND2_X1   g393(.A1(KEYINPUT99), .A2(KEYINPUT33), .ZN(new_n580));
  NOR2_X1   g394(.A1(KEYINPUT99), .A2(KEYINPUT33), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n516), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n580), .B1(new_n513), .B2(new_n515), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n577), .B(new_n579), .C1(new_n585), .C2(new_n518), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n481), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n570), .A2(new_n575), .A3(new_n490), .A4(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT34), .B(G104), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(KEYINPUT100), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n588), .B(new_n590), .ZN(G6));
  INV_X1    g405(.A(KEYINPUT102), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n478), .A2(KEYINPUT101), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n592), .B1(new_n478), .B2(KEYINPUT101), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n474), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n478), .A2(KEYINPUT101), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT102), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n598), .A2(KEYINPUT20), .A3(new_n473), .A4(new_n593), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n517), .B(new_n519), .ZN(new_n600));
  INV_X1    g414(.A(new_n466), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n596), .A2(new_n599), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(new_n489), .B(KEYINPUT103), .Z(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n575), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(KEYINPUT104), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT104), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n575), .A2(new_n603), .A3(new_n608), .A4(new_n605), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n570), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT35), .B(G107), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G9));
  INV_X1    g427(.A(new_n339), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(KEYINPUT36), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n333), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n352), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n349), .A2(new_n351), .A3(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n309), .A2(new_n563), .A3(new_n568), .A4(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT37), .B(G110), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT105), .B(KEYINPUT106), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G12));
  INV_X1    g437(.A(G900), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n484), .B1(new_n488), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n602), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n562), .B1(new_n415), .B2(new_n431), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n626), .A2(new_n575), .A3(new_n627), .A4(new_n618), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G128), .ZN(G30));
  NAND2_X1  g443(.A1(new_n573), .A2(new_n574), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT38), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n625), .B(KEYINPUT39), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n562), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT40), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n618), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n481), .A2(new_n571), .A3(new_n520), .ZN(new_n636));
  INV_X1    g450(.A(new_n390), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n407), .B1(new_n637), .B2(new_n417), .ZN(new_n638));
  OR2_X1    g452(.A1(new_n638), .A2(KEYINPUT107), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(KEYINPUT107), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n639), .A2(new_n400), .A3(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(G472), .B1(new_n641), .B2(G902), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n415), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n633), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n643), .B1(new_n644), .B2(KEYINPUT40), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n631), .A2(new_n635), .A3(new_n636), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G143), .ZN(G45));
  NOR3_X1   g461(.A1(new_n481), .A2(new_n586), .A3(new_n625), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n575), .A2(new_n648), .A3(new_n627), .A4(new_n618), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G146), .ZN(G48));
  NOR2_X1   g464(.A1(new_n551), .A2(new_n553), .ZN(new_n651));
  OAI21_X1  g465(.A(G469), .B1(new_n651), .B2(G902), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n652), .A2(new_n561), .A3(new_n554), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n432), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n654), .A2(new_n575), .A3(new_n490), .A4(new_n587), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT41), .B(G113), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G15));
  INV_X1    g471(.A(new_n654), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n658), .B1(new_n607), .B2(new_n609), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT108), .B(G116), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G18));
  NAND2_X1  g475(.A1(new_n415), .A2(new_n431), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n575), .A2(new_n662), .A3(new_n618), .A4(new_n653), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(new_n521), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(new_n227), .ZN(G21));
  AND2_X1   g479(.A1(new_n636), .A2(new_n630), .ZN(new_n666));
  INV_X1    g480(.A(new_n354), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n410), .B1(new_n423), .B2(new_n399), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n400), .A2(KEYINPUT31), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n412), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n670), .A2(KEYINPUT109), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(KEYINPUT109), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n566), .A2(G472), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n667), .A2(new_n671), .A3(new_n672), .A4(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n604), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n666), .A2(new_n653), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT110), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G122), .ZN(G24));
  AND4_X1   g492(.A1(new_n618), .A2(new_n671), .A3(new_n672), .A4(new_n673), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n575), .A2(new_n648), .A3(new_n679), .A4(new_n653), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G125), .ZN(G27));
  NOR2_X1   g495(.A1(new_n302), .A2(new_n304), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n432), .A2(new_n682), .A3(new_n187), .ZN(new_n683));
  INV_X1    g497(.A(new_n562), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n683), .A2(KEYINPUT42), .A3(new_n684), .A4(new_n648), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT42), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n432), .A2(new_n682), .A3(new_n187), .A4(new_n684), .ZN(new_n687));
  INV_X1    g501(.A(new_n648), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT111), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n685), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n690), .B1(new_n685), .B2(new_n689), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n360), .ZN(G33));
  NOR3_X1   g508(.A1(new_n687), .A2(new_n602), .A3(new_n625), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT112), .B(G134), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G36));
  INV_X1    g511(.A(new_n586), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n481), .ZN(new_n699));
  XOR2_X1   g513(.A(new_n699), .B(KEYINPUT43), .Z(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(KEYINPUT114), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n699), .B(KEYINPUT43), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT114), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n701), .A2(new_n569), .A3(new_n618), .A4(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n706));
  OR2_X1    g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n630), .A2(new_n571), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n555), .B1(new_n556), .B2(new_n540), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT45), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(G469), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n558), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT46), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n712), .A2(KEYINPUT113), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n554), .B1(new_n712), .B2(new_n713), .ZN(new_n715));
  AOI21_X1  g529(.A(KEYINPUT113), .B1(new_n712), .B2(new_n713), .ZN(new_n716));
  OR3_X1    g530(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n561), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n632), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n705), .A2(new_n706), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n707), .A2(new_n708), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G137), .ZN(G39));
  INV_X1    g536(.A(KEYINPUT47), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n718), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n717), .A2(KEYINPUT47), .A3(new_n561), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n708), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n727), .A2(new_n662), .A3(new_n667), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n726), .A2(new_n648), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G140), .ZN(G42));
  AND3_X1   g544(.A1(new_n708), .A2(new_n484), .A3(new_n653), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(new_n667), .A3(new_n643), .ZN(new_n732));
  INV_X1    g546(.A(new_n587), .ZN(new_n733));
  OAI211_X1 g547(.A(G952), .B(new_n218), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n674), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n700), .A2(new_n484), .A3(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT119), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n653), .A2(new_n571), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n631), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n737), .B(new_n740), .C1(new_n738), .C2(new_n739), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT50), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n700), .A2(new_n731), .A3(new_n679), .ZN(new_n744));
  INV_X1    g558(.A(new_n481), .ZN(new_n745));
  OR3_X1    g559(.A1(new_n732), .A2(new_n745), .A3(new_n698), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n743), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT51), .ZN(new_n749));
  INV_X1    g563(.A(new_n726), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n652), .A2(new_n554), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n560), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n736), .A2(new_n727), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n749), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n734), .B1(new_n748), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n752), .B(KEYINPUT118), .ZN(new_n757));
  AOI211_X1 g571(.A(new_n727), .B(new_n736), .C1(new_n750), .C2(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n749), .B1(new_n747), .B2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT116), .ZN(new_n760));
  INV_X1    g574(.A(new_n570), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n745), .A2(new_n520), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT91), .B1(new_n630), .B2(new_n187), .ZN(new_n763));
  INV_X1    g577(.A(new_n308), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n605), .B(new_n762), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT115), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n604), .B1(new_n307), .B2(new_n308), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n768), .A3(new_n762), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n761), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n309), .A2(new_n570), .A3(new_n587), .A4(new_n605), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n619), .A2(new_n771), .A3(new_n564), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n760), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  AND4_X1   g587(.A1(new_n768), .A2(new_n309), .A3(new_n605), .A4(new_n762), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n768), .B1(new_n767), .B2(new_n762), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n570), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n619), .A2(new_n771), .A3(new_n564), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(KEYINPUT116), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n773), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n664), .B1(new_n610), .B2(new_n654), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n676), .A2(new_n655), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n695), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n662), .A2(new_n520), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n596), .A2(new_n599), .A3(new_n601), .ZN(new_n788));
  OAI22_X1  g602(.A1(new_n733), .A2(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n562), .A2(new_n625), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n789), .A2(new_n618), .A3(new_n708), .A4(new_n790), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n785), .B(new_n791), .C1(new_n691), .C2(new_n692), .ZN(new_n792));
  INV_X1    g606(.A(new_n625), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n349), .A2(new_n351), .A3(new_n617), .A4(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n794), .B1(new_n415), .B2(new_n642), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n636), .A2(new_n795), .A3(new_n630), .A4(new_n684), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n628), .A2(new_n649), .A3(new_n680), .A4(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT52), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n792), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n779), .A2(new_n784), .A3(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n783), .B1(new_n773), .B2(new_n778), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT53), .B1(new_n803), .B2(new_n799), .ZN(new_n804));
  OAI21_X1  g618(.A(KEYINPUT54), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n800), .A2(new_n801), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n685), .A2(new_n689), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n798), .A2(new_n808), .A3(new_n695), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT117), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n810), .B1(new_n780), .B2(new_n782), .ZN(new_n811));
  NOR4_X1   g625(.A1(new_n659), .A2(new_n781), .A3(KEYINPUT117), .A4(new_n664), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n791), .A2(KEYINPUT53), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n779), .A2(new_n809), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n806), .A2(new_n807), .A3(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n756), .A2(new_n759), .A3(new_n805), .A4(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n700), .A2(new_n731), .A3(new_n432), .ZN(new_n818));
  XOR2_X1   g632(.A(new_n818), .B(KEYINPUT48), .Z(new_n819));
  NAND3_X1  g633(.A1(new_n737), .A2(new_n575), .A3(new_n653), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(KEYINPUT120), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n817), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(G952), .A2(G953), .ZN(new_n823));
  XOR2_X1   g637(.A(new_n751), .B(KEYINPUT49), .Z(new_n824));
  NOR4_X1   g638(.A1(new_n631), .A2(new_n824), .A3(new_n354), .A4(new_n560), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n187), .A3(new_n643), .ZN(new_n826));
  OAI22_X1  g640(.A1(new_n822), .A2(new_n823), .B1(new_n699), .B2(new_n826), .ZN(G75));
  AOI21_X1  g641(.A(new_n299), .B1(new_n806), .B2(new_n815), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(G210), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT56), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n286), .A2(new_n287), .B1(new_n269), .B2(new_n270), .ZN(new_n831));
  XOR2_X1   g645(.A(new_n831), .B(new_n220), .Z(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT55), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n829), .A2(new_n830), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n833), .B1(new_n829), .B2(new_n830), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n218), .A2(G952), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(G51));
  XOR2_X1   g651(.A(new_n558), .B(KEYINPUT57), .Z(new_n838));
  AND4_X1   g652(.A1(new_n779), .A2(new_n809), .A3(new_n813), .A4(new_n814), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n839), .A2(new_n804), .A3(KEYINPUT54), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n807), .B1(new_n806), .B2(new_n815), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n838), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n651), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n842), .A2(KEYINPUT121), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n845));
  INV_X1    g659(.A(new_n838), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT54), .B1(new_n839), .B2(new_n804), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n846), .B1(new_n847), .B2(new_n816), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n845), .B1(new_n848), .B2(new_n651), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n828), .A2(G469), .A3(new_n710), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n844), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n836), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(G54));
  NAND3_X1  g667(.A1(new_n828), .A2(KEYINPUT58), .A3(G475), .ZN(new_n854));
  INV_X1    g668(.A(new_n472), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n854), .A2(KEYINPUT122), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT122), .B1(new_n854), .B2(new_n855), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(G60));
  XNOR2_X1  g673(.A(new_n578), .B(KEYINPUT59), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n860), .B1(new_n805), .B2(new_n816), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n852), .B1(new_n861), .B2(new_n585), .ZN(new_n862));
  INV_X1    g676(.A(new_n585), .ZN(new_n863));
  AOI211_X1 g677(.A(new_n863), .B(new_n860), .C1(new_n847), .C2(new_n816), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n862), .A2(new_n864), .ZN(G63));
  NAND2_X1  g679(.A1(new_n806), .A2(new_n815), .ZN(new_n866));
  NAND2_X1  g680(.A1(G217), .A2(G902), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT60), .Z(new_n868));
  NAND3_X1  g682(.A1(new_n866), .A2(new_n616), .A3(new_n868), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n869), .A2(KEYINPUT123), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n866), .A2(new_n868), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n836), .B1(new_n871), .B2(new_n341), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n869), .A2(KEYINPUT123), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n870), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n870), .A2(KEYINPUT61), .A3(new_n872), .A4(new_n873), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(G66));
  INV_X1    g692(.A(G224), .ZN(new_n879));
  OAI21_X1  g693(.A(G953), .B1(new_n486), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n880), .B1(new_n803), .B2(G953), .ZN(new_n881));
  INV_X1    g695(.A(new_n831), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n882), .B1(G898), .B2(new_n218), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n881), .B(new_n883), .ZN(G69));
  NAND2_X1  g698(.A1(new_n624), .A2(G953), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n628), .A2(new_n649), .A3(new_n680), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT124), .Z(new_n887));
  NAND3_X1  g701(.A1(new_n721), .A2(new_n729), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n719), .A2(new_n432), .A3(new_n666), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n889), .B(new_n785), .C1(new_n692), .C2(new_n691), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n885), .B1(new_n891), .B2(G953), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n380), .A2(new_n387), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(new_n468), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(G953), .B1(new_n538), .B2(new_n624), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT127), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n683), .B(new_n633), .C1(new_n587), .C2(new_n762), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT126), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n721), .A2(new_n729), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n887), .A2(new_n646), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n902), .A2(KEYINPUT125), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n902), .A2(KEYINPUT125), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n901), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n901), .A2(new_n903), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n900), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n894), .B1(new_n907), .B2(new_n218), .ZN(new_n908));
  OR3_X1    g722(.A1(new_n895), .A2(new_n897), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n897), .B1(new_n895), .B2(new_n908), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(G72));
  NAND2_X1  g725(.A1(G472), .A2(G902), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT63), .Z(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n907), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n914), .B1(new_n915), .B2(new_n803), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n388), .A2(new_n390), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n399), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n852), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n891), .A2(new_n803), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n429), .B1(new_n920), .B2(new_n913), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n802), .A2(new_n804), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n918), .A2(new_n429), .A3(new_n913), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n919), .A2(new_n921), .A3(new_n924), .ZN(G57));
endmodule


