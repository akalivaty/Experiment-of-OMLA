//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1286, new_n1287, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1295, new_n1296, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g0005(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n206));
  NAND3_X1  g0006(.A1(new_n205), .A2(G50), .A3(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(KEYINPUT65), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n222), .A2(KEYINPUT65), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n213), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n212), .B(new_n216), .C1(new_n228), .C2(KEYINPUT1), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(G226), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n235), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n244), .B(new_n248), .ZN(G351));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n209), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT8), .B(G58), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G20), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n254), .A2(new_n256), .B1(G150), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n203), .ZN(new_n259));
  OAI21_X1  g0059(.A(G20), .B1(new_n259), .B2(G50), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n252), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G1), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(G13), .A3(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(new_n251), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n262), .A2(G20), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(G50), .A3(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G50), .B2(new_n263), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n261), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT9), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT71), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  AOI21_X1  g0073(.A(G1), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G1), .A3(G13), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(new_n276), .A3(G274), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(KEYINPUT69), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT69), .ZN(new_n279));
  INV_X1    g0079(.A(G274), .ZN(new_n280));
  INV_X1    g0080(.A(new_n209), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n280), .B1(new_n281), .B2(new_n275), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n279), .B1(new_n282), .B2(new_n274), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n278), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n262), .B1(G41), .B2(G45), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n276), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n284), .B1(G226), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT3), .B(G33), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(G222), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G77), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(G1698), .ZN(new_n293));
  INV_X1    g0093(.A(G223), .ZN(new_n294));
  OAI221_X1 g0094(.A(new_n291), .B1(new_n292), .B2(new_n289), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n288), .A2(G190), .A3(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n269), .A2(KEYINPUT9), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n288), .A2(new_n297), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n299), .B1(G200), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n271), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n271), .A2(new_n304), .A3(new_n298), .A4(new_n301), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G169), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n269), .B1(new_n300), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(G179), .B2(new_n300), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n265), .A2(G68), .A3(new_n266), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n311), .B(KEYINPUT73), .ZN(new_n312));
  INV_X1    g0112(.A(G68), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n257), .A2(G50), .B1(G20), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n210), .A2(G33), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n314), .B1(new_n292), .B2(new_n315), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n316), .A2(new_n251), .ZN(new_n317));
  OR2_X1    g0117(.A1(new_n317), .A2(KEYINPUT11), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n264), .A2(new_n313), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n319), .B(KEYINPUT12), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n317), .A2(KEYINPUT11), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n312), .A2(new_n318), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n289), .A2(G226), .A3(new_n290), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n289), .A2(G232), .A3(G1698), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G33), .A2(G97), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT72), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT72), .A4(new_n325), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(new_n296), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n277), .A2(KEYINPUT69), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n282), .A2(new_n279), .A3(new_n274), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n331), .A2(new_n332), .B1(G238), .B2(new_n287), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT13), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT13), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n330), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G179), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n335), .A2(new_n337), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT14), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(new_n341), .A3(G169), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n341), .B1(new_n340), .B2(G169), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n322), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n340), .A2(G200), .ZN(new_n346));
  INV_X1    g0146(.A(new_n322), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n335), .A2(G190), .A3(new_n337), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G58), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(new_n313), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n352), .A2(new_n203), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n353), .A2(G20), .B1(G159), .B2(new_n257), .ZN(new_n354));
  OR2_X1    g0154(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n355));
  NAND2_X1  g0155(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(G33), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT7), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(new_n360), .A3(new_n210), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G68), .ZN(new_n362));
  AOI21_X1  g0162(.A(G20), .B1(new_n357), .B2(new_n358), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(new_n360), .ZN(new_n364));
  OAI211_X1 g0164(.A(KEYINPUT16), .B(new_n354), .C1(new_n362), .C2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT16), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n360), .A2(G20), .ZN(new_n367));
  AOI21_X1  g0167(.A(G33), .B1(new_n355), .B2(new_n356), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT3), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G33), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n367), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n360), .B1(new_n289), .B2(G20), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n313), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n353), .A2(G20), .ZN(new_n375));
  INV_X1    g0175(.A(G159), .ZN(new_n376));
  INV_X1    g0176(.A(new_n257), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n366), .B1(new_n374), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n365), .A2(new_n379), .A3(new_n251), .ZN(new_n380));
  INV_X1    g0180(.A(new_n265), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n254), .A2(new_n266), .ZN(new_n382));
  OAI22_X1  g0182(.A1(new_n381), .A2(new_n382), .B1(new_n263), .B2(new_n254), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n331), .A2(new_n332), .B1(G232), .B2(new_n287), .ZN(new_n386));
  MUX2_X1   g0186(.A(G223), .B(G226), .S(G1698), .Z(new_n387));
  NAND3_X1  g0187(.A1(new_n387), .A2(new_n357), .A3(new_n358), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G33), .A2(G87), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n386), .B1(new_n390), .B2(new_n276), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G169), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n386), .B(G179), .C1(new_n390), .C2(new_n276), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n385), .A2(KEYINPUT18), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT75), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n385), .A2(KEYINPUT75), .A3(KEYINPUT18), .A4(new_n394), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n385), .A2(new_n394), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT18), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n397), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n287), .A2(G232), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(new_n278), .B2(new_n283), .ZN(new_n404));
  INV_X1    g0204(.A(G190), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n276), .B1(new_n388), .B2(new_n389), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n407), .B1(G200), .B2(new_n391), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n408), .A2(new_n380), .A3(new_n384), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT17), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n408), .A2(KEYINPUT17), .A3(new_n380), .A4(new_n384), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n402), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n266), .A2(G77), .ZN(new_n415));
  OAI22_X1  g0215(.A1(new_n381), .A2(new_n415), .B1(G77), .B2(new_n263), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n254), .A2(new_n257), .B1(G20), .B2(G77), .ZN(new_n417));
  XNOR2_X1  g0217(.A(KEYINPUT15), .B(G87), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n417), .B1(new_n315), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n416), .B1(new_n419), .B2(new_n251), .ZN(new_n420));
  XOR2_X1   g0220(.A(new_n420), .B(KEYINPUT70), .Z(new_n421));
  AOI21_X1  g0221(.A(new_n284), .B1(G244), .B2(new_n287), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n289), .A2(G232), .A3(new_n290), .ZN(new_n423));
  INV_X1    g0223(.A(G107), .ZN(new_n424));
  INV_X1    g0224(.A(G238), .ZN(new_n425));
  OAI221_X1 g0225(.A(new_n423), .B1(new_n424), .B2(new_n289), .C1(new_n293), .C2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n296), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(G200), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n422), .A2(G190), .A3(new_n427), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n421), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n428), .A2(new_n307), .ZN(new_n432));
  INV_X1    g0232(.A(G179), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n422), .A2(new_n433), .A3(new_n427), .ZN(new_n434));
  INV_X1    g0234(.A(new_n420), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n431), .A2(new_n436), .ZN(new_n437));
  NOR4_X1   g0237(.A1(new_n310), .A2(new_n350), .A3(new_n414), .A4(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT81), .ZN(new_n439));
  INV_X1    g0239(.A(G244), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(G1698), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n357), .A2(new_n358), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT4), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n358), .A2(new_n370), .A3(G250), .A4(G1698), .ZN(new_n445));
  AND2_X1   g0245(.A1(KEYINPUT4), .A2(G244), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n358), .A2(new_n370), .A3(new_n446), .A4(new_n290), .ZN(new_n447));
  NAND2_X1  g0247(.A1(G33), .A2(G283), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT78), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT78), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(G33), .A3(G283), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n445), .A2(new_n447), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT79), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n444), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n454), .B1(new_n444), .B2(new_n453), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n296), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(KEYINPUT5), .A2(G41), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(KEYINPUT5), .A2(G41), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n273), .A2(G1), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n296), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G257), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n262), .A2(G45), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n465), .B1(new_n459), .B2(new_n460), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n282), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(G179), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n457), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n424), .B1(new_n372), .B2(new_n373), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT6), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n472), .A2(new_n220), .A3(G107), .ZN(new_n473));
  XNOR2_X1  g0273(.A(G97), .B(G107), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n473), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  OAI22_X1  g0275(.A1(new_n475), .A2(new_n210), .B1(new_n292), .B2(new_n377), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n251), .B1(new_n471), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n262), .A2(G33), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n252), .A2(KEYINPUT76), .A3(new_n263), .A4(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n263), .A2(new_n478), .A3(new_n209), .A4(new_n250), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT76), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G97), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n264), .A2(G97), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT77), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n220), .B1(new_n479), .B2(new_n482), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT77), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n488), .A2(new_n489), .A3(new_n485), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n477), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n470), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n468), .ZN(new_n493));
  AOI21_X1  g0293(.A(G169), .B1(new_n457), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n439), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n484), .A2(KEYINPUT77), .A3(new_n486), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n489), .B1(new_n488), .B2(new_n485), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n477), .A2(new_n498), .B1(new_n457), .B2(new_n469), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n444), .A2(new_n453), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT79), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n444), .A2(new_n453), .A3(new_n454), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n276), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n307), .B1(new_n503), .B2(new_n468), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n499), .A2(KEYINPUT81), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n495), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(G200), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n507), .B1(new_n457), .B2(new_n493), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT80), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n457), .A2(G190), .A3(new_n493), .ZN(new_n511));
  XNOR2_X1  g0311(.A(KEYINPUT74), .B(KEYINPUT3), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n371), .B1(new_n512), .B2(new_n255), .ZN(new_n513));
  INV_X1    g0313(.A(new_n367), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n373), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G107), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n474), .A2(new_n472), .ZN(new_n517));
  INV_X1    g0317(.A(new_n473), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n519), .A2(G20), .B1(G77), .B2(new_n257), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n252), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n521), .B1(new_n497), .B2(new_n496), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n509), .A2(new_n510), .A3(new_n511), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n511), .A2(new_n522), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT80), .B1(new_n524), .B2(new_n508), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n506), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n479), .A2(new_n482), .A3(G87), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT82), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n479), .A2(new_n482), .A3(KEYINPUT82), .A4(G87), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(G238), .A2(G1698), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n440), .B2(G1698), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n533), .A2(new_n357), .A3(new_n358), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G116), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n276), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n462), .A2(new_n219), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n282), .A2(new_n462), .B1(new_n537), .B2(new_n276), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(G200), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n535), .ZN(new_n541));
  INV_X1    g0341(.A(new_n358), .ZN(new_n542));
  AND2_X1   g0342(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n543));
  NOR2_X1   g0343(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n542), .B1(new_n545), .B2(G33), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n541), .B1(new_n546), .B2(new_n533), .ZN(new_n547));
  OAI211_X1 g0347(.A(G190), .B(new_n538), .C1(new_n547), .C2(new_n276), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n357), .A2(new_n210), .A3(G68), .A4(new_n358), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT19), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n256), .A2(new_n550), .A3(G97), .ZN(new_n551));
  NOR2_X1   g0351(.A1(G97), .A2(G107), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n552), .A2(new_n218), .B1(new_n325), .B2(new_n210), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n551), .B1(new_n553), .B2(new_n550), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n555), .A2(new_n251), .B1(new_n264), .B2(new_n418), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n531), .A2(new_n540), .A3(new_n548), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n251), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n418), .A2(new_n264), .ZN(new_n559));
  INV_X1    g0359(.A(new_n418), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n479), .A2(new_n482), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n558), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n307), .B1(new_n536), .B2(new_n539), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n433), .B(new_n538), .C1(new_n547), .C2(new_n276), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n557), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(G257), .A2(G1698), .ZN(new_n567));
  INV_X1    g0367(.A(G264), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n567), .B1(new_n568), .B2(G1698), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n569), .A2(new_n357), .A3(new_n358), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n358), .A2(new_n370), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G303), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n296), .ZN(new_n574));
  INV_X1    g0374(.A(new_n460), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n462), .B1(new_n575), .B2(new_n458), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n576), .A2(G270), .A3(new_n276), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n467), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n307), .B1(new_n574), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n210), .B1(new_n220), .B2(G33), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n452), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(G116), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G20), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n582), .A2(KEYINPUT20), .A3(new_n251), .A4(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT20), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n580), .B1(new_n451), .B2(new_n449), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n251), .A2(new_n584), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n480), .A2(G116), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n263), .A2(new_n583), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT21), .B1(new_n579), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n585), .A2(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n574), .A2(G179), .A3(new_n578), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT21), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n598), .A2(new_n307), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n276), .B1(new_n570), .B2(new_n572), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n467), .A2(new_n577), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n596), .B1(new_n597), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n595), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n600), .A2(new_n601), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(G190), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n606), .B(new_n596), .C1(new_n507), .C2(new_n605), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n566), .A2(new_n604), .A3(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(G250), .A2(G1698), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n609), .B1(new_n221), .B2(G1698), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n610), .A2(new_n357), .A3(new_n358), .ZN(new_n611));
  NAND2_X1  g0411(.A1(G33), .A2(G294), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n276), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n467), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n466), .A2(new_n568), .A3(new_n296), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n433), .ZN(new_n617));
  INV_X1    g0417(.A(new_n616), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n307), .ZN(new_n619));
  OAI21_X1  g0419(.A(KEYINPUT23), .B1(new_n210), .B2(G107), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT23), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n621), .A2(new_n424), .A3(G20), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n620), .B(new_n622), .C1(new_n583), .C2(new_n315), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT83), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n256), .A2(G116), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n626), .A2(KEYINPUT83), .A3(new_n622), .A4(new_n620), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT22), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n629), .A2(new_n218), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n357), .A2(new_n210), .A3(new_n358), .A4(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n210), .A2(G87), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n629), .B1(new_n571), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT24), .B1(new_n628), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n634), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT24), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n625), .A2(new_n627), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n252), .B1(new_n635), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n479), .A2(new_n482), .A3(G107), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n263), .A2(G107), .ZN(new_n642));
  XNOR2_X1  g0442(.A(new_n642), .B(KEYINPUT25), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n617), .B(new_n619), .C1(new_n640), .C2(new_n644), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n628), .A2(KEYINPUT24), .A3(new_n634), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n637), .B1(new_n636), .B2(new_n638), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n251), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n644), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n611), .A2(new_n612), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n296), .ZN(new_n651));
  INV_X1    g0451(.A(new_n615), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n651), .A2(new_n405), .A3(new_n467), .A4(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(new_n616), .B2(G200), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n648), .A2(new_n649), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n645), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n608), .A2(new_n656), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n438), .A2(new_n526), .A3(new_n657), .ZN(G372));
  NAND2_X1  g0458(.A1(new_n566), .A2(new_n655), .ZN(new_n659));
  INV_X1    g0459(.A(new_n603), .ZN(new_n660));
  OAI21_X1  g0460(.A(G169), .B1(new_n600), .B2(new_n601), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n598), .B1(new_n661), .B2(new_n596), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n660), .A2(KEYINPUT84), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT84), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n595), .B2(new_n603), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n659), .B1(new_n666), .B2(new_n645), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n492), .A2(new_n439), .A3(new_n494), .ZN(new_n668));
  AOI21_X1  g0468(.A(KEYINPUT81), .B1(new_n499), .B2(new_n504), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n525), .A2(new_n523), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n566), .B1(new_n668), .B2(new_n669), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(KEYINPUT26), .ZN(new_n674));
  INV_X1    g0474(.A(new_n565), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n557), .A2(new_n565), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n492), .A2(new_n676), .A3(new_n494), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT26), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n675), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n672), .A2(new_n674), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n438), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n309), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n401), .A2(new_n395), .ZN(new_n683));
  OAI21_X1  g0483(.A(KEYINPUT14), .B1(new_n338), .B2(new_n307), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n684), .A2(new_n339), .A3(new_n342), .ZN(new_n685));
  INV_X1    g0485(.A(new_n436), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n685), .A2(new_n322), .B1(new_n349), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n411), .A2(new_n412), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n683), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n682), .B1(new_n689), .B2(new_n306), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n681), .A2(new_n690), .ZN(G369));
  INV_X1    g0491(.A(G13), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G1), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT27), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(new_n694), .A3(new_n210), .ZN(new_n695));
  XOR2_X1   g0495(.A(new_n695), .B(KEYINPUT85), .Z(new_n696));
  INV_X1    g0496(.A(G213), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n693), .A2(new_n210), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n697), .B1(new_n698), .B2(KEYINPUT27), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT86), .ZN(new_n701));
  INV_X1    g0501(.A(G343), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n594), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT87), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n705), .A2(new_n604), .A3(new_n607), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n666), .B2(new_n705), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n707), .A2(G330), .ZN(new_n708));
  INV_X1    g0508(.A(new_n656), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n648), .A2(new_n649), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n703), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n709), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n645), .B2(new_n712), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n708), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n703), .A2(new_n604), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n709), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n645), .B2(new_n703), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n715), .A2(new_n719), .ZN(G399));
  INV_X1    g0520(.A(new_n214), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G41), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n552), .A2(new_n218), .A3(new_n583), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n722), .A2(new_n262), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n724), .B1(new_n208), .B2(new_n722), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT88), .ZN(new_n726));
  XOR2_X1   g0526(.A(new_n726), .B(KEYINPUT28), .Z(new_n727));
  NAND4_X1  g0527(.A1(new_n670), .A2(new_n657), .A3(new_n671), .A4(new_n712), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n536), .A2(new_n539), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n613), .A2(new_n615), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n597), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT30), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(KEYINPUT89), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n732), .A2(new_n493), .A3(new_n457), .A4(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n457), .A2(new_n493), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n729), .A2(new_n605), .A3(G179), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n736), .A2(new_n618), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n736), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n734), .B1(new_n740), .B2(new_n732), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n703), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT31), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI211_X1 g0544(.A(KEYINPUT31), .B(new_n703), .C1(new_n739), .C2(new_n741), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n728), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n746), .A2(G330), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n680), .A2(new_n712), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT90), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT29), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n680), .A2(KEYINPUT90), .A3(new_n712), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n673), .A2(KEYINPUT91), .A3(new_n678), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT91), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n676), .B1(new_n495), .B2(new_n505), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n755), .B1(new_n756), .B2(KEYINPUT26), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n677), .A2(KEYINPUT26), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n754), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n659), .B1(new_n645), .B2(new_n604), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n675), .B1(new_n526), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n703), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(KEYINPUT29), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n747), .B1(new_n753), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n727), .B1(new_n764), .B2(G1), .ZN(G364));
  NOR2_X1   g0565(.A1(new_n692), .A2(G20), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n262), .B1(new_n766), .B2(G45), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n722), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n708), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(G330), .B2(new_n707), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n721), .A2(new_n571), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT92), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n772), .B1(new_n773), .B2(G355), .ZN(new_n774));
  AND2_X1   g0574(.A1(G355), .A2(new_n773), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n774), .A2(new_n775), .B1(G116), .B2(new_n214), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n546), .A2(new_n721), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n778), .B1(new_n273), .B2(new_n208), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n248), .A2(G45), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n776), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G13), .A2(G33), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G20), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n209), .B1(G20), .B2(new_n307), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n769), .B1(new_n781), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(G20), .A2(G179), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT93), .Z(new_n790));
  NAND3_X1  g0590(.A1(new_n790), .A2(new_n405), .A3(G200), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT96), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(KEYINPUT33), .B(G317), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR4_X1   g0598(.A1(new_n210), .A2(new_n405), .A3(new_n507), .A4(G179), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n289), .B1(new_n799), .B2(G303), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT98), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n790), .A2(new_n405), .A3(new_n507), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n801), .B1(G311), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n405), .A2(G20), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT95), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n807), .A2(G179), .A3(G200), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n405), .A2(G179), .A3(G200), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n210), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n808), .A2(G329), .B1(G294), .B2(new_n811), .ZN(new_n812));
  NOR3_X1   g0612(.A1(new_n807), .A2(G179), .A3(new_n507), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G283), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n790), .A2(G190), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(G200), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n790), .A2(G190), .A3(G200), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(KEYINPUT97), .B(G326), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G322), .A2(new_n817), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n798), .A2(new_n804), .A3(new_n815), .A4(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n799), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n289), .B1(new_n823), .B2(new_n218), .ZN(new_n824));
  INV_X1    g0624(.A(new_n813), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(new_n424), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n824), .B(new_n826), .C1(G97), .C2(new_n811), .ZN(new_n827));
  INV_X1    g0627(.A(new_n817), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n828), .A2(new_n351), .B1(new_n292), .B2(new_n802), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(KEYINPUT94), .ZN(new_n830));
  INV_X1    g0630(.A(new_n808), .ZN(new_n831));
  OAI21_X1  g0631(.A(KEYINPUT32), .B1(new_n831), .B2(new_n376), .ZN(new_n832));
  NOR3_X1   g0632(.A1(new_n831), .A2(KEYINPUT32), .A3(new_n376), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(G50), .B2(new_n819), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n827), .A2(new_n830), .A3(new_n832), .A4(new_n834), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n829), .A2(KEYINPUT94), .B1(new_n795), .B2(new_n313), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n822), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n788), .B1(new_n837), .B2(new_n785), .ZN(new_n838));
  INV_X1    g0638(.A(new_n784), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n838), .B1(new_n707), .B2(new_n839), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n771), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G396));
  NAND2_X1  g0642(.A1(new_n703), .A2(new_n435), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n431), .A2(new_n843), .A3(new_n436), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(KEYINPUT99), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n686), .A2(new_n703), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT99), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n431), .A2(new_n843), .A3(new_n436), .A4(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n750), .A2(new_n752), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n845), .A2(new_n848), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n680), .A2(new_n712), .A3(new_n852), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NOR3_X1   g0654(.A1(new_n854), .A2(KEYINPUT100), .A3(new_n747), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n769), .ZN(new_n857));
  OAI21_X1  g0657(.A(KEYINPUT100), .B1(new_n854), .B2(new_n747), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n854), .A2(new_n747), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n856), .A2(new_n857), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n785), .ZN(new_n861));
  AOI22_X1  g0661(.A1(G137), .A2(new_n819), .B1(new_n803), .B2(G159), .ZN(new_n862));
  INV_X1    g0662(.A(G143), .ZN(new_n863));
  INV_X1    g0663(.A(G150), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n862), .B1(new_n863), .B2(new_n828), .C1(new_n795), .C2(new_n864), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT34), .ZN(new_n866));
  INV_X1    g0666(.A(G50), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n546), .B1(new_n351), .B2(new_n810), .C1(new_n823), .C2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n825), .A2(new_n313), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n868), .B(new_n869), .C1(G132), .C2(new_n808), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n571), .B1(new_n220), .B2(new_n810), .C1(new_n823), .C2(new_n424), .ZN(new_n872));
  INV_X1    g0672(.A(G311), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n831), .A2(new_n873), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n872), .B(new_n874), .C1(G87), .C2(new_n813), .ZN(new_n875));
  INV_X1    g0675(.A(G303), .ZN(new_n876));
  OAI22_X1  g0676(.A1(new_n583), .A2(new_n802), .B1(new_n818), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(G294), .B2(new_n817), .ZN(new_n878));
  INV_X1    g0678(.A(G283), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n875), .B(new_n878), .C1(new_n879), .C2(new_n795), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n861), .B1(new_n871), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n785), .A2(new_n782), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n857), .B(new_n881), .C1(new_n292), .C2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n783), .B2(new_n849), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n860), .A2(new_n884), .ZN(G384));
  OR2_X1    g0685(.A1(new_n519), .A2(KEYINPUT35), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n519), .A2(KEYINPUT35), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n886), .A2(G116), .A3(new_n211), .A4(new_n887), .ZN(new_n888));
  XOR2_X1   g0688(.A(KEYINPUT101), .B(KEYINPUT36), .Z(new_n889));
  XNOR2_X1  g0689(.A(new_n888), .B(new_n889), .ZN(new_n890));
  OR3_X1    g0690(.A1(new_n207), .A2(new_n292), .A3(new_n352), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n867), .A2(G68), .ZN(new_n892));
  AOI211_X1 g0692(.A(new_n262), .B(G13), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(G330), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n365), .A2(new_n251), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n354), .B1(new_n362), .B2(new_n364), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n366), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n383), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n409), .B1(new_n899), .B2(new_n701), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n392), .A2(new_n393), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT37), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n700), .B(KEYINPUT86), .Z(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n385), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT37), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n905), .A2(new_n399), .A3(new_n409), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT18), .B1(new_n385), .B2(new_n394), .ZN(new_n909));
  AOI221_X4 g0709(.A(new_n400), .B1(new_n392), .B2(new_n393), .C1(new_n380), .C2(new_n384), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n909), .B1(new_n910), .B2(KEYINPUT75), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n688), .B1(new_n911), .B2(new_n397), .ZN(new_n912));
  INV_X1    g0712(.A(new_n899), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n904), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n908), .B(KEYINPUT38), .C1(new_n912), .C2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT103), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n914), .B1(new_n402), .B2(new_n413), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n919), .A2(KEYINPUT103), .A3(KEYINPUT38), .A4(new_n908), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT38), .ZN(new_n921));
  INV_X1    g0721(.A(new_n908), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n921), .B1(new_n922), .B2(new_n918), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n917), .A2(new_n920), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n746), .A2(new_n849), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n703), .A2(new_n322), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n345), .A2(new_n349), .A3(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n349), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n322), .B(new_n703), .C1(new_n685), .C2(new_n928), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n925), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT40), .B1(new_n924), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n905), .A2(new_n399), .A3(new_n409), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(new_n906), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n905), .B1(new_n413), .B2(new_n683), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n921), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n937), .A2(new_n915), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n927), .A2(new_n929), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n939), .A2(new_n746), .A3(KEYINPUT40), .A4(new_n849), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n933), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n438), .A2(new_n746), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT104), .Z(new_n944));
  AOI21_X1  g0744(.A(new_n895), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n942), .B2(new_n944), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n683), .A2(new_n904), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n436), .A2(new_n703), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT102), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n930), .B1(new_n853), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n947), .B1(new_n950), .B2(new_n924), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n937), .A2(new_n915), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n952), .A2(KEYINPUT39), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(KEYINPUT39), .B2(new_n924), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n685), .A2(new_n322), .A3(new_n712), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n951), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n753), .A2(new_n438), .A3(new_n763), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n690), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n956), .B(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n946), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n262), .B2(new_n766), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n946), .A2(new_n959), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n894), .B1(new_n961), .B2(new_n962), .ZN(G367));
  NOR2_X1   g0763(.A1(new_n239), .A2(new_n778), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n786), .B1(new_n214), .B2(new_n418), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n769), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AOI22_X1  g0766(.A1(G303), .A2(new_n817), .B1(new_n803), .B2(G283), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n873), .B2(new_n818), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n825), .A2(new_n220), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n799), .A2(G116), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT46), .Z(new_n971));
  NOR2_X1   g0771(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n546), .B1(G107), .B2(new_n811), .ZN(new_n973));
  INV_X1    g0773(.A(G317), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n972), .B(new_n973), .C1(new_n974), .C2(new_n831), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n968), .B(new_n975), .C1(G294), .C2(new_n796), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n808), .A2(G137), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n813), .A2(G77), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n811), .A2(G68), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n571), .B1(new_n799), .B2(G58), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n977), .A2(new_n978), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  AOI22_X1  g0781(.A1(G50), .A2(new_n803), .B1(new_n819), .B2(G143), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n864), .B2(new_n828), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n981), .B(new_n983), .C1(G159), .C2(new_n796), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n976), .A2(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT47), .Z(new_n986));
  AOI21_X1  g0786(.A(new_n966), .B1(new_n986), .B2(new_n785), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n531), .A2(new_n556), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n703), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n566), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n565), .B2(new_n989), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n987), .B1(new_n839), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n526), .B1(new_n522), .B2(new_n712), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n703), .A2(new_n504), .A3(new_n499), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n717), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT42), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n994), .A2(new_n995), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n670), .B1(new_n999), .B2(new_n645), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n998), .B1(new_n1000), .B2(new_n712), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n996), .A2(new_n997), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1002), .A2(KEYINPUT105), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT105), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(new_n996), .B2(new_n997), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1001), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(KEYINPUT106), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT106), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1010), .A2(new_n1011), .A3(new_n1007), .A4(new_n1001), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n715), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n994), .A2(new_n995), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1006), .A2(new_n1008), .A3(new_n1018), .ZN(new_n1019));
  AND3_X1   g0819(.A1(new_n1013), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1017), .B1(new_n1013), .B2(new_n1019), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n994), .A2(new_n718), .A3(new_n995), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT44), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT45), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1026), .B(new_n718), .C1(new_n994), .C2(new_n995), .ZN(new_n1027));
  AOI21_X1  g0827(.A(KEYINPUT45), .B1(new_n1015), .B2(new_n719), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n1014), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1025), .B(new_n715), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n717), .B1(new_n714), .B2(new_n716), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n708), .B(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n764), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n764), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n722), .B(KEYINPUT41), .Z(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n768), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n993), .B1(new_n1022), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(G387));
  AOI22_X1  g0842(.A1(new_n772), .A2(new_n723), .B1(new_n424), .B2(new_n721), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n235), .A2(new_n273), .ZN(new_n1044));
  AOI211_X1 g0844(.A(G45), .B(new_n723), .C1(G68), .C2(G77), .ZN(new_n1045));
  AND3_X1   g0845(.A1(new_n254), .A2(KEYINPUT50), .A3(new_n867), .ZN(new_n1046));
  AOI21_X1  g0846(.A(KEYINPUT50), .B1(new_n254), .B2(new_n867), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n777), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1043), .B1(new_n1044), .B2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1050), .A2(KEYINPUT107), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(KEYINPUT107), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n786), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n769), .B1(new_n1051), .B2(new_n1053), .C1(new_n714), .C2(new_n839), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n811), .A2(new_n560), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n799), .A2(G77), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1055), .A2(new_n546), .A3(new_n1056), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1057), .B(new_n969), .C1(G150), .C2(new_n808), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n828), .A2(new_n867), .B1(new_n376), .B2(new_n818), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G68), .B2(new_n803), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1058), .B(new_n1060), .C1(new_n253), .C2(new_n795), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G303), .A2(new_n803), .B1(new_n819), .B2(G322), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n974), .B2(new_n828), .C1(new_n795), .C2(new_n873), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT48), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n811), .A2(G283), .B1(new_n799), .B2(G294), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT108), .Z(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(KEYINPUT49), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n359), .B1(new_n825), .B2(new_n583), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n808), .B2(new_n820), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1069), .A2(KEYINPUT49), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1061), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1054), .B1(new_n1075), .B2(new_n785), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n1034), .B2(new_n768), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1035), .A2(new_n722), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1034), .A2(new_n764), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1077), .B1(new_n1078), .B2(new_n1079), .ZN(G393));
  INV_X1    g0880(.A(KEYINPUT109), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1030), .A2(new_n1081), .A3(new_n1031), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1029), .A2(KEYINPUT109), .A3(new_n1014), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n767), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1015), .A2(new_n839), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT110), .Z(new_n1086));
  OAI221_X1 g0886(.A(new_n786), .B1(new_n220), .B2(new_n214), .C1(new_n243), .C2(new_n778), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1087), .A2(KEYINPUT111), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(KEYINPUT111), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1088), .A2(new_n769), .A3(new_n1089), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n546), .B1(new_n292), .B2(new_n810), .C1(new_n823), .C2(new_n313), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n218), .A2(new_n825), .B1(new_n831), .B2(new_n863), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1091), .B(new_n1092), .C1(new_n254), .C2(new_n803), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n828), .A2(new_n376), .B1(new_n864), .B2(new_n818), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT51), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1093), .B(new_n1095), .C1(new_n867), .C2(new_n795), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n1096), .A2(KEYINPUT112), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n826), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n808), .A2(G322), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n811), .A2(G116), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n289), .B1(new_n799), .B2(G283), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G294), .B2(new_n803), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(G311), .A2(new_n817), .B1(new_n819), .B2(G317), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1104), .B(new_n1105), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1103), .B(new_n1106), .C1(new_n876), .C2(new_n795), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1096), .A2(KEYINPUT112), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1097), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1090), .B1(new_n1109), .B2(new_n785), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1084), .B1(new_n1086), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1082), .A2(new_n1035), .A3(new_n1083), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1112), .B(new_n722), .C1(new_n1035), .C2(new_n1032), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1111), .A2(new_n1113), .ZN(G390));
  NAND2_X1  g0914(.A1(new_n924), .A2(KEYINPUT39), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n953), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n955), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1115), .B(new_n1116), .C1(new_n1117), .C2(new_n950), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n939), .A2(new_n746), .A3(G330), .A4(new_n849), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n938), .A2(new_n1117), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n948), .B1(new_n762), .B2(new_n852), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT114), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n939), .B(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1120), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1118), .A2(new_n1119), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1119), .B1(new_n1118), .B2(new_n1124), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1125), .A2(new_n1126), .A3(new_n767), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n954), .A2(new_n782), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n571), .B1(new_n292), .B2(new_n810), .C1(new_n823), .C2(new_n218), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1129), .B(new_n869), .C1(G294), .C2(new_n808), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n828), .A2(new_n583), .B1(new_n879), .B2(new_n818), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(G97), .B2(new_n803), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1130), .B(new_n1132), .C1(new_n424), .C2(new_n795), .ZN(new_n1133));
  INV_X1    g0933(.A(G137), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n795), .A2(new_n1134), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n289), .B1(new_n810), .B2(new_n376), .C1(new_n825), .C2(new_n867), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(G125), .B2(new_n808), .ZN(new_n1137));
  INV_X1    g0937(.A(G132), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT54), .B(G143), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n828), .A2(new_n1138), .B1(new_n802), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(G128), .B2(new_n819), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n799), .A2(G150), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT117), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT53), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1137), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1133), .B1(new_n1135), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n861), .B1(new_n1146), .B2(KEYINPUT118), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(KEYINPUT118), .B2(new_n1146), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n857), .B1(new_n253), .B2(new_n882), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1128), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(KEYINPUT119), .B1(new_n1127), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT119), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n950), .A2(new_n1117), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1124), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1119), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1118), .A2(new_n1119), .A3(new_n1124), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1153), .B(new_n1150), .C1(new_n1160), .C2(new_n767), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1152), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT120), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n722), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n438), .A2(new_n747), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n957), .A2(new_n690), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(KEYINPUT115), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n939), .B(KEYINPUT114), .ZN(new_n1168));
  AND4_X1   g0968(.A1(new_n671), .A2(new_n670), .A3(new_n657), .A4(new_n712), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n744), .A2(new_n745), .ZN(new_n1170));
  OAI211_X1 g0970(.A(G330), .B(new_n849), .C1(new_n1169), .C2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1121), .B(new_n1119), .C1(new_n1168), .C2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1171), .A2(new_n930), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n1119), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n853), .A2(new_n949), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n1175), .A2(KEYINPUT116), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(KEYINPUT116), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1173), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT115), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n957), .A2(new_n1180), .A3(new_n690), .A4(new_n1165), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1167), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1164), .B1(new_n1160), .B2(new_n1182), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n1167), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n1162), .A2(new_n1163), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1163), .B1(new_n1162), .B2(new_n1187), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1188), .A2(new_n1189), .ZN(G378));
  XNOR2_X1  g0990(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n701), .A2(new_n269), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n306), .A2(new_n309), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1194), .B1(new_n306), .B2(new_n309), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1192), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1197), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1199), .A2(new_n1195), .A3(new_n1191), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(G330), .B1(new_n938), .B2(new_n940), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1202), .B1(new_n932), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n932), .A2(new_n1203), .A3(new_n1202), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n956), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1203), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n933), .A2(new_n1208), .A3(new_n1201), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1154), .A2(new_n1117), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1209), .A2(new_n1210), .A3(new_n1204), .A4(new_n951), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1207), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1202), .A2(new_n782), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n882), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n769), .B1(new_n1214), .B2(G50), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n359), .A2(new_n272), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n813), .A2(G58), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1217), .A2(new_n979), .A3(new_n1056), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1216), .B(new_n1218), .C1(G283), .C2(new_n808), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n828), .A2(new_n424), .B1(new_n583), .B2(new_n818), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n560), .B2(new_n803), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1219), .B(new_n1221), .C1(new_n220), .C2(new_n795), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT58), .ZN(new_n1223));
  AOI21_X1  g1023(.A(G50), .B1(new_n255), .B2(new_n272), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1222), .A2(new_n1223), .B1(new_n1216), .B2(new_n1224), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(G128), .A2(new_n817), .B1(new_n803), .B2(G137), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n823), .A2(new_n1139), .B1(new_n864), .B2(new_n810), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n819), .B2(G125), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1226), .B(new_n1228), .C1(new_n795), .C2(new_n1138), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1229), .A2(KEYINPUT59), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(KEYINPUT59), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n255), .B(new_n272), .C1(new_n825), .C2(new_n376), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(G124), .B2(new_n808), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1225), .B1(new_n1223), .B2(new_n1222), .C1(new_n1230), .C2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1215), .B1(new_n1235), .B2(new_n785), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1212), .A2(new_n768), .B1(new_n1213), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT121), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1167), .A2(new_n1238), .A3(new_n1181), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1238), .B1(new_n1167), .B2(new_n1181), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n1239), .A2(new_n1240), .B1(new_n1160), .B2(new_n1182), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT57), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n1207), .B2(new_n1211), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1164), .B1(new_n1241), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT122), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1207), .A2(new_n1211), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1167), .A2(new_n1181), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(KEYINPUT121), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1167), .A2(new_n1238), .A3(new_n1181), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1246), .B1(new_n1250), .B2(new_n1186), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n1244), .A2(new_n1245), .B1(new_n1251), .B2(KEYINPUT57), .ZN(new_n1252));
  AOI211_X1 g1052(.A(KEYINPUT122), .B(new_n1164), .C1(new_n1241), .C2(new_n1243), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1237), .B1(new_n1252), .B2(new_n1253), .ZN(G375));
  NAND2_X1  g1054(.A1(new_n808), .A2(G303), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n289), .B1(new_n799), .B2(G97), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n978), .A2(new_n1255), .A3(new_n1055), .A4(new_n1256), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n828), .A2(new_n879), .B1(new_n424), .B2(new_n802), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n1257), .B(new_n1258), .C1(G294), .C2(new_n819), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n796), .A2(G116), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n795), .A2(new_n1139), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n808), .A2(G128), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n811), .A2(G50), .B1(new_n799), .B2(G159), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1262), .B(new_n1263), .C1(new_n1138), .C2(new_n818), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n828), .A2(new_n1134), .B1(new_n864), .B2(new_n802), .ZN(new_n1265));
  NOR3_X1   g1065(.A1(new_n1261), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1217), .A2(new_n546), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(KEYINPUT123), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1259), .A2(new_n1260), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1269));
  OAI221_X1 g1069(.A(new_n769), .B1(G68), .B2(new_n1214), .C1(new_n1269), .C2(new_n861), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1270), .B1(new_n1123), .B2(new_n782), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(new_n1179), .B2(new_n768), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT124), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1272), .B(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1179), .B1(new_n1167), .B2(new_n1181), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1182), .A2(new_n1038), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1274), .B1(new_n1275), .B2(new_n1276), .ZN(G381));
  OR2_X1    g1077(.A1(G393), .A2(G396), .ZN(new_n1278));
  OR3_X1    g1078(.A1(G381), .A2(G384), .A3(new_n1278), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1150), .B1(new_n1160), .B2(new_n767), .ZN(new_n1281));
  OR2_X1    g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(G390), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1041), .A2(new_n1283), .ZN(new_n1284));
  OR4_X1    g1084(.A1(G375), .A2(new_n1279), .A3(new_n1282), .A4(new_n1284), .ZN(G407));
  INV_X1    g1085(.A(new_n1237), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT57), .B1(new_n1241), .B2(new_n1212), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1248), .A2(new_n1249), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1243), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n722), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1287), .B1(new_n1290), .B2(KEYINPUT122), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1253), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1286), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1282), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n697), .A2(G343), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1293), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(G407), .A2(G213), .A3(new_n1296), .ZN(G409));
  NAND2_X1  g1097(.A1(new_n1251), .A2(new_n1038), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1237), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1294), .A2(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1300), .B1(G375), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1295), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1179), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1247), .A2(KEYINPUT60), .A3(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n722), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1275), .B1(KEYINPUT60), .B2(new_n1182), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1274), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(G384), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  OAI211_X1 g1110(.A(new_n1274), .B(G384), .C1(new_n1307), .C2(new_n1306), .ZN(new_n1311));
  AND3_X1   g1111(.A1(new_n1310), .A2(new_n1311), .A3(KEYINPUT125), .ZN(new_n1312));
  AOI21_X1  g1112(.A(KEYINPUT125), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1302), .A2(new_n1303), .A3(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(KEYINPUT62), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT125), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1310), .A2(new_n1311), .A3(KEYINPUT125), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1295), .A2(G2897), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1319), .A2(new_n1320), .A3(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1317), .A2(G2897), .A3(new_n1295), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1282), .B1(new_n1237), .B2(new_n1298), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1324), .B1(new_n1293), .B2(G378), .ZN(new_n1325));
  OAI211_X1 g1125(.A(new_n1322), .B(new_n1323), .C1(new_n1325), .C2(new_n1295), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT61), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT62), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1302), .A2(new_n1314), .A3(new_n1328), .A4(new_n1303), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1316), .A2(new_n1326), .A3(new_n1327), .A4(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT126), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(G393), .A2(G396), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1278), .A2(new_n1332), .ZN(new_n1333));
  NOR3_X1   g1133(.A1(new_n1020), .A2(new_n1039), .A3(new_n1021), .ZN(new_n1334));
  OAI21_X1  g1134(.A(G390), .B1(new_n1334), .B2(new_n993), .ZN(new_n1335));
  AOI211_X1 g1135(.A(new_n1331), .B(new_n1333), .C1(new_n1284), .C2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1333), .A2(new_n1331), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1333), .A2(new_n1331), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  AND4_X1   g1139(.A1(new_n1284), .A2(new_n1335), .A3(new_n1337), .A4(new_n1339), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1336), .A2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1330), .A2(new_n1342), .ZN(new_n1343));
  AND2_X1   g1143(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1345));
  AOI21_X1  g1145(.A(KEYINPUT61), .B1(new_n1344), .B2(new_n1345), .ZN(new_n1346));
  NAND4_X1  g1146(.A1(new_n1302), .A2(new_n1314), .A3(KEYINPUT63), .A4(new_n1303), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT63), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1315), .A2(new_n1348), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1346), .A2(new_n1347), .A3(new_n1341), .A4(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1343), .A2(new_n1350), .ZN(G405));
  INV_X1    g1151(.A(KEYINPUT127), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1352), .B1(new_n1336), .B2(new_n1340), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1284), .A2(new_n1335), .A3(new_n1337), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1354), .A2(new_n1338), .ZN(new_n1355));
  NAND4_X1  g1155(.A1(new_n1284), .A2(new_n1335), .A3(new_n1337), .A4(new_n1339), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1355), .A2(KEYINPUT127), .A3(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1353), .A2(new_n1357), .ZN(new_n1358));
  NOR2_X1   g1158(.A1(new_n1293), .A2(new_n1282), .ZN(new_n1359));
  NOR2_X1   g1159(.A1(G375), .A2(new_n1301), .ZN(new_n1360));
  NOR2_X1   g1160(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1361), .A2(new_n1317), .ZN(new_n1362));
  OAI21_X1  g1162(.A(new_n1314), .B1(new_n1359), .B2(new_n1360), .ZN(new_n1363));
  AND3_X1   g1163(.A1(new_n1358), .A2(new_n1362), .A3(new_n1363), .ZN(new_n1364));
  AOI21_X1  g1164(.A(new_n1358), .B1(new_n1362), .B2(new_n1363), .ZN(new_n1365));
  NOR2_X1   g1165(.A1(new_n1364), .A2(new_n1365), .ZN(G402));
endmodule


