

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U551 ( .A(n720), .ZN(n734) );
  NOR2_X1 U552 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X2 U553 ( .A(KEYINPUT17), .B(n522), .Z(n988) );
  NOR2_X1 U554 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U555 ( .A1(n734), .A2(n867), .ZN(n697) );
  AND2_X1 U556 ( .A1(n693), .A2(n788), .ZN(n720) );
  INV_X1 U557 ( .A(KEYINPUT26), .ZN(n515) );
  XNOR2_X1 U558 ( .A(n697), .B(n515), .ZN(n699) );
  NOR2_X2 U559 ( .A1(G2105), .A2(n523), .ZN(n990) );
  XNOR2_X1 U560 ( .A(n516), .B(KEYINPUT23), .ZN(n517) );
  INV_X1 U561 ( .A(KEYINPUT64), .ZN(n516) );
  INV_X1 U562 ( .A(G2104), .ZN(n523) );
  NOR2_X1 U563 ( .A1(G651), .A2(n535), .ZN(n651) );
  XNOR2_X1 U564 ( .A(n518), .B(n517), .ZN(n521) );
  NOR2_X1 U565 ( .A1(n527), .A2(n526), .ZN(G160) );
  NAND2_X1 U566 ( .A1(G101), .A2(n990), .ZN(n518) );
  NAND2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n519) );
  XNOR2_X1 U568 ( .A(n519), .B(KEYINPUT65), .ZN(n996) );
  NAND2_X1 U569 ( .A1(G113), .A2(n996), .ZN(n520) );
  NAND2_X1 U570 ( .A1(n521), .A2(n520), .ZN(n527) );
  NOR2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  NAND2_X1 U572 ( .A1(G137), .A2(n988), .ZN(n525) );
  AND2_X1 U573 ( .A1(n523), .A2(G2105), .ZN(n997) );
  NAND2_X1 U574 ( .A1(G125), .A2(n997), .ZN(n524) );
  NAND2_X1 U575 ( .A1(n525), .A2(n524), .ZN(n526) );
  INV_X1 U576 ( .A(G651), .ZN(n536) );
  NOR2_X1 U577 ( .A1(G543), .A2(n536), .ZN(n528) );
  XOR2_X1 U578 ( .A(KEYINPUT68), .B(n528), .Z(n529) );
  XNOR2_X1 U579 ( .A(KEYINPUT1), .B(n529), .ZN(n658) );
  NAND2_X1 U580 ( .A1(G63), .A2(n658), .ZN(n530) );
  XOR2_X1 U581 ( .A(KEYINPUT79), .B(n530), .Z(n532) );
  XOR2_X1 U582 ( .A(G543), .B(KEYINPUT0), .Z(n535) );
  NAND2_X1 U583 ( .A1(n651), .A2(G51), .ZN(n531) );
  NAND2_X1 U584 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U585 ( .A(KEYINPUT6), .B(n533), .ZN(n543) );
  NOR2_X1 U586 ( .A1(G543), .A2(G651), .ZN(n639) );
  NAND2_X1 U587 ( .A1(n639), .A2(G89), .ZN(n534) );
  XNOR2_X1 U588 ( .A(n534), .B(KEYINPUT4), .ZN(n539) );
  OR2_X1 U589 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X2 U590 ( .A(n537), .B(KEYINPUT67), .ZN(n642) );
  NAND2_X1 U591 ( .A1(G76), .A2(n642), .ZN(n538) );
  NAND2_X1 U592 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U593 ( .A(KEYINPUT78), .B(n540), .Z(n541) );
  XNOR2_X1 U594 ( .A(KEYINPUT5), .B(n541), .ZN(n542) );
  NOR2_X1 U595 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U596 ( .A(KEYINPUT7), .B(n544), .Z(G168) );
  XOR2_X1 U597 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U598 ( .A(G2427), .B(G2446), .Z(n546) );
  XNOR2_X1 U599 ( .A(G1348), .B(G2430), .ZN(n545) );
  XNOR2_X1 U600 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U601 ( .A(n547), .B(G2435), .Z(n549) );
  XNOR2_X1 U602 ( .A(G1341), .B(G2438), .ZN(n548) );
  XNOR2_X1 U603 ( .A(n549), .B(n548), .ZN(n553) );
  XOR2_X1 U604 ( .A(G2454), .B(G2451), .Z(n551) );
  XNOR2_X1 U605 ( .A(KEYINPUT104), .B(G2443), .ZN(n550) );
  XNOR2_X1 U606 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U607 ( .A(n553), .B(n552), .Z(n554) );
  AND2_X1 U608 ( .A1(G14), .A2(n554), .ZN(G401) );
  NAND2_X1 U609 ( .A1(G52), .A2(n651), .ZN(n556) );
  NAND2_X1 U610 ( .A1(G64), .A2(n658), .ZN(n555) );
  NAND2_X1 U611 ( .A1(n556), .A2(n555), .ZN(n561) );
  NAND2_X1 U612 ( .A1(G90), .A2(n639), .ZN(n558) );
  NAND2_X1 U613 ( .A1(G77), .A2(n642), .ZN(n557) );
  NAND2_X1 U614 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U615 ( .A(KEYINPUT9), .B(n559), .Z(n560) );
  NOR2_X1 U616 ( .A1(n561), .A2(n560), .ZN(G171) );
  AND2_X1 U617 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U618 ( .A1(G111), .A2(n996), .ZN(n562) );
  XNOR2_X1 U619 ( .A(n562), .B(KEYINPUT82), .ZN(n569) );
  NAND2_X1 U620 ( .A1(G99), .A2(n990), .ZN(n564) );
  NAND2_X1 U621 ( .A1(G135), .A2(n988), .ZN(n563) );
  NAND2_X1 U622 ( .A1(n564), .A2(n563), .ZN(n567) );
  NAND2_X1 U623 ( .A1(n997), .A2(G123), .ZN(n565) );
  XOR2_X1 U624 ( .A(KEYINPUT18), .B(n565), .Z(n566) );
  NOR2_X1 U625 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U626 ( .A1(n569), .A2(n568), .ZN(n976) );
  XNOR2_X1 U627 ( .A(G2096), .B(n976), .ZN(n570) );
  OR2_X1 U628 ( .A1(G2100), .A2(n570), .ZN(G156) );
  INV_X1 U629 ( .A(G132), .ZN(G219) );
  NAND2_X1 U630 ( .A1(G91), .A2(n639), .ZN(n572) );
  NAND2_X1 U631 ( .A1(G78), .A2(n642), .ZN(n571) );
  NAND2_X1 U632 ( .A1(n572), .A2(n571), .ZN(n577) );
  NAND2_X1 U633 ( .A1(G53), .A2(n651), .ZN(n574) );
  NAND2_X1 U634 ( .A1(G65), .A2(n658), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U636 ( .A(KEYINPUT70), .B(n575), .ZN(n576) );
  NOR2_X1 U637 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U638 ( .A(n578), .B(KEYINPUT71), .ZN(G299) );
  NAND2_X1 U639 ( .A1(G7), .A2(G661), .ZN(n579) );
  XNOR2_X1 U640 ( .A(n579), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U641 ( .A(KEYINPUT11), .B(KEYINPUT74), .Z(n581) );
  INV_X1 U642 ( .A(G223), .ZN(n822) );
  NAND2_X1 U643 ( .A1(G567), .A2(n822), .ZN(n580) );
  XNOR2_X1 U644 ( .A(n581), .B(n580), .ZN(G234) );
  NAND2_X1 U645 ( .A1(n639), .A2(G81), .ZN(n582) );
  XNOR2_X1 U646 ( .A(KEYINPUT12), .B(n582), .ZN(n586) );
  NAND2_X1 U647 ( .A1(n642), .A2(G68), .ZN(n584) );
  INV_X1 U648 ( .A(KEYINPUT75), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n585) );
  NAND2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(n587), .B(KEYINPUT13), .ZN(n589) );
  NAND2_X1 U652 ( .A1(G43), .A2(n651), .ZN(n588) );
  NAND2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U654 ( .A1(n658), .A2(G56), .ZN(n590) );
  XOR2_X1 U655 ( .A(KEYINPUT14), .B(n590), .Z(n591) );
  XOR2_X2 U656 ( .A(n593), .B(KEYINPUT76), .Z(n952) );
  INV_X1 U657 ( .A(n952), .ZN(n594) );
  NAND2_X1 U658 ( .A1(G860), .A2(n594), .ZN(G153) );
  INV_X1 U659 ( .A(G171), .ZN(G301) );
  NAND2_X1 U660 ( .A1(G868), .A2(G301), .ZN(n604) );
  NAND2_X1 U661 ( .A1(G79), .A2(n642), .ZN(n596) );
  NAND2_X1 U662 ( .A1(G54), .A2(n651), .ZN(n595) );
  NAND2_X1 U663 ( .A1(n596), .A2(n595), .ZN(n601) );
  NAND2_X1 U664 ( .A1(G92), .A2(n639), .ZN(n598) );
  NAND2_X1 U665 ( .A1(G66), .A2(n658), .ZN(n597) );
  NAND2_X1 U666 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U667 ( .A(KEYINPUT77), .B(n599), .Z(n600) );
  NOR2_X1 U668 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U669 ( .A(KEYINPUT15), .B(n602), .ZN(n706) );
  INV_X1 U670 ( .A(G868), .ZN(n671) );
  NAND2_X1 U671 ( .A1(n706), .A2(n671), .ZN(n603) );
  NAND2_X1 U672 ( .A1(n604), .A2(n603), .ZN(G284) );
  XNOR2_X1 U673 ( .A(KEYINPUT80), .B(n671), .ZN(n605) );
  NOR2_X1 U674 ( .A1(G286), .A2(n605), .ZN(n607) );
  NOR2_X1 U675 ( .A1(G868), .A2(G299), .ZN(n606) );
  NOR2_X1 U676 ( .A1(n607), .A2(n606), .ZN(G297) );
  INV_X1 U677 ( .A(G559), .ZN(n608) );
  NOR2_X1 U678 ( .A1(G860), .A2(n608), .ZN(n609) );
  XNOR2_X1 U679 ( .A(KEYINPUT81), .B(n609), .ZN(n610) );
  INV_X1 U680 ( .A(n706), .ZN(n948) );
  NAND2_X1 U681 ( .A1(n610), .A2(n948), .ZN(n611) );
  XNOR2_X1 U682 ( .A(n611), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U683 ( .A1(n952), .A2(G868), .ZN(n614) );
  NAND2_X1 U684 ( .A1(G868), .A2(n948), .ZN(n612) );
  NOR2_X1 U685 ( .A1(G559), .A2(n612), .ZN(n613) );
  NOR2_X1 U686 ( .A1(n614), .A2(n613), .ZN(G282) );
  NAND2_X1 U687 ( .A1(G93), .A2(n639), .ZN(n616) );
  NAND2_X1 U688 ( .A1(G80), .A2(n642), .ZN(n615) );
  NAND2_X1 U689 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U690 ( .A(KEYINPUT83), .B(n617), .ZN(n622) );
  NAND2_X1 U691 ( .A1(G55), .A2(n651), .ZN(n619) );
  NAND2_X1 U692 ( .A1(G67), .A2(n658), .ZN(n618) );
  NAND2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U694 ( .A(KEYINPUT84), .B(n620), .Z(n621) );
  NAND2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n670) );
  NAND2_X1 U696 ( .A1(G559), .A2(n948), .ZN(n623) );
  XNOR2_X1 U697 ( .A(n623), .B(n952), .ZN(n668) );
  NOR2_X1 U698 ( .A1(n668), .A2(G860), .ZN(n624) );
  XOR2_X1 U699 ( .A(n670), .B(n624), .Z(G145) );
  NAND2_X1 U700 ( .A1(G88), .A2(n639), .ZN(n626) );
  NAND2_X1 U701 ( .A1(G75), .A2(n642), .ZN(n625) );
  NAND2_X1 U702 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U703 ( .A1(G50), .A2(n651), .ZN(n628) );
  NAND2_X1 U704 ( .A1(G62), .A2(n658), .ZN(n627) );
  NAND2_X1 U705 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U706 ( .A1(n630), .A2(n629), .ZN(G166) );
  NAND2_X1 U707 ( .A1(G60), .A2(n658), .ZN(n637) );
  NAND2_X1 U708 ( .A1(n651), .A2(G47), .ZN(n632) );
  NAND2_X1 U709 ( .A1(n642), .A2(G72), .ZN(n631) );
  NAND2_X1 U710 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U711 ( .A1(G85), .A2(n639), .ZN(n633) );
  XOR2_X1 U712 ( .A(KEYINPUT66), .B(n633), .Z(n634) );
  NOR2_X1 U713 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U714 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U715 ( .A(KEYINPUT69), .B(n638), .Z(G290) );
  NAND2_X1 U716 ( .A1(G86), .A2(n639), .ZN(n641) );
  NAND2_X1 U717 ( .A1(G61), .A2(n658), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n641), .A2(n640), .ZN(n647) );
  XOR2_X1 U719 ( .A(KEYINPUT89), .B(KEYINPUT2), .Z(n644) );
  NAND2_X1 U720 ( .A1(G73), .A2(n642), .ZN(n643) );
  XNOR2_X1 U721 ( .A(n644), .B(n643), .ZN(n645) );
  XOR2_X1 U722 ( .A(KEYINPUT88), .B(n645), .Z(n646) );
  NOR2_X1 U723 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U724 ( .A(n648), .B(KEYINPUT90), .ZN(n650) );
  NAND2_X1 U725 ( .A1(G48), .A2(n651), .ZN(n649) );
  NAND2_X1 U726 ( .A1(n650), .A2(n649), .ZN(G305) );
  NAND2_X1 U727 ( .A1(n651), .A2(G49), .ZN(n652) );
  XOR2_X1 U728 ( .A(KEYINPUT85), .B(n652), .Z(n654) );
  NAND2_X1 U729 ( .A1(G651), .A2(G74), .ZN(n653) );
  NAND2_X1 U730 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U731 ( .A(KEYINPUT86), .B(n655), .Z(n660) );
  NAND2_X1 U732 ( .A1(G87), .A2(n535), .ZN(n656) );
  XNOR2_X1 U733 ( .A(KEYINPUT87), .B(n656), .ZN(n657) );
  NOR2_X1 U734 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U735 ( .A1(n660), .A2(n659), .ZN(G288) );
  XOR2_X1 U736 ( .A(KEYINPUT19), .B(KEYINPUT92), .Z(n662) );
  XNOR2_X1 U737 ( .A(G166), .B(KEYINPUT91), .ZN(n661) );
  XNOR2_X1 U738 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U739 ( .A(n663), .B(G290), .ZN(n666) );
  XNOR2_X1 U740 ( .A(G305), .B(G288), .ZN(n664) );
  XNOR2_X1 U741 ( .A(n664), .B(n670), .ZN(n665) );
  XNOR2_X1 U742 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U743 ( .A(n667), .B(G299), .ZN(n951) );
  XNOR2_X1 U744 ( .A(n668), .B(n951), .ZN(n669) );
  NAND2_X1 U745 ( .A1(n669), .A2(G868), .ZN(n673) );
  NAND2_X1 U746 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U747 ( .A1(n673), .A2(n672), .ZN(G295) );
  NAND2_X1 U748 ( .A1(G2078), .A2(G2084), .ZN(n674) );
  XOR2_X1 U749 ( .A(KEYINPUT20), .B(n674), .Z(n675) );
  NAND2_X1 U750 ( .A1(G2090), .A2(n675), .ZN(n676) );
  XNOR2_X1 U751 ( .A(KEYINPUT21), .B(n676), .ZN(n677) );
  NAND2_X1 U752 ( .A1(n677), .A2(G2072), .ZN(G158) );
  XOR2_X1 U753 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  XNOR2_X1 U754 ( .A(KEYINPUT73), .B(G82), .ZN(G220) );
  XNOR2_X1 U755 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U756 ( .A1(G108), .A2(G120), .ZN(n678) );
  NOR2_X1 U757 ( .A1(G237), .A2(n678), .ZN(n679) );
  NAND2_X1 U758 ( .A1(G69), .A2(n679), .ZN(n946) );
  NAND2_X1 U759 ( .A1(n946), .A2(G567), .ZN(n685) );
  NOR2_X1 U760 ( .A1(G219), .A2(G220), .ZN(n681) );
  XNOR2_X1 U761 ( .A(KEYINPUT22), .B(KEYINPUT93), .ZN(n680) );
  XNOR2_X1 U762 ( .A(n681), .B(n680), .ZN(n682) );
  NOR2_X1 U763 ( .A1(n682), .A2(G218), .ZN(n683) );
  NAND2_X1 U764 ( .A1(G96), .A2(n683), .ZN(n947) );
  NAND2_X1 U765 ( .A1(n947), .A2(G2106), .ZN(n684) );
  NAND2_X1 U766 ( .A1(n685), .A2(n684), .ZN(n1014) );
  NAND2_X1 U767 ( .A1(G661), .A2(G483), .ZN(n686) );
  NOR2_X1 U768 ( .A1(n1014), .A2(n686), .ZN(n825) );
  NAND2_X1 U769 ( .A1(n825), .A2(G36), .ZN(G176) );
  NAND2_X1 U770 ( .A1(G102), .A2(n990), .ZN(n688) );
  NAND2_X1 U771 ( .A1(G138), .A2(n988), .ZN(n687) );
  NAND2_X1 U772 ( .A1(n688), .A2(n687), .ZN(n692) );
  NAND2_X1 U773 ( .A1(G114), .A2(n996), .ZN(n690) );
  NAND2_X1 U774 ( .A1(G126), .A2(n997), .ZN(n689) );
  NAND2_X1 U775 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U776 ( .A1(n692), .A2(n691), .ZN(G164) );
  INV_X1 U777 ( .A(G166), .ZN(G303) );
  XOR2_X1 U778 ( .A(G1981), .B(G305), .Z(n889) );
  NAND2_X1 U779 ( .A1(G160), .A2(G40), .ZN(n789) );
  INV_X1 U780 ( .A(n789), .ZN(n693) );
  NOR2_X1 U781 ( .A1(G164), .A2(G1384), .ZN(n788) );
  NAND2_X1 U782 ( .A1(G8), .A2(n734), .ZN(n766) );
  INV_X1 U783 ( .A(n766), .ZN(n760) );
  NOR2_X1 U784 ( .A1(G288), .A2(G1976), .ZN(n694) );
  XOR2_X1 U785 ( .A(n694), .B(KEYINPUT99), .Z(n903) );
  AND2_X1 U786 ( .A1(n760), .A2(n903), .ZN(n695) );
  NAND2_X1 U787 ( .A1(KEYINPUT33), .A2(n695), .ZN(n696) );
  NAND2_X1 U788 ( .A1(n889), .A2(n696), .ZN(n758) );
  INV_X1 U789 ( .A(G1996), .ZN(n867) );
  NAND2_X1 U790 ( .A1(n734), .A2(G1341), .ZN(n698) );
  NAND2_X1 U791 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U792 ( .A1(n952), .A2(n700), .ZN(n704) );
  NAND2_X1 U793 ( .A1(G1348), .A2(n734), .ZN(n702) );
  NAND2_X1 U794 ( .A1(G2067), .A2(n720), .ZN(n701) );
  NAND2_X1 U795 ( .A1(n702), .A2(n701), .ZN(n705) );
  NOR2_X1 U796 ( .A1(n706), .A2(n705), .ZN(n703) );
  NOR2_X1 U797 ( .A1(n704), .A2(n703), .ZN(n708) );
  AND2_X1 U798 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U799 ( .A1(n708), .A2(n707), .ZN(n714) );
  NAND2_X1 U800 ( .A1(n720), .A2(G2072), .ZN(n709) );
  XOR2_X1 U801 ( .A(KEYINPUT27), .B(n709), .Z(n711) );
  NAND2_X1 U802 ( .A1(G1956), .A2(n734), .ZN(n710) );
  NAND2_X1 U803 ( .A1(n711), .A2(n710), .ZN(n715) );
  NOR2_X1 U804 ( .A1(G299), .A2(n715), .ZN(n712) );
  XNOR2_X1 U805 ( .A(n712), .B(KEYINPUT98), .ZN(n713) );
  NOR2_X1 U806 ( .A1(n714), .A2(n713), .ZN(n718) );
  NAND2_X1 U807 ( .A1(G299), .A2(n715), .ZN(n716) );
  XOR2_X1 U808 ( .A(KEYINPUT28), .B(n716), .Z(n717) );
  XNOR2_X1 U809 ( .A(n719), .B(KEYINPUT29), .ZN(n724) );
  INV_X1 U810 ( .A(G1961), .ZN(n911) );
  NAND2_X1 U811 ( .A1(n734), .A2(n911), .ZN(n722) );
  XNOR2_X1 U812 ( .A(G2078), .B(KEYINPUT25), .ZN(n865) );
  NAND2_X1 U813 ( .A1(n720), .A2(n865), .ZN(n721) );
  NAND2_X1 U814 ( .A1(n722), .A2(n721), .ZN(n728) );
  NAND2_X1 U815 ( .A1(G171), .A2(n728), .ZN(n723) );
  NAND2_X1 U816 ( .A1(n724), .A2(n723), .ZN(n733) );
  NOR2_X1 U817 ( .A1(G1966), .A2(n766), .ZN(n746) );
  NOR2_X1 U818 ( .A1(G2084), .A2(n734), .ZN(n742) );
  NOR2_X1 U819 ( .A1(n746), .A2(n742), .ZN(n725) );
  NAND2_X1 U820 ( .A1(G8), .A2(n725), .ZN(n726) );
  XNOR2_X1 U821 ( .A(KEYINPUT30), .B(n726), .ZN(n727) );
  NOR2_X1 U822 ( .A1(G168), .A2(n727), .ZN(n730) );
  NOR2_X1 U823 ( .A1(G171), .A2(n728), .ZN(n729) );
  NOR2_X1 U824 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U825 ( .A(KEYINPUT31), .B(n731), .Z(n732) );
  NAND2_X1 U826 ( .A1(n733), .A2(n732), .ZN(n744) );
  NAND2_X1 U827 ( .A1(n744), .A2(G286), .ZN(n739) );
  NOR2_X1 U828 ( .A1(G1971), .A2(n766), .ZN(n736) );
  NOR2_X1 U829 ( .A1(G2090), .A2(n734), .ZN(n735) );
  NOR2_X1 U830 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U831 ( .A1(n737), .A2(G303), .ZN(n738) );
  NAND2_X1 U832 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U833 ( .A1(n740), .A2(G8), .ZN(n741) );
  XNOR2_X1 U834 ( .A(n741), .B(KEYINPUT32), .ZN(n750) );
  NAND2_X1 U835 ( .A1(G8), .A2(n742), .ZN(n743) );
  XOR2_X1 U836 ( .A(KEYINPUT97), .B(n743), .Z(n748) );
  INV_X1 U837 ( .A(n744), .ZN(n745) );
  NOR2_X1 U838 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U839 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U840 ( .A1(n750), .A2(n749), .ZN(n762) );
  NOR2_X1 U841 ( .A1(G1971), .A2(G303), .ZN(n751) );
  NOR2_X1 U842 ( .A1(n903), .A2(n751), .ZN(n752) );
  NAND2_X1 U843 ( .A1(n762), .A2(n752), .ZN(n753) );
  NAND2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n896) );
  NAND2_X1 U845 ( .A1(n753), .A2(n896), .ZN(n754) );
  XNOR2_X1 U846 ( .A(n754), .B(KEYINPUT100), .ZN(n755) );
  NOR2_X1 U847 ( .A1(n766), .A2(n755), .ZN(n756) );
  NOR2_X1 U848 ( .A1(KEYINPUT33), .A2(n756), .ZN(n757) );
  NOR2_X1 U849 ( .A1(n758), .A2(n757), .ZN(n770) );
  NOR2_X1 U850 ( .A1(G1981), .A2(G305), .ZN(n759) );
  XNOR2_X1 U851 ( .A(KEYINPUT24), .B(n759), .ZN(n761) );
  NAND2_X1 U852 ( .A1(n761), .A2(n760), .ZN(n768) );
  NOR2_X1 U853 ( .A1(G2090), .A2(G303), .ZN(n763) );
  NAND2_X1 U854 ( .A1(G8), .A2(n763), .ZN(n764) );
  NAND2_X1 U855 ( .A1(n762), .A2(n764), .ZN(n765) );
  NAND2_X1 U856 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U857 ( .A1(n768), .A2(n767), .ZN(n769) );
  NOR2_X1 U858 ( .A1(n770), .A2(n769), .ZN(n803) );
  XOR2_X1 U859 ( .A(G1986), .B(G290), .Z(n892) );
  NAND2_X1 U860 ( .A1(G95), .A2(n990), .ZN(n771) );
  XNOR2_X1 U861 ( .A(n771), .B(KEYINPUT96), .ZN(n774) );
  NAND2_X1 U862 ( .A1(G119), .A2(n997), .ZN(n772) );
  XOR2_X1 U863 ( .A(KEYINPUT95), .B(n772), .Z(n773) );
  NAND2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n778) );
  NAND2_X1 U865 ( .A1(G107), .A2(n996), .ZN(n776) );
  NAND2_X1 U866 ( .A1(G131), .A2(n988), .ZN(n775) );
  NAND2_X1 U867 ( .A1(n776), .A2(n775), .ZN(n777) );
  OR2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n980) );
  AND2_X1 U869 ( .A1(n980), .A2(G1991), .ZN(n787) );
  NAND2_X1 U870 ( .A1(n990), .A2(G105), .ZN(n779) );
  XNOR2_X1 U871 ( .A(n779), .B(KEYINPUT38), .ZN(n781) );
  NAND2_X1 U872 ( .A1(G117), .A2(n996), .ZN(n780) );
  NAND2_X1 U873 ( .A1(n781), .A2(n780), .ZN(n785) );
  NAND2_X1 U874 ( .A1(G141), .A2(n988), .ZN(n783) );
  NAND2_X1 U875 ( .A1(G129), .A2(n997), .ZN(n782) );
  NAND2_X1 U876 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U877 ( .A1(n785), .A2(n784), .ZN(n979) );
  NOR2_X1 U878 ( .A1(n867), .A2(n979), .ZN(n786) );
  NOR2_X1 U879 ( .A1(n787), .A2(n786), .ZN(n851) );
  NAND2_X1 U880 ( .A1(n892), .A2(n851), .ZN(n790) );
  NOR2_X1 U881 ( .A1(n789), .A2(n788), .ZN(n817) );
  NAND2_X1 U882 ( .A1(n790), .A2(n817), .ZN(n801) );
  NAND2_X1 U883 ( .A1(G104), .A2(n990), .ZN(n792) );
  NAND2_X1 U884 ( .A1(G140), .A2(n988), .ZN(n791) );
  NAND2_X1 U885 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U886 ( .A(KEYINPUT34), .B(n793), .ZN(n798) );
  NAND2_X1 U887 ( .A1(G116), .A2(n996), .ZN(n795) );
  NAND2_X1 U888 ( .A1(G128), .A2(n997), .ZN(n794) );
  NAND2_X1 U889 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U890 ( .A(KEYINPUT35), .B(n796), .Z(n797) );
  NOR2_X1 U891 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U892 ( .A(KEYINPUT36), .B(n799), .Z(n1004) );
  XOR2_X1 U893 ( .A(G2067), .B(KEYINPUT37), .Z(n805) );
  AND2_X1 U894 ( .A1(n1004), .A2(n805), .ZN(n853) );
  NAND2_X1 U895 ( .A1(n853), .A2(n817), .ZN(n800) );
  XNOR2_X1 U896 ( .A(n800), .B(KEYINPUT94), .ZN(n806) );
  NAND2_X1 U897 ( .A1(n801), .A2(n806), .ZN(n802) );
  NOR2_X2 U898 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U899 ( .A(n804), .B(KEYINPUT101), .ZN(n820) );
  NOR2_X1 U900 ( .A1(n1004), .A2(n805), .ZN(n857) );
  INV_X1 U901 ( .A(n806), .ZN(n813) );
  AND2_X1 U902 ( .A1(n867), .A2(n979), .ZN(n844) );
  INV_X1 U903 ( .A(n851), .ZN(n809) );
  NOR2_X1 U904 ( .A1(G1986), .A2(G290), .ZN(n807) );
  NOR2_X1 U905 ( .A1(G1991), .A2(n980), .ZN(n848) );
  NOR2_X1 U906 ( .A1(n807), .A2(n848), .ZN(n808) );
  NOR2_X1 U907 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U908 ( .A1(n844), .A2(n810), .ZN(n811) );
  XOR2_X1 U909 ( .A(KEYINPUT39), .B(n811), .Z(n812) );
  NOR2_X1 U910 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U911 ( .A(n814), .B(KEYINPUT102), .ZN(n815) );
  NOR2_X1 U912 ( .A1(n857), .A2(n815), .ZN(n816) );
  XNOR2_X1 U913 ( .A(KEYINPUT103), .B(n816), .ZN(n818) );
  NAND2_X1 U914 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U915 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U916 ( .A(n821), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n822), .ZN(G217) );
  AND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n823) );
  NAND2_X1 U919 ( .A1(G661), .A2(n823), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U921 ( .A1(n825), .A2(n824), .ZN(G188) );
  XNOR2_X1 U922 ( .A(G96), .B(KEYINPUT105), .ZN(G221) );
  NAND2_X1 U924 ( .A1(G124), .A2(n997), .ZN(n826) );
  XNOR2_X1 U925 ( .A(n826), .B(KEYINPUT44), .ZN(n828) );
  NAND2_X1 U926 ( .A1(n996), .A2(G112), .ZN(n827) );
  NAND2_X1 U927 ( .A1(n828), .A2(n827), .ZN(n832) );
  NAND2_X1 U928 ( .A1(G100), .A2(n990), .ZN(n830) );
  NAND2_X1 U929 ( .A1(G136), .A2(n988), .ZN(n829) );
  NAND2_X1 U930 ( .A1(n830), .A2(n829), .ZN(n831) );
  NOR2_X1 U931 ( .A1(n832), .A2(n831), .ZN(G162) );
  NAND2_X1 U932 ( .A1(G103), .A2(n990), .ZN(n834) );
  NAND2_X1 U933 ( .A1(G139), .A2(n988), .ZN(n833) );
  NAND2_X1 U934 ( .A1(n834), .A2(n833), .ZN(n839) );
  NAND2_X1 U935 ( .A1(G115), .A2(n996), .ZN(n836) );
  NAND2_X1 U936 ( .A1(G127), .A2(n997), .ZN(n835) );
  NAND2_X1 U937 ( .A1(n836), .A2(n835), .ZN(n837) );
  XOR2_X1 U938 ( .A(KEYINPUT47), .B(n837), .Z(n838) );
  NOR2_X1 U939 ( .A1(n839), .A2(n838), .ZN(n985) );
  XOR2_X1 U940 ( .A(G2072), .B(n985), .Z(n841) );
  XOR2_X1 U941 ( .A(G164), .B(G2078), .Z(n840) );
  NOR2_X1 U942 ( .A1(n841), .A2(n840), .ZN(n842) );
  XOR2_X1 U943 ( .A(KEYINPUT50), .B(n842), .Z(n860) );
  XOR2_X1 U944 ( .A(G2090), .B(G162), .Z(n843) );
  NOR2_X1 U945 ( .A1(n844), .A2(n843), .ZN(n845) );
  XOR2_X1 U946 ( .A(KEYINPUT51), .B(n845), .Z(n855) );
  XNOR2_X1 U947 ( .A(G160), .B(G2084), .ZN(n846) );
  NAND2_X1 U948 ( .A1(n846), .A2(n976), .ZN(n847) );
  NOR2_X1 U949 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n849), .B(KEYINPUT116), .ZN(n850) );
  NAND2_X1 U951 ( .A1(n851), .A2(n850), .ZN(n852) );
  NOR2_X1 U952 ( .A1(n853), .A2(n852), .ZN(n854) );
  NAND2_X1 U953 ( .A1(n855), .A2(n854), .ZN(n856) );
  NOR2_X1 U954 ( .A1(n857), .A2(n856), .ZN(n858) );
  XNOR2_X1 U955 ( .A(KEYINPUT117), .B(n858), .ZN(n859) );
  NOR2_X1 U956 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U957 ( .A(KEYINPUT52), .B(n861), .ZN(n862) );
  INV_X1 U958 ( .A(KEYINPUT55), .ZN(n885) );
  NAND2_X1 U959 ( .A1(n862), .A2(n885), .ZN(n863) );
  NAND2_X1 U960 ( .A1(n863), .A2(G29), .ZN(n944) );
  XNOR2_X1 U961 ( .A(G2084), .B(G34), .ZN(n864) );
  XNOR2_X1 U962 ( .A(n864), .B(KEYINPUT54), .ZN(n880) );
  XNOR2_X1 U963 ( .A(G27), .B(n865), .ZN(n872) );
  XOR2_X1 U964 ( .A(G25), .B(G1991), .Z(n866) );
  NAND2_X1 U965 ( .A1(n866), .A2(G28), .ZN(n870) );
  XOR2_X1 U966 ( .A(G32), .B(n867), .Z(n868) );
  XNOR2_X1 U967 ( .A(KEYINPUT120), .B(n868), .ZN(n869) );
  NOR2_X1 U968 ( .A1(n870), .A2(n869), .ZN(n871) );
  NAND2_X1 U969 ( .A1(n872), .A2(n871), .ZN(n877) );
  XNOR2_X1 U970 ( .A(G2067), .B(G26), .ZN(n874) );
  XNOR2_X1 U971 ( .A(G2072), .B(G33), .ZN(n873) );
  NOR2_X1 U972 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U973 ( .A(n875), .B(KEYINPUT119), .ZN(n876) );
  NOR2_X1 U974 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U975 ( .A(n878), .B(KEYINPUT53), .ZN(n879) );
  NOR2_X1 U976 ( .A1(n880), .A2(n879), .ZN(n883) );
  XOR2_X1 U977 ( .A(G2090), .B(KEYINPUT118), .Z(n881) );
  XNOR2_X1 U978 ( .A(G35), .B(n881), .ZN(n882) );
  NAND2_X1 U979 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U980 ( .A(n885), .B(n884), .ZN(n887) );
  INV_X1 U981 ( .A(G29), .ZN(n886) );
  NAND2_X1 U982 ( .A1(n887), .A2(n886), .ZN(n888) );
  NAND2_X1 U983 ( .A1(G11), .A2(n888), .ZN(n942) );
  XNOR2_X1 U984 ( .A(G16), .B(KEYINPUT56), .ZN(n910) );
  XNOR2_X1 U985 ( .A(G1966), .B(G168), .ZN(n890) );
  NAND2_X1 U986 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U987 ( .A(n891), .B(KEYINPUT57), .ZN(n908) );
  XNOR2_X1 U988 ( .A(n952), .B(G1341), .ZN(n906) );
  XNOR2_X1 U989 ( .A(n948), .B(G1348), .ZN(n893) );
  NAND2_X1 U990 ( .A1(n893), .A2(n892), .ZN(n895) );
  XNOR2_X1 U991 ( .A(G1971), .B(G303), .ZN(n894) );
  NOR2_X1 U992 ( .A1(n895), .A2(n894), .ZN(n901) );
  XNOR2_X1 U993 ( .A(G171), .B(G1961), .ZN(n897) );
  NAND2_X1 U994 ( .A1(n897), .A2(n896), .ZN(n899) );
  XNOR2_X1 U995 ( .A(G1956), .B(G299), .ZN(n898) );
  NOR2_X1 U996 ( .A1(n899), .A2(n898), .ZN(n900) );
  NAND2_X1 U997 ( .A1(n901), .A2(n900), .ZN(n902) );
  NOR2_X1 U998 ( .A1(n903), .A2(n902), .ZN(n904) );
  XNOR2_X1 U999 ( .A(KEYINPUT121), .B(n904), .ZN(n905) );
  NOR2_X1 U1000 ( .A1(n906), .A2(n905), .ZN(n907) );
  NAND2_X1 U1001 ( .A1(n908), .A2(n907), .ZN(n909) );
  NAND2_X1 U1002 ( .A1(n910), .A2(n909), .ZN(n940) );
  INV_X1 U1003 ( .A(G16), .ZN(n938) );
  XNOR2_X1 U1004 ( .A(G5), .B(n911), .ZN(n920) );
  XOR2_X1 U1005 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n918) );
  XNOR2_X1 U1006 ( .A(G1986), .B(G24), .ZN(n913) );
  XNOR2_X1 U1007 ( .A(G1971), .B(G22), .ZN(n912) );
  NOR2_X1 U1008 ( .A1(n913), .A2(n912), .ZN(n916) );
  XNOR2_X1 U1009 ( .A(G1976), .B(KEYINPUT125), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(n914), .B(G23), .ZN(n915) );
  NAND2_X1 U1011 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1012 ( .A(n918), .B(n917), .ZN(n919) );
  NAND2_X1 U1013 ( .A1(n920), .A2(n919), .ZN(n935) );
  XOR2_X1 U1014 ( .A(G1966), .B(G21), .Z(n933) );
  XNOR2_X1 U1015 ( .A(G1341), .B(G19), .ZN(n922) );
  XNOR2_X1 U1016 ( .A(G1981), .B(G6), .ZN(n921) );
  NOR2_X1 U1017 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1018 ( .A(KEYINPUT123), .B(n923), .Z(n927) );
  XNOR2_X1 U1019 ( .A(KEYINPUT59), .B(KEYINPUT124), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(n924), .B(G4), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(G1348), .B(n925), .ZN(n926) );
  NAND2_X1 U1022 ( .A1(n927), .A2(n926), .ZN(n930) );
  XNOR2_X1 U1023 ( .A(KEYINPUT122), .B(G1956), .ZN(n928) );
  XNOR2_X1 U1024 ( .A(G20), .B(n928), .ZN(n929) );
  NOR2_X1 U1025 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1026 ( .A(KEYINPUT60), .B(n931), .ZN(n932) );
  NAND2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1028 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1029 ( .A(KEYINPUT61), .B(n936), .ZN(n937) );
  NAND2_X1 U1030 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1031 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1032 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1033 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1034 ( .A(KEYINPUT62), .B(n945), .Z(G311) );
  XNOR2_X1 U1035 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1036 ( .A(G120), .ZN(G236) );
  INV_X1 U1037 ( .A(G108), .ZN(G238) );
  INV_X1 U1038 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1039 ( .A1(n947), .A2(n946), .ZN(G325) );
  INV_X1 U1040 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1041 ( .A(KEYINPUT114), .B(G286), .Z(n950) );
  XNOR2_X1 U1042 ( .A(G171), .B(n948), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(n950), .B(n949), .ZN(n954) );
  XNOR2_X1 U1044 ( .A(n952), .B(n951), .ZN(n953) );
  XNOR2_X1 U1045 ( .A(n954), .B(n953), .ZN(n955) );
  NOR2_X1 U1046 ( .A1(G37), .A2(n955), .ZN(G397) );
  XNOR2_X1 U1047 ( .A(G1966), .B(G1961), .ZN(n965) );
  XOR2_X1 U1048 ( .A(G1971), .B(G1956), .Z(n957) );
  XNOR2_X1 U1049 ( .A(G1996), .B(G1986), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(n957), .B(n956), .ZN(n961) );
  XOR2_X1 U1051 ( .A(KEYINPUT108), .B(G2474), .Z(n959) );
  XNOR2_X1 U1052 ( .A(G1991), .B(G1981), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(n959), .B(n958), .ZN(n960) );
  XOR2_X1 U1054 ( .A(n961), .B(n960), .Z(n963) );
  XNOR2_X1 U1055 ( .A(G1976), .B(KEYINPUT41), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(n963), .B(n962), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(n965), .B(n964), .ZN(G229) );
  XOR2_X1 U1058 ( .A(KEYINPUT107), .B(KEYINPUT106), .Z(n967) );
  XNOR2_X1 U1059 ( .A(G2072), .B(G2090), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(n967), .B(n966), .ZN(n971) );
  XOR2_X1 U1061 ( .A(KEYINPUT43), .B(G2678), .Z(n969) );
  XNOR2_X1 U1062 ( .A(G2067), .B(KEYINPUT42), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(n969), .B(n968), .ZN(n970) );
  XOR2_X1 U1064 ( .A(n971), .B(n970), .Z(n973) );
  XNOR2_X1 U1065 ( .A(G2096), .B(G2100), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(n973), .B(n972), .ZN(n975) );
  XOR2_X1 U1067 ( .A(G2078), .B(G2084), .Z(n974) );
  XNOR2_X1 U1068 ( .A(n975), .B(n974), .ZN(G227) );
  XNOR2_X1 U1069 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(n976), .B(KEYINPUT113), .ZN(n977) );
  XNOR2_X1 U1071 ( .A(n978), .B(n977), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(n980), .B(n979), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(G160), .B(G164), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(n982), .B(n981), .ZN(n983) );
  XOR2_X1 U1075 ( .A(n984), .B(n983), .Z(n987) );
  XNOR2_X1 U1076 ( .A(n985), .B(G162), .ZN(n986) );
  XNOR2_X1 U1077 ( .A(n987), .B(n986), .ZN(n1006) );
  XNOR2_X1 U1078 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n995) );
  NAND2_X1 U1079 ( .A1(n988), .A2(G142), .ZN(n989) );
  XNOR2_X1 U1080 ( .A(n989), .B(KEYINPUT110), .ZN(n992) );
  NAND2_X1 U1081 ( .A1(G106), .A2(n990), .ZN(n991) );
  NAND2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1083 ( .A(n993), .B(KEYINPUT45), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(n995), .B(n994), .ZN(n1002) );
  NAND2_X1 U1085 ( .A1(G118), .A2(n996), .ZN(n999) );
  NAND2_X1 U1086 ( .A1(G130), .A2(n997), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1088 ( .A(KEYINPUT109), .B(n1000), .Z(n1001) );
  NOR2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1090 ( .A(n1004), .B(n1003), .Z(n1005) );
  XNOR2_X1 U1091 ( .A(n1006), .B(n1005), .ZN(n1007) );
  NOR2_X1 U1092 ( .A1(G37), .A2(n1007), .ZN(G395) );
  NOR2_X1 U1093 ( .A1(G401), .A2(n1014), .ZN(n1011) );
  NOR2_X1 U1094 ( .A1(G229), .A2(G227), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(KEYINPUT49), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1096 ( .A1(G397), .A2(n1009), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1098 ( .A1(n1012), .A2(G395), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(n1013), .B(KEYINPUT115), .ZN(G225) );
  INV_X1 U1100 ( .A(G225), .ZN(G308) );
  INV_X1 U1101 ( .A(n1014), .ZN(G319) );
endmodule

