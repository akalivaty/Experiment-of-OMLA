//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 0 1 0 1 1 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n565,
    new_n566, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  XOR2_X1   g016(.A(KEYINPUT67), .B(G57), .Z(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT68), .Z(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G137), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n465), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AND2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(KEYINPUT69), .ZN(new_n480));
  INV_X1    g055(.A(G2105), .ZN(new_n481));
  XNOR2_X1  g056(.A(KEYINPUT3), .B(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G125), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n481), .B1(new_n483), .B2(new_n473), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n472), .B1(new_n480), .B2(new_n486), .ZN(G160));
  NAND2_X1  g062(.A1(new_n468), .A2(G136), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n481), .B1(new_n466), .B2(new_n467), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  OR2_X1    g065(.A1(G100), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G112), .C2(new_n481), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n488), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  NAND3_X1  g069(.A1(new_n482), .A2(G126), .A3(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(G114), .B2(new_n481), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g074(.A(G138), .B(new_n481), .C1(new_n474), .C2(new_n475), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n468), .A2(new_n502), .A3(G138), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n499), .B1(new_n501), .B2(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT70), .B1(new_n511), .B2(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n513), .A2(new_n514), .A3(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n506), .B1(KEYINPUT6), .B2(new_n511), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G50), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n510), .A2(new_n511), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n507), .A2(new_n508), .B1(KEYINPUT6), .B2(new_n511), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n522));
  AND3_X1   g097(.A1(new_n521), .A2(new_n522), .A3(new_n516), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n522), .B1(new_n521), .B2(new_n516), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n520), .B1(new_n525), .B2(G88), .ZN(G166));
  INV_X1    g101(.A(new_n518), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n531));
  AND2_X1   g106(.A1(G63), .A2(G651), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n530), .A2(new_n531), .B1(new_n509), .B2(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n525), .A2(G89), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(G168));
  NAND2_X1  g111(.A1(new_n525), .A2(G90), .ZN(new_n537));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  XOR2_X1   g113(.A(KEYINPUT5), .B(G543), .Z(new_n539));
  INV_X1    g114(.A(G64), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(G52), .A2(new_n527), .B1(new_n541), .B2(G651), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n537), .A2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n545), .B1(new_n507), .B2(new_n508), .ZN(new_n546));
  AND2_X1   g121(.A1(G68), .A2(G543), .ZN(new_n547));
  OR3_X1    g122(.A1(new_n546), .A2(KEYINPUT72), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g123(.A(KEYINPUT72), .B1(new_n546), .B2(new_n547), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n548), .A2(G651), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n527), .A2(G43), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n521), .A2(new_n516), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(KEYINPUT71), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n521), .A2(new_n516), .A3(new_n522), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(G81), .ZN(new_n556));
  OAI211_X1 g131(.A(new_n550), .B(new_n551), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(KEYINPUT73), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n525), .A2(G81), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT73), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n559), .A2(new_n560), .A3(new_n550), .A4(new_n551), .ZN(new_n561));
  AND2_X1   g136(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  NAND3_X1  g142(.A1(new_n516), .A2(G53), .A3(new_n517), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT9), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n553), .A2(G91), .A3(new_n554), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n509), .A2(G65), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  XOR2_X1   g147(.A(new_n572), .B(KEYINPUT74), .Z(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n569), .A2(new_n570), .A3(new_n574), .ZN(G299));
  NAND2_X1  g150(.A1(new_n534), .A2(new_n535), .ZN(G286));
  INV_X1    g151(.A(G166), .ZN(G303));
  OR2_X1    g152(.A1(new_n509), .A2(G74), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n527), .A2(G49), .B1(new_n578), .B2(G651), .ZN(new_n579));
  INV_X1    g154(.A(G87), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n555), .B2(new_n580), .ZN(G288));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n539), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(G48), .A2(new_n527), .B1(new_n584), .B2(G651), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n553), .A2(G86), .A3(new_n554), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT75), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n553), .A2(KEYINPUT75), .A3(G86), .A4(new_n554), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n586), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(G72), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G60), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n539), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(G47), .A2(new_n527), .B1(new_n595), .B2(G651), .ZN(new_n596));
  INV_X1    g171(.A(G85), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n555), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT76), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n598), .B(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  XOR2_X1   g176(.A(KEYINPUT77), .B(G66), .Z(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(new_n509), .B1(G79), .B2(G543), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n603), .A2(new_n511), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n527), .A2(G54), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n555), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n525), .A2(KEYINPUT10), .A3(G92), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n601), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n601), .B1(new_n611), .B2(G868), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  INV_X1    g189(.A(G299), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(G868), .B2(new_n615), .ZN(G297));
  OAI21_X1  g191(.A(new_n614), .B1(G868), .B2(new_n615), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n609), .A2(new_n610), .ZN(new_n620));
  INV_X1    g195(.A(new_n606), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(G868), .B1(new_n622), .B2(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n562), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n468), .A2(G135), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT79), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  INV_X1    g203(.A(G111), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(G2105), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(G123), .B2(new_n489), .ZN(new_n631));
  AND2_X1   g206(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(G2096), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n482), .A2(new_n470), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT78), .B(KEYINPUT13), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(G2100), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(G2100), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n633), .A2(G2096), .ZN(new_n641));
  NAND4_X1  g216(.A1(new_n634), .A2(new_n639), .A3(new_n640), .A4(new_n641), .ZN(G156));
  XOR2_X1   g217(.A(KEYINPUT15), .B(G2435), .Z(new_n643));
  XOR2_X1   g218(.A(KEYINPUT80), .B(G2438), .Z(new_n644));
  XOR2_X1   g219(.A(new_n643), .B(new_n644), .Z(new_n645));
  XNOR2_X1  g220(.A(G2427), .B(G2430), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(KEYINPUT14), .ZN(new_n648));
  AND2_X1   g223(.A1(new_n648), .A2(KEYINPUT81), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n648), .A2(KEYINPUT81), .ZN(new_n650));
  OAI22_X1  g225(.A1(new_n649), .A2(new_n650), .B1(new_n646), .B2(new_n645), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n653), .A2(new_n655), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT82), .ZN(new_n661));
  INV_X1    g236(.A(G14), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n656), .A2(new_n659), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n662), .B1(new_n663), .B2(new_n657), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(G401));
  INV_X1    g241(.A(KEYINPUT18), .ZN(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(KEYINPUT17), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n668), .A2(new_n669), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n667), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G2100), .ZN(new_n674));
  XOR2_X1   g249(.A(G2072), .B(G2078), .Z(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n670), .B2(KEYINPUT18), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G2096), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n674), .B(new_n677), .ZN(G227));
  XOR2_X1   g253(.A(G1971), .B(G1976), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  AND2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT20), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n681), .A2(new_n682), .ZN(new_n686));
  NOR3_X1   g261(.A1(new_n680), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(new_n680), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G1981), .B(G1986), .Z(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n690), .B(new_n691), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n689), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT83), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT84), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n693), .B(new_n696), .ZN(G229));
  XNOR2_X1  g272(.A(KEYINPUT96), .B(KEYINPUT26), .ZN(new_n698));
  AND3_X1   g273(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  AOI22_X1  g276(.A1(new_n700), .A2(new_n701), .B1(G105), .B2(new_n470), .ZN(new_n702));
  AOI22_X1  g277(.A1(G129), .A2(new_n489), .B1(new_n468), .B2(G141), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G29), .ZN(new_n706));
  NOR2_X1   g281(.A1(G29), .A2(G32), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(KEYINPUT97), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(KEYINPUT97), .B2(new_n706), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT27), .B(G1996), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G21), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G168), .B2(new_n712), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n711), .B1(G1966), .B2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT24), .ZN(new_n716));
  INV_X1    g291(.A(G34), .ZN(new_n717));
  AOI21_X1  g292(.A(G29), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(new_n716), .B2(new_n717), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(G160), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n721), .A2(G2084), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT98), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n714), .A2(G1966), .B1(G2084), .B2(new_n721), .ZN(new_n724));
  INV_X1    g299(.A(G1961), .ZN(new_n725));
  NOR2_X1   g300(.A1(G171), .A2(new_n712), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G5), .B2(new_n712), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n723), .B(new_n724), .C1(new_n725), .C2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n725), .ZN(new_n729));
  NOR2_X1   g304(.A1(G29), .A2(G35), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G162), .B2(G29), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT99), .B(KEYINPUT29), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n729), .B1(G2090), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT31), .B(G11), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT30), .B(G28), .Z(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(G29), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n632), .B2(G29), .ZN(new_n738));
  INV_X1    g313(.A(G2072), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n720), .A2(G33), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT95), .B(KEYINPUT25), .Z(new_n741));
  NAND3_X1  g316(.A1(new_n481), .A2(G103), .A3(G2104), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n468), .A2(G139), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n482), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n743), .B(new_n744), .C1(new_n481), .C2(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n740), .B1(new_n746), .B2(G29), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n738), .B1(new_n739), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n739), .B2(new_n747), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n720), .A2(G27), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G164), .B2(new_n720), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G2078), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n733), .B2(G2090), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n720), .A2(G26), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT28), .Z(new_n755));
  OAI21_X1  g330(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n756));
  INV_X1    g331(.A(G116), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(G2105), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT94), .ZN(new_n759));
  AOI22_X1  g334(.A1(G128), .A2(new_n489), .B1(new_n468), .B2(G140), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n755), .B1(new_n761), .B2(G29), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G2067), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n749), .A2(new_n753), .A3(new_n763), .ZN(new_n764));
  NOR4_X1   g339(.A1(new_n715), .A2(new_n728), .A3(new_n734), .A4(new_n764), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT89), .B(G16), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G20), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT23), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n615), .B2(new_n712), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(G1956), .Z(new_n770));
  NOR2_X1   g345(.A1(G4), .A2(G16), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n611), .B2(G16), .ZN(new_n772));
  INV_X1    g347(.A(G1348), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n765), .A2(new_n770), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n766), .A2(G19), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n562), .B2(new_n766), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT93), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1341), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n712), .A2(G23), .ZN(new_n782));
  INV_X1    g357(.A(G288), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n712), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT33), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1976), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n712), .A2(G6), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n591), .B2(new_n712), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT32), .B(G1981), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n788), .B(new_n789), .Z(new_n790));
  INV_X1    g365(.A(new_n766), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(G22), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G166), .B2(new_n791), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT91), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1971), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n786), .A2(new_n790), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n796), .A2(KEYINPUT34), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n791), .A2(G24), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n598), .B(KEYINPUT76), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(new_n791), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT90), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n802), .A2(G1986), .A3(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT35), .B(G1991), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT87), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT88), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT86), .ZN(new_n809));
  AOI22_X1  g384(.A1(G119), .A2(new_n489), .B1(new_n468), .B2(G131), .ZN(new_n810));
  OAI21_X1  g385(.A(KEYINPUT85), .B1(G95), .B2(G2105), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  NOR3_X1   g387(.A1(KEYINPUT85), .A2(G95), .A3(G2105), .ZN(new_n813));
  OAI221_X1 g388(.A(G2104), .B1(G107), .B2(new_n481), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  MUX2_X1   g390(.A(G25), .B(new_n815), .S(G29), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n809), .B(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(G1986), .B1(new_n802), .B2(new_n803), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n805), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT92), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT34), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n786), .A2(new_n821), .A3(new_n790), .A4(new_n795), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n819), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n820), .B1(new_n819), .B2(new_n822), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n797), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(KEYINPUT36), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n819), .A2(new_n822), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT92), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(new_n823), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT36), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n830), .A2(new_n831), .A3(new_n797), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n781), .B1(new_n827), .B2(new_n832), .ZN(G311));
  AOI21_X1  g408(.A(new_n831), .B1(new_n830), .B2(new_n797), .ZN(new_n834));
  INV_X1    g409(.A(new_n797), .ZN(new_n835));
  AOI211_X1 g410(.A(KEYINPUT36), .B(new_n835), .C1(new_n829), .C2(new_n823), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n780), .B1(new_n834), .B2(new_n836), .ZN(G150));
  NAND2_X1  g412(.A1(G80), .A2(G543), .ZN(new_n838));
  INV_X1    g413(.A(G67), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n539), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(G651), .ZN(new_n841));
  INV_X1    g416(.A(G55), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n842), .B2(new_n518), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(new_n525), .B2(G93), .ZN(new_n844));
  INV_X1    g419(.A(G860), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT37), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n611), .A2(G559), .ZN(new_n848));
  XNOR2_X1  g423(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n844), .B1(new_n558), .B2(new_n561), .ZN(new_n851));
  INV_X1    g426(.A(G93), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n555), .A2(new_n852), .ZN(new_n853));
  NOR3_X1   g428(.A1(new_n557), .A2(new_n853), .A3(new_n843), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n850), .B(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT39), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT101), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n845), .B1(new_n857), .B2(KEYINPUT39), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n847), .B1(new_n859), .B2(new_n860), .ZN(G145));
  XNOR2_X1  g436(.A(new_n746), .B(new_n704), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n489), .A2(G130), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n481), .A2(G118), .ZN(new_n864));
  OAI21_X1  g439(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n866), .B1(G142), .B2(new_n468), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n636), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n862), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n761), .B(G164), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n815), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n869), .B(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(G160), .B(G162), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n633), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n872), .A2(new_n874), .ZN(new_n876));
  NOR3_X1   g451(.A1(new_n875), .A2(new_n876), .A3(G37), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n877), .B(KEYINPUT40), .Z(G395));
  XNOR2_X1  g453(.A(new_n591), .B(G303), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(G290), .A2(G288), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n799), .A2(new_n783), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n880), .B1(new_n883), .B2(KEYINPUT104), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(KEYINPUT104), .B2(new_n883), .ZN(new_n885));
  OR3_X1    g460(.A1(new_n883), .A2(KEYINPUT104), .A3(new_n879), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(KEYINPUT42), .B1(new_n888), .B2(KEYINPUT105), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n622), .A2(new_n615), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n611), .A2(G299), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n890), .A2(KEYINPUT102), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT41), .ZN(new_n893));
  OR3_X1    g468(.A1(new_n611), .A2(KEYINPUT102), .A3(G299), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n895), .A2(KEYINPUT103), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n890), .A2(new_n891), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  AOI22_X1  g473(.A1(new_n895), .A2(KEYINPUT103), .B1(KEYINPUT41), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n622), .A2(G559), .ZN(new_n901));
  XOR2_X1   g476(.A(new_n855), .B(new_n901), .Z(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(new_n898), .B2(new_n902), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT42), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n887), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n889), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n904), .B1(new_n889), .B2(new_n907), .ZN(new_n909));
  OAI21_X1  g484(.A(G868), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n910), .B1(G868), .B2(new_n844), .ZN(G295));
  OAI21_X1  g486(.A(new_n910), .B1(G868), .B2(new_n844), .ZN(G331));
  XNOR2_X1  g487(.A(G168), .B(G301), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n855), .A2(KEYINPUT106), .A3(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(G286), .B(G301), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(new_n851), .B2(new_n854), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT106), .B1(new_n855), .B2(new_n913), .ZN(new_n918));
  NOR3_X1   g493(.A1(new_n917), .A2(new_n898), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n855), .A2(new_n913), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n916), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n919), .B1(new_n900), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(G37), .B1(new_n922), .B2(new_n888), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n917), .A2(new_n918), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n893), .B1(new_n892), .B2(new_n894), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI22_X1  g502(.A1(new_n925), .A2(new_n926), .B1(new_n893), .B2(new_n897), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n924), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n920), .A2(new_n897), .A3(new_n916), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n930), .B(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n887), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n923), .A2(KEYINPUT43), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n900), .A2(new_n921), .ZN(new_n935));
  INV_X1    g510(.A(new_n919), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(new_n887), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT43), .B1(new_n923), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT44), .B1(new_n934), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n942));
  INV_X1    g517(.A(G37), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n888), .A2(new_n935), .A3(new_n936), .ZN(new_n944));
  AND4_X1   g519(.A1(new_n942), .A2(new_n933), .A3(new_n943), .A4(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n942), .B1(new_n923), .B2(new_n938), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n941), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n940), .A2(new_n947), .ZN(G397));
  INV_X1    g523(.A(G2067), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n761), .B(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n950), .B(KEYINPUT110), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n705), .ZN(new_n952));
  INV_X1    g527(.A(G1996), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  XOR2_X1   g529(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(G164), .B2(G1384), .ZN(new_n956));
  INV_X1    g531(.A(new_n472), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n484), .A2(new_n485), .ZN(new_n958));
  AOI211_X1 g533(.A(KEYINPUT69), .B(new_n481), .C1(new_n483), .C2(new_n473), .ZN(new_n959));
  OAI211_X1 g534(.A(G40), .B(new_n957), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n956), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n952), .A2(new_n954), .A3(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n961), .A2(new_n953), .A3(new_n705), .ZN(new_n963));
  INV_X1    g538(.A(new_n961), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n815), .B(new_n807), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT111), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n962), .B(new_n963), .C1(new_n964), .C2(new_n966), .ZN(new_n967));
  OR2_X1    g542(.A1(G290), .A2(G1986), .ZN(new_n968));
  NAND2_X1  g543(.A1(G290), .A2(G1986), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n964), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G8), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n503), .A2(new_n501), .ZN(new_n973));
  INV_X1    g548(.A(G114), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n496), .B1(new_n974), .B2(G2105), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n975), .B1(G126), .B2(new_n489), .ZN(new_n976));
  AOI21_X1  g551(.A(G1384), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT50), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT113), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT113), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n980), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n960), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n977), .A2(new_n978), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT112), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT112), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n977), .A2(new_n985), .A3(new_n978), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G2090), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n982), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G1971), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n977), .A2(KEYINPUT45), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n956), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n990), .B1(new_n992), .B2(new_n960), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n972), .B1(new_n989), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(G166), .A2(new_n972), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT55), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G2084), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n982), .A2(new_n987), .A3(new_n998), .ZN(new_n999));
  OR2_X1    g574(.A1(new_n977), .A2(KEYINPUT45), .ZN(new_n1000));
  INV_X1    g575(.A(G40), .ZN(new_n1001));
  AOI211_X1 g576(.A(new_n1001), .B(new_n472), .C1(new_n480), .C2(new_n486), .ZN(new_n1002));
  INV_X1    g577(.A(new_n955), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n977), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1000), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1966), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n999), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1008), .A2(G8), .A3(G168), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n997), .A2(new_n1010), .A3(KEYINPUT63), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n973), .A2(new_n976), .ZN(new_n1012));
  INV_X1    g587(.A(G1384), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n960), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(new_n972), .ZN(new_n1016));
  INV_X1    g591(.A(G1981), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1017), .B1(new_n585), .B2(new_n587), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT75), .B1(new_n525), .B2(G86), .ZN(new_n1019));
  INV_X1    g594(.A(new_n590), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1017), .B(new_n585), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT117), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n591), .A2(KEYINPUT117), .A3(new_n1017), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1018), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1016), .B1(new_n1025), .B2(KEYINPUT49), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT49), .ZN(new_n1027));
  AOI211_X1 g602(.A(new_n1027), .B(new_n1018), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT118), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1018), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT117), .B1(new_n591), .B2(new_n1017), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n1027), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1025), .A2(KEYINPUT49), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1016), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1029), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n1039));
  XOR2_X1   g614(.A(KEYINPUT115), .B(G1976), .Z(new_n1040));
  OAI21_X1  g615(.A(new_n1039), .B1(new_n783), .B2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1041), .B(KEYINPUT116), .ZN(new_n1042));
  INV_X1    g617(.A(G1976), .ZN(new_n1043));
  OAI221_X1 g618(.A(G8), .B1(G288), .B2(new_n1043), .C1(new_n960), .C2(new_n1014), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1044), .A2(KEYINPUT114), .A3(KEYINPUT52), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT114), .B1(new_n1044), .B2(KEYINPUT52), .ZN(new_n1046));
  OAI22_X1  g621(.A1(new_n1042), .A2(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  OR2_X1    g623(.A1(new_n994), .A2(new_n996), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1011), .A2(new_n1038), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1014), .A2(KEYINPUT50), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1002), .A2(new_n983), .A3(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n993), .B1(G2090), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n996), .B1(new_n1054), .B2(G8), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1055), .B1(new_n996), .B2(new_n994), .ZN(new_n1056));
  AND4_X1   g631(.A1(new_n1038), .A2(new_n1048), .A3(new_n1056), .A4(new_n1010), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT63), .B1(new_n1057), .B2(KEYINPUT120), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT120), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1038), .A2(new_n1048), .A3(new_n1056), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1059), .B1(new_n1060), .B2(new_n1009), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1051), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1062));
  AOI211_X1 g637(.A(new_n997), .B(new_n1047), .C1(new_n1029), .C2(new_n1037), .ZN(new_n1063));
  NOR2_X1   g638(.A1(G288), .A2(G1976), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1016), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1065), .B1(new_n1033), .B2(new_n1027), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1036), .B1(new_n1066), .B2(new_n1035), .ZN(new_n1067));
  NOR3_X1   g642(.A1(new_n1026), .A2(KEYINPUT118), .A3(new_n1028), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1064), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  XOR2_X1   g646(.A(new_n1016), .B(KEYINPUT119), .Z(new_n1072));
  AOI21_X1  g647(.A(new_n1063), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n980), .B1(new_n1014), .B2(KEYINPUT50), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n977), .A2(KEYINPUT113), .A3(new_n978), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1002), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n986), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n985), .B1(new_n977), .B2(new_n978), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n725), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G2078), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT53), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n1005), .A2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1002), .A2(new_n1081), .A3(new_n956), .A4(new_n991), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1080), .A2(new_n1083), .A3(new_n1086), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n1087), .A2(G301), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n999), .A2(G168), .A3(new_n1007), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1089), .A2(new_n1090), .A3(G8), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1008), .A2(G286), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1092), .A2(G8), .A3(new_n1089), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1091), .B1(new_n1093), .B2(KEYINPUT51), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT62), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1088), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1093), .A2(KEYINPUT51), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1091), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT62), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT122), .B(KEYINPUT57), .ZN(new_n1101));
  XNOR2_X1  g676(.A(G299), .B(new_n1101), .ZN(new_n1102));
  XOR2_X1   g677(.A(KEYINPUT121), .B(G1956), .Z(new_n1103));
  NAND2_X1  g678(.A1(new_n1053), .A2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT123), .B(KEYINPUT56), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1105), .B(new_n739), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1002), .A2(new_n956), .A3(new_n991), .A4(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1102), .B1(new_n1104), .B2(new_n1107), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1104), .A2(new_n1102), .A3(new_n1107), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1109), .A2(new_n622), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n773), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1015), .A2(new_n949), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1108), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1111), .A2(KEYINPUT60), .A3(new_n1112), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n611), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1111), .A2(KEYINPUT60), .A3(new_n622), .A4(new_n1112), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT60), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1116), .A2(new_n1117), .B1(new_n1118), .B2(new_n1113), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT61), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(new_n1109), .B2(new_n1108), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1002), .A2(new_n953), .A3(new_n956), .A4(new_n991), .ZN(new_n1122));
  XNOR2_X1  g697(.A(KEYINPUT124), .B(KEYINPUT58), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1123), .B(G1341), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n960), .B2(new_n1014), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT125), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1127), .B1(new_n1128), .B2(KEYINPUT59), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1129), .B1(new_n1127), .B2(KEYINPUT59), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1126), .A2(new_n562), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1129), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1132), .B1(new_n1126), .B2(new_n562), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1102), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1103), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n960), .B1(KEYINPUT50), .B2(new_n1014), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1136), .B1(new_n1137), .B2(new_n983), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1107), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1135), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1104), .A2(new_n1102), .A3(new_n1107), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1140), .A2(KEYINPUT61), .A3(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1121), .A2(new_n1134), .A3(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1114), .B1(new_n1119), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT54), .ZN(new_n1145));
  XNOR2_X1  g720(.A(G301), .B(new_n1145), .ZN(new_n1146));
  NOR4_X1   g721(.A1(new_n472), .A2(new_n484), .A3(new_n1001), .A4(new_n1082), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n956), .A2(new_n991), .A3(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1080), .A2(new_n1086), .A3(new_n1146), .A4(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(new_n1087), .B2(new_n1146), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1150), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1151));
  AOI22_X1  g726(.A1(new_n1096), .A2(new_n1100), .B1(new_n1144), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1073), .B1(new_n1152), .B2(new_n1060), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n971), .B1(new_n1062), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n952), .A2(new_n961), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n961), .A2(new_n953), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1156), .B(KEYINPUT46), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(new_n1158), .B(KEYINPUT47), .Z(new_n1159));
  INV_X1    g734(.A(KEYINPUT127), .ZN(new_n1160));
  AND2_X1   g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n968), .A2(new_n964), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1163), .B(KEYINPUT48), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1164), .A2(new_n967), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n962), .A2(new_n963), .ZN(new_n1166));
  OR2_X1    g741(.A1(new_n815), .A2(new_n807), .ZN(new_n1167));
  OAI22_X1  g742(.A1(new_n1166), .A2(new_n1167), .B1(G2067), .B2(new_n761), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1168), .A2(new_n961), .ZN(new_n1169));
  NOR4_X1   g744(.A1(new_n1161), .A2(new_n1162), .A3(new_n1165), .A4(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1154), .A2(new_n1170), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g746(.A1(new_n877), .A2(new_n462), .A3(G227), .A4(G229), .ZN(new_n1173));
  OAI211_X1 g747(.A(new_n665), .B(new_n1173), .C1(new_n945), .C2(new_n946), .ZN(G225));
  INV_X1    g748(.A(G225), .ZN(G308));
endmodule


