

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594;

  XNOR2_X1 U326 ( .A(n450), .B(n449), .ZN(n451) );
  NOR2_X1 U327 ( .A1(n578), .A2(n442), .ZN(n559) );
  XNOR2_X1 U328 ( .A(KEYINPUT102), .B(KEYINPUT37), .ZN(n455) );
  XNOR2_X1 U329 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U330 ( .A(n483), .B(KEYINPUT123), .ZN(n484) );
  XNOR2_X1 U331 ( .A(n345), .B(n344), .ZN(n569) );
  NOR2_X1 U332 ( .A1(n502), .A2(n515), .ZN(n508) );
  XOR2_X1 U333 ( .A(KEYINPUT93), .B(n414), .Z(n294) );
  XOR2_X1 U334 ( .A(n467), .B(KEYINPUT45), .Z(n295) );
  XOR2_X1 U335 ( .A(G99GAT), .B(KEYINPUT78), .Z(n296) );
  XOR2_X1 U336 ( .A(n425), .B(n424), .Z(n297) );
  XOR2_X1 U337 ( .A(KEYINPUT54), .B(n481), .Z(n298) );
  XNOR2_X1 U338 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U339 ( .A(n427), .B(n296), .ZN(n428) );
  INV_X1 U340 ( .A(KEYINPUT98), .ZN(n449) );
  XOR2_X1 U341 ( .A(n335), .B(KEYINPUT72), .Z(n337) );
  XNOR2_X1 U342 ( .A(n429), .B(n428), .ZN(n433) );
  NOR2_X1 U343 ( .A1(n528), .A2(n298), .ZN(n576) );
  XNOR2_X1 U344 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U345 ( .A(n400), .B(n399), .ZN(n402) );
  XNOR2_X1 U346 ( .A(n485), .B(n484), .ZN(n486) );
  NOR2_X1 U347 ( .A1(n578), .A2(n577), .ZN(n589) );
  INV_X1 U348 ( .A(G29GAT), .ZN(n462) );
  XNOR2_X1 U349 ( .A(n493), .B(G190GAT), .ZN(n494) );
  XNOR2_X1 U350 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U351 ( .A(n495), .B(n494), .ZN(G1351GAT) );
  XNOR2_X1 U352 ( .A(n461), .B(n460), .ZN(G1330GAT) );
  XOR2_X1 U353 ( .A(G113GAT), .B(G15GAT), .Z(n300) );
  XNOR2_X1 U354 ( .A(G197GAT), .B(G141GAT), .ZN(n299) );
  XNOR2_X1 U355 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U356 ( .A(KEYINPUT64), .B(KEYINPUT65), .Z(n302) );
  XNOR2_X1 U357 ( .A(G169GAT), .B(G8GAT), .ZN(n301) );
  XNOR2_X1 U358 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U359 ( .A(n304), .B(n303), .ZN(n316) );
  XOR2_X1 U360 ( .A(G1GAT), .B(KEYINPUT67), .Z(n358) );
  XOR2_X1 U361 ( .A(G22GAT), .B(G50GAT), .Z(n306) );
  XNOR2_X1 U362 ( .A(G43GAT), .B(G36GAT), .ZN(n305) );
  XNOR2_X1 U363 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U364 ( .A(n358), .B(n307), .Z(n309) );
  NAND2_X1 U365 ( .A1(G229GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U366 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U367 ( .A(n310), .B(KEYINPUT30), .Z(n314) );
  XOR2_X1 U368 ( .A(G29GAT), .B(KEYINPUT7), .Z(n312) );
  XNOR2_X1 U369 ( .A(KEYINPUT66), .B(KEYINPUT8), .ZN(n311) );
  XNOR2_X1 U370 ( .A(n312), .B(n311), .ZN(n334) );
  XNOR2_X1 U371 ( .A(n334), .B(KEYINPUT29), .ZN(n313) );
  XNOR2_X1 U372 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U373 ( .A(n316), .B(n315), .Z(n560) );
  INV_X1 U374 ( .A(n560), .ZN(n579) );
  XNOR2_X1 U375 ( .A(G57GAT), .B(KEYINPUT68), .ZN(n317) );
  XOR2_X1 U376 ( .A(n317), .B(KEYINPUT13), .Z(n348) );
  XOR2_X1 U377 ( .A(G92GAT), .B(G85GAT), .Z(n319) );
  XNOR2_X1 U378 ( .A(G99GAT), .B(G106GAT), .ZN(n318) );
  XNOR2_X1 U379 ( .A(n319), .B(n318), .ZN(n339) );
  XNOR2_X1 U380 ( .A(n348), .B(n339), .ZN(n324) );
  XNOR2_X1 U381 ( .A(G78GAT), .B(KEYINPUT70), .ZN(n320) );
  XNOR2_X1 U382 ( .A(n320), .B(G148GAT), .ZN(n415) );
  XOR2_X1 U383 ( .A(G64GAT), .B(KEYINPUT71), .Z(n322) );
  XNOR2_X1 U384 ( .A(G176GAT), .B(G204GAT), .ZN(n321) );
  XNOR2_X1 U385 ( .A(n322), .B(n321), .ZN(n396) );
  XNOR2_X1 U386 ( .A(n415), .B(n396), .ZN(n323) );
  XNOR2_X1 U387 ( .A(n324), .B(n323), .ZN(n331) );
  XOR2_X1 U388 ( .A(G120GAT), .B(G71GAT), .Z(n427) );
  XOR2_X1 U389 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n326) );
  XNOR2_X1 U390 ( .A(KEYINPUT69), .B(KEYINPUT32), .ZN(n325) );
  XNOR2_X1 U391 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U392 ( .A(n427), .B(n327), .Z(n329) );
  NAND2_X1 U393 ( .A1(G230GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U394 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U395 ( .A(n331), .B(n330), .Z(n466) );
  NAND2_X1 U396 ( .A1(n579), .A2(n466), .ZN(n502) );
  INV_X1 U397 ( .A(KEYINPUT36), .ZN(n346) );
  XOR2_X1 U398 ( .A(G36GAT), .B(G218GAT), .Z(n397) );
  AND2_X1 U399 ( .A1(G232GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U400 ( .A(n397), .B(n332), .ZN(n333) );
  XOR2_X1 U401 ( .A(G50GAT), .B(G162GAT), .Z(n405) );
  XNOR2_X1 U402 ( .A(n405), .B(KEYINPUT74), .ZN(n336) );
  XNOR2_X1 U403 ( .A(n337), .B(n336), .ZN(n345) );
  XNOR2_X1 U404 ( .A(G43GAT), .B(G190GAT), .ZN(n338) );
  XNOR2_X1 U405 ( .A(n338), .B(G134GAT), .ZN(n435) );
  XNOR2_X1 U406 ( .A(n435), .B(n339), .ZN(n343) );
  XOR2_X1 U407 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n341) );
  XNOR2_X1 U408 ( .A(KEYINPUT73), .B(KEYINPUT10), .ZN(n340) );
  XOR2_X1 U409 ( .A(n341), .B(n340), .Z(n342) );
  XNOR2_X1 U410 ( .A(n569), .B(KEYINPUT75), .ZN(n491) );
  XNOR2_X1 U411 ( .A(n346), .B(n491), .ZN(n591) );
  XNOR2_X1 U412 ( .A(G15GAT), .B(G183GAT), .ZN(n347) );
  XNOR2_X1 U413 ( .A(n347), .B(G127GAT), .ZN(n434) );
  XNOR2_X1 U414 ( .A(n434), .B(n348), .ZN(n362) );
  XOR2_X1 U415 ( .A(G8GAT), .B(G211GAT), .Z(n401) );
  XOR2_X1 U416 ( .A(G22GAT), .B(G155GAT), .Z(n404) );
  XOR2_X1 U417 ( .A(n401), .B(n404), .Z(n350) );
  NAND2_X1 U418 ( .A1(G231GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U419 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U420 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n352) );
  XNOR2_X1 U421 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n351) );
  XNOR2_X1 U422 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U423 ( .A(n354), .B(n353), .Z(n360) );
  XOR2_X1 U424 ( .A(KEYINPUT12), .B(G64GAT), .Z(n356) );
  XNOR2_X1 U425 ( .A(G71GAT), .B(G78GAT), .ZN(n355) );
  XNOR2_X1 U426 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U427 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U428 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U429 ( .A(n362), .B(n361), .Z(n587) );
  INV_X1 U430 ( .A(n587), .ZN(n498) );
  XOR2_X1 U431 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n364) );
  XNOR2_X1 U432 ( .A(G120GAT), .B(G57GAT), .ZN(n363) );
  XNOR2_X1 U433 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U434 ( .A(KEYINPUT73), .B(G155GAT), .Z(n366) );
  XNOR2_X1 U435 ( .A(G127GAT), .B(G148GAT), .ZN(n365) );
  XNOR2_X1 U436 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U437 ( .A(n368), .B(n367), .ZN(n387) );
  XOR2_X1 U438 ( .A(KEYINPUT88), .B(KEYINPUT6), .Z(n370) );
  XNOR2_X1 U439 ( .A(KEYINPUT89), .B(KEYINPUT1), .ZN(n369) );
  XNOR2_X1 U440 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U441 ( .A(KEYINPUT5), .B(KEYINPUT92), .Z(n372) );
  XNOR2_X1 U442 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n371) );
  XNOR2_X1 U443 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U444 ( .A(n374), .B(n373), .Z(n385) );
  XOR2_X1 U445 ( .A(KEYINPUT2), .B(KEYINPUT87), .Z(n376) );
  XNOR2_X1 U446 ( .A(KEYINPUT3), .B(KEYINPUT86), .ZN(n375) );
  XNOR2_X1 U447 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U448 ( .A(G141GAT), .B(n377), .Z(n422) );
  XOR2_X1 U449 ( .A(G113GAT), .B(KEYINPUT0), .Z(n424) );
  XOR2_X1 U450 ( .A(G85GAT), .B(G162GAT), .Z(n379) );
  XNOR2_X1 U451 ( .A(G29GAT), .B(G134GAT), .ZN(n378) );
  XNOR2_X1 U452 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U453 ( .A(n424), .B(n380), .Z(n382) );
  NAND2_X1 U454 ( .A1(G225GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U455 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U456 ( .A(n422), .B(n383), .ZN(n384) );
  XNOR2_X1 U457 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U458 ( .A(n387), .B(n386), .Z(n541) );
  INV_X1 U459 ( .A(n541), .ZN(n528) );
  XNOR2_X1 U460 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n388) );
  XNOR2_X1 U461 ( .A(n388), .B(KEYINPUT85), .ZN(n414) );
  NAND2_X1 U462 ( .A1(G226GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U463 ( .A(n294), .B(n389), .ZN(n393) );
  XOR2_X1 U464 ( .A(KEYINPUT94), .B(G92GAT), .Z(n391) );
  XNOR2_X1 U465 ( .A(G190GAT), .B(G183GAT), .ZN(n390) );
  XNOR2_X1 U466 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U467 ( .A(n393), .B(n392), .Z(n400) );
  XOR2_X1 U468 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n395) );
  XNOR2_X1 U469 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n394) );
  XNOR2_X1 U470 ( .A(n395), .B(n394), .ZN(n425) );
  XNOR2_X1 U471 ( .A(n425), .B(n396), .ZN(n398) );
  XOR2_X1 U472 ( .A(n402), .B(n401), .Z(n480) );
  INV_X1 U473 ( .A(n480), .ZN(n531) );
  XOR2_X1 U474 ( .A(KEYINPUT27), .B(KEYINPUT95), .Z(n403) );
  XOR2_X1 U475 ( .A(n531), .B(n403), .Z(n442) );
  XOR2_X1 U476 ( .A(G106GAT), .B(G218GAT), .Z(n407) );
  XNOR2_X1 U477 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U478 ( .A(n407), .B(n406), .ZN(n419) );
  XOR2_X1 U479 ( .A(KEYINPUT84), .B(KEYINPUT24), .Z(n409) );
  XNOR2_X1 U480 ( .A(G204GAT), .B(KEYINPUT23), .ZN(n408) );
  XNOR2_X1 U481 ( .A(n409), .B(n408), .ZN(n413) );
  XOR2_X1 U482 ( .A(G211GAT), .B(KEYINPUT22), .Z(n411) );
  XNOR2_X1 U483 ( .A(KEYINPUT83), .B(KEYINPUT82), .ZN(n410) );
  XNOR2_X1 U484 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U485 ( .A(n413), .B(n412), .Z(n417) );
  XNOR2_X1 U486 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U487 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U488 ( .A(n419), .B(n418), .Z(n421) );
  NAND2_X1 U489 ( .A1(G228GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U490 ( .A(n421), .B(n420), .ZN(n423) );
  XOR2_X1 U491 ( .A(n423), .B(n422), .Z(n482) );
  XOR2_X1 U492 ( .A(n482), .B(KEYINPUT28), .Z(n536) );
  OR2_X1 U493 ( .A1(n442), .A2(n536), .ZN(n544) );
  NAND2_X1 U494 ( .A1(G227GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U495 ( .A(n297), .B(n426), .ZN(n429) );
  XOR2_X1 U496 ( .A(G176GAT), .B(KEYINPUT80), .Z(n431) );
  XNOR2_X1 U497 ( .A(KEYINPUT79), .B(KEYINPUT20), .ZN(n430) );
  XNOR2_X1 U498 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U499 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U500 ( .A(n435), .B(n434), .Z(n436) );
  XNOR2_X1 U501 ( .A(n437), .B(n436), .ZN(n443) );
  INV_X1 U502 ( .A(n443), .ZN(n542) );
  XOR2_X1 U503 ( .A(KEYINPUT81), .B(n542), .Z(n438) );
  NOR2_X1 U504 ( .A1(n544), .A2(n438), .ZN(n439) );
  NAND2_X1 U505 ( .A1(n528), .A2(n439), .ZN(n440) );
  XNOR2_X1 U506 ( .A(KEYINPUT96), .B(n440), .ZN(n452) );
  NOR2_X1 U507 ( .A1(n482), .A2(n542), .ZN(n441) );
  XOR2_X1 U508 ( .A(KEYINPUT26), .B(n441), .Z(n578) );
  NOR2_X1 U509 ( .A1(n443), .A2(n480), .ZN(n444) );
  XNOR2_X1 U510 ( .A(n444), .B(KEYINPUT97), .ZN(n445) );
  NAND2_X1 U511 ( .A1(n445), .A2(n482), .ZN(n446) );
  XNOR2_X1 U512 ( .A(n446), .B(KEYINPUT25), .ZN(n447) );
  NOR2_X1 U513 ( .A1(n559), .A2(n447), .ZN(n448) );
  NOR2_X1 U514 ( .A1(n528), .A2(n448), .ZN(n450) );
  NAND2_X1 U515 ( .A1(n452), .A2(n451), .ZN(n500) );
  NAND2_X1 U516 ( .A1(n498), .A2(n500), .ZN(n453) );
  XOR2_X1 U517 ( .A(n453), .B(KEYINPUT101), .Z(n454) );
  NOR2_X1 U518 ( .A1(n591), .A2(n454), .ZN(n456) );
  XNOR2_X1 U519 ( .A(n456), .B(n455), .ZN(n527) );
  NOR2_X1 U520 ( .A1(n502), .A2(n527), .ZN(n457) );
  XNOR2_X1 U521 ( .A(n457), .B(KEYINPUT38), .ZN(n511) );
  NAND2_X1 U522 ( .A1(n511), .A2(n542), .ZN(n461) );
  XOR2_X1 U523 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n459) );
  XNOR2_X1 U524 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n458) );
  NAND2_X1 U525 ( .A1(n528), .A2(n511), .ZN(n465) );
  XOR2_X1 U526 ( .A(KEYINPUT39), .B(KEYINPUT103), .Z(n463) );
  XNOR2_X1 U527 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U528 ( .A(n465), .B(n464), .ZN(G1328GAT) );
  INV_X1 U529 ( .A(KEYINPUT118), .ZN(n469) );
  INV_X1 U530 ( .A(n466), .ZN(n584) );
  NOR2_X1 U531 ( .A1(n498), .A2(n591), .ZN(n467) );
  NOR2_X1 U532 ( .A1(n584), .A2(n295), .ZN(n468) );
  XNOR2_X1 U533 ( .A(n469), .B(n468), .ZN(n470) );
  NOR2_X1 U534 ( .A1(n579), .A2(n470), .ZN(n478) );
  XOR2_X1 U535 ( .A(KEYINPUT116), .B(KEYINPUT46), .Z(n472) );
  XOR2_X1 U536 ( .A(KEYINPUT41), .B(n584), .Z(n562) );
  NAND2_X1 U537 ( .A1(n579), .A2(n562), .ZN(n471) );
  XNOR2_X1 U538 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U539 ( .A(KEYINPUT115), .B(n587), .Z(n573) );
  NOR2_X1 U540 ( .A1(n473), .A2(n573), .ZN(n474) );
  NAND2_X1 U541 ( .A1(n569), .A2(n474), .ZN(n475) );
  XNOR2_X1 U542 ( .A(KEYINPUT117), .B(n475), .ZN(n476) );
  XOR2_X1 U543 ( .A(n476), .B(KEYINPUT47), .Z(n477) );
  NOR2_X1 U544 ( .A1(n478), .A2(n477), .ZN(n479) );
  XNOR2_X1 U545 ( .A(KEYINPUT48), .B(n479), .ZN(n540) );
  NOR2_X1 U546 ( .A1(n480), .A2(n540), .ZN(n481) );
  AND2_X1 U547 ( .A1(n576), .A2(n482), .ZN(n485) );
  INV_X1 U548 ( .A(KEYINPUT55), .ZN(n483) );
  NOR2_X1 U549 ( .A1(n443), .A2(n486), .ZN(n574) );
  XOR2_X1 U550 ( .A(KEYINPUT107), .B(n562), .Z(n546) );
  NAND2_X1 U551 ( .A1(n574), .A2(n546), .ZN(n490) );
  XOR2_X1 U552 ( .A(G176GAT), .B(KEYINPUT56), .Z(n488) );
  XNOR2_X1 U553 ( .A(KEYINPUT57), .B(KEYINPUT124), .ZN(n487) );
  XNOR2_X1 U554 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U555 ( .A(n490), .B(n489), .ZN(G1349GAT) );
  INV_X1 U556 ( .A(n491), .ZN(n492) );
  INV_X1 U557 ( .A(n492), .ZN(n553) );
  NAND2_X1 U558 ( .A1(n574), .A2(n553), .ZN(n495) );
  XOR2_X1 U559 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n493) );
  XNOR2_X1 U560 ( .A(G1GAT), .B(KEYINPUT100), .ZN(n496) );
  XNOR2_X1 U561 ( .A(n496), .B(KEYINPUT34), .ZN(n497) );
  XOR2_X1 U562 ( .A(KEYINPUT99), .B(n497), .Z(n504) );
  NOR2_X1 U563 ( .A1(n498), .A2(n553), .ZN(n499) );
  XNOR2_X1 U564 ( .A(n499), .B(KEYINPUT16), .ZN(n501) );
  NAND2_X1 U565 ( .A1(n501), .A2(n500), .ZN(n515) );
  NAND2_X1 U566 ( .A1(n508), .A2(n528), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(G1324GAT) );
  NAND2_X1 U568 ( .A1(n508), .A2(n531), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n505), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U570 ( .A(G15GAT), .B(KEYINPUT35), .Z(n507) );
  NAND2_X1 U571 ( .A1(n508), .A2(n542), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n507), .B(n506), .ZN(G1326GAT) );
  NAND2_X1 U573 ( .A1(n508), .A2(n536), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n509), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U575 ( .A1(n531), .A2(n511), .ZN(n510) );
  XNOR2_X1 U576 ( .A(G36GAT), .B(n510), .ZN(G1329GAT) );
  NAND2_X1 U577 ( .A1(n511), .A2(n536), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n512), .B(KEYINPUT106), .ZN(n513) );
  XNOR2_X1 U579 ( .A(G50GAT), .B(n513), .ZN(G1331GAT) );
  XNOR2_X1 U580 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n517) );
  NAND2_X1 U581 ( .A1(n546), .A2(n560), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n514), .B(KEYINPUT108), .ZN(n526) );
  NOR2_X1 U583 ( .A1(n526), .A2(n515), .ZN(n521) );
  NAND2_X1 U584 ( .A1(n528), .A2(n521), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n517), .B(n516), .ZN(G1332GAT) );
  XOR2_X1 U586 ( .A(G64GAT), .B(KEYINPUT109), .Z(n519) );
  NAND2_X1 U587 ( .A1(n521), .A2(n531), .ZN(n518) );
  XNOR2_X1 U588 ( .A(n519), .B(n518), .ZN(G1333GAT) );
  NAND2_X1 U589 ( .A1(n542), .A2(n521), .ZN(n520) );
  XNOR2_X1 U590 ( .A(n520), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n523) );
  NAND2_X1 U592 ( .A1(n521), .A2(n536), .ZN(n522) );
  XNOR2_X1 U593 ( .A(n523), .B(n522), .ZN(n525) );
  XOR2_X1 U594 ( .A(G78GAT), .B(KEYINPUT111), .Z(n524) );
  XNOR2_X1 U595 ( .A(n525), .B(n524), .ZN(G1335GAT) );
  NOR2_X1 U596 ( .A1(n527), .A2(n526), .ZN(n537) );
  NAND2_X1 U597 ( .A1(n537), .A2(n528), .ZN(n529) );
  XNOR2_X1 U598 ( .A(n529), .B(KEYINPUT112), .ZN(n530) );
  XNOR2_X1 U599 ( .A(G85GAT), .B(n530), .ZN(G1336GAT) );
  XOR2_X1 U600 ( .A(G92GAT), .B(KEYINPUT113), .Z(n533) );
  NAND2_X1 U601 ( .A1(n537), .A2(n531), .ZN(n532) );
  XNOR2_X1 U602 ( .A(n533), .B(n532), .ZN(G1337GAT) );
  NAND2_X1 U603 ( .A1(n542), .A2(n537), .ZN(n534) );
  XNOR2_X1 U604 ( .A(n534), .B(KEYINPUT114), .ZN(n535) );
  XNOR2_X1 U605 ( .A(G99GAT), .B(n535), .ZN(G1338GAT) );
  NAND2_X1 U606 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n538), .B(KEYINPUT44), .ZN(n539) );
  XNOR2_X1 U608 ( .A(G106GAT), .B(n539), .ZN(G1339GAT) );
  NOR2_X1 U609 ( .A1(n541), .A2(n540), .ZN(n558) );
  NAND2_X1 U610 ( .A1(n558), .A2(n542), .ZN(n543) );
  NOR2_X1 U611 ( .A1(n544), .A2(n543), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n554), .A2(n579), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n545), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT49), .B(KEYINPUT119), .Z(n548) );
  NAND2_X1 U615 ( .A1(n554), .A2(n546), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U617 ( .A(G120GAT), .B(n549), .Z(G1341GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT50), .B(KEYINPUT120), .Z(n551) );
  NAND2_X1 U619 ( .A1(n554), .A2(n573), .ZN(n550) );
  XNOR2_X1 U620 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U621 ( .A(G127GAT), .B(n552), .Z(G1342GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT121), .B(KEYINPUT51), .Z(n556) );
  NAND2_X1 U623 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U625 ( .A(G134GAT), .B(n557), .Z(G1343GAT) );
  NAND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n568) );
  NOR2_X1 U627 ( .A1(n560), .A2(n568), .ZN(n561) );
  XOR2_X1 U628 ( .A(G141GAT), .B(n561), .Z(G1344GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n564) );
  INV_X1 U630 ( .A(n568), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n566), .A2(n562), .ZN(n563) );
  XNOR2_X1 U632 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U633 ( .A(G148GAT), .B(n565), .ZN(G1345GAT) );
  NAND2_X1 U634 ( .A1(n566), .A2(n587), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n567), .B(G155GAT), .ZN(G1346GAT) );
  NOR2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U637 ( .A(KEYINPUT122), .B(n570), .Z(n571) );
  XNOR2_X1 U638 ( .A(G162GAT), .B(n571), .ZN(G1347GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n579), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n572), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n575), .B(G183GAT), .ZN(G1350GAT) );
  INV_X1 U643 ( .A(n576), .ZN(n577) );
  NAND2_X1 U644 ( .A1(n589), .A2(n579), .ZN(n583) );
  XOR2_X1 U645 ( .A(KEYINPUT59), .B(KEYINPUT126), .Z(n581) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1352GAT) );
  XOR2_X1 U649 ( .A(G204GAT), .B(KEYINPUT61), .Z(n586) );
  NAND2_X1 U650 ( .A1(n589), .A2(n584), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  NAND2_X1 U652 ( .A1(n587), .A2(n589), .ZN(n588) );
  XNOR2_X1 U653 ( .A(G211GAT), .B(n588), .ZN(G1354GAT) );
  INV_X1 U654 ( .A(n589), .ZN(n590) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n593) );
  XNOR2_X1 U656 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(n594), .B(G218GAT), .ZN(G1355GAT) );
endmodule

