//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G137), .ZN(new_n188));
  AND2_X1   g002(.A1(KEYINPUT66), .A2(G134), .ZN(new_n189));
  NOR2_X1   g003(.A1(KEYINPUT66), .A2(G134), .ZN(new_n190));
  OAI211_X1 g004(.A(new_n187), .B(new_n188), .C1(new_n189), .C2(new_n190), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n187), .B1(G134), .B2(new_n188), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n189), .A2(new_n190), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G137), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G131), .ZN(new_n198));
  AOI21_X1  g012(.A(G131), .B1(new_n195), .B2(G137), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n194), .A2(new_n199), .A3(KEYINPUT67), .ZN(new_n200));
  AOI21_X1  g014(.A(KEYINPUT67), .B1(new_n194), .B2(new_n199), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n198), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT0), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(new_n204), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n206), .B(new_n207), .C1(new_n209), .C2(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT65), .B1(new_n208), .B2(G146), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(new_n210), .A3(G143), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n208), .A2(G146), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n205), .A2(new_n213), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n202), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G134), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G137), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n222), .B1(new_n195), .B2(G137), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n224), .B1(G143), .B2(new_n210), .ZN(new_n225));
  OAI22_X1  g039(.A1(new_n225), .A2(new_n204), .B1(new_n209), .B2(new_n211), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n213), .A2(new_n215), .A3(new_n216), .A4(new_n227), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n223), .A2(G131), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(new_n200), .B2(new_n201), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT70), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n232), .B(new_n229), .C1(new_n200), .C2(new_n201), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n220), .A2(new_n231), .A3(KEYINPUT30), .A4(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G131), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n235), .B1(new_n194), .B2(new_n196), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n221), .ZN(new_n239));
  NAND2_X1  g053(.A1(KEYINPUT66), .A2(G134), .ZN(new_n240));
  AOI21_X1  g054(.A(G137), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n192), .B1(new_n241), .B2(new_n187), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n240), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n235), .B1(new_n243), .B2(new_n188), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n237), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n194), .A2(new_n199), .A3(KEYINPUT67), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n236), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n230), .B1(new_n247), .B2(new_n218), .ZN(new_n248));
  XOR2_X1   g062(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OR2_X1    g064(.A1(KEYINPUT2), .A2(G113), .ZN(new_n251));
  AND3_X1   g065(.A1(KEYINPUT68), .A2(KEYINPUT2), .A3(G113), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G119), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G116), .ZN(new_n256));
  INV_X1    g070(.A(G116), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G119), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n254), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(G116), .B(G119), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n261), .B(new_n251), .C1(new_n253), .C2(new_n252), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n260), .A2(new_n262), .A3(KEYINPUT69), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n254), .A2(new_n264), .A3(new_n259), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n234), .A2(new_n250), .A3(new_n267), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n220), .A2(new_n231), .A3(new_n266), .A4(new_n233), .ZN(new_n269));
  NOR2_X1   g083(.A1(G237), .A2(G953), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G210), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n271), .B(KEYINPUT27), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT26), .B(G101), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n272), .B(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT31), .B1(new_n268), .B2(new_n275), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n266), .B(new_n230), .C1(new_n247), .C2(new_n218), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT28), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n248), .A2(new_n267), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n279), .B(new_n280), .C1(new_n269), .C2(new_n278), .ZN(new_n281));
  INV_X1    g095(.A(new_n274), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n234), .A2(new_n250), .A3(new_n267), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT31), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n284), .A2(new_n285), .A3(new_n274), .A4(new_n269), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n276), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(G472), .A2(G902), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT71), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT32), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n287), .A2(KEYINPUT71), .A3(new_n288), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n287), .A2(KEYINPUT32), .A3(new_n288), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G472), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n281), .A2(new_n274), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n284), .A2(new_n282), .A3(new_n269), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT29), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n279), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n220), .A2(new_n231), .A3(new_n233), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n267), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n269), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n303), .B1(new_n306), .B2(KEYINPUT28), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n282), .A2(new_n301), .ZN(new_n308));
  AOI21_X1  g122(.A(G902), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n297), .B1(new_n302), .B2(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n296), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n294), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT25), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT16), .ZN(new_n314));
  INV_X1    g128(.A(G140), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(new_n315), .A3(G125), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(G125), .ZN(new_n317));
  INV_X1    g131(.A(G125), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n316), .B1(new_n320), .B2(new_n314), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n321), .A2(new_n210), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n317), .A2(new_n319), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n210), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n204), .A2(G119), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT23), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n204), .A2(KEYINPUT23), .A3(G119), .ZN(new_n329));
  INV_X1    g143(.A(G110), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n255), .A2(G128), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n328), .A2(new_n329), .A3(new_n330), .A4(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n326), .A2(new_n331), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT24), .B(G110), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n332), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n333), .B1(new_n332), .B2(new_n336), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n323), .B(new_n325), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  OR3_X1    g153(.A1(new_n334), .A2(new_n335), .A3(KEYINPUT73), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT73), .B1(new_n334), .B2(new_n335), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n328), .A2(new_n329), .A3(new_n331), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G110), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n321), .A2(new_n210), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n342), .B(new_n344), .C1(new_n346), .C2(new_n322), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n339), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT22), .B(G137), .ZN(new_n349));
  INV_X1    g163(.A(G953), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(G221), .A3(G234), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n349), .B(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT75), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n348), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n339), .A2(new_n347), .A3(KEYINPUT75), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n352), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n354), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n313), .B1(new_n360), .B2(G902), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n339), .A2(new_n347), .A3(KEYINPUT75), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT75), .B1(new_n339), .B2(new_n347), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n359), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n353), .ZN(new_n365));
  INV_X1    g179(.A(G902), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(KEYINPUT25), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n361), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G234), .ZN(new_n369));
  OAI21_X1  g183(.A(G217), .B1(new_n369), .B2(G902), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n370), .B(KEYINPUT72), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n366), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n373), .B(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  AOI22_X1  g190(.A1(new_n368), .A2(new_n372), .B1(new_n376), .B2(new_n365), .ZN(new_n377));
  OAI21_X1  g191(.A(G214), .B1(G237), .B2(G902), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n226), .A2(new_n228), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n379), .A2(G125), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n318), .B1(new_n212), .B2(new_n217), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n350), .A2(G224), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n383), .B(KEYINPUT84), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n382), .B(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(KEYINPUT80), .B(G101), .ZN(new_n386));
  INV_X1    g200(.A(G104), .ZN(new_n387));
  OAI21_X1  g201(.A(KEYINPUT3), .B1(new_n387), .B2(G107), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT3), .ZN(new_n389));
  INV_X1    g203(.A(G107), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(G104), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n387), .A2(G107), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n386), .A2(new_n388), .A3(new_n391), .A4(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n388), .A2(new_n391), .A3(new_n392), .ZN(new_n394));
  AOI22_X1  g208(.A1(new_n393), .A2(KEYINPUT4), .B1(G101), .B2(new_n394), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n394), .A2(KEYINPUT4), .A3(G101), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n265), .B(new_n263), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G101), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n390), .A2(G104), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n398), .B1(new_n399), .B2(new_n392), .ZN(new_n400));
  INV_X1    g214(.A(new_n394), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n400), .B1(new_n401), .B2(new_n386), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT5), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n259), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(G113), .B1(new_n256), .B2(KEYINPUT5), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n402), .B(new_n262), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n397), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT83), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT6), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n397), .A2(new_n406), .A3(KEYINPUT83), .ZN(new_n411));
  XNOR2_X1  g225(.A(G110), .B(G122), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n409), .A2(new_n410), .A3(new_n411), .A4(new_n413), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n397), .A2(new_n406), .A3(KEYINPUT83), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT83), .B1(new_n397), .B2(new_n406), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n415), .A2(new_n416), .A3(new_n412), .ZN(new_n417));
  OAI21_X1  g231(.A(KEYINPUT6), .B1(new_n407), .B2(new_n413), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n385), .B(new_n414), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n407), .A2(new_n413), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n387), .A2(G107), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n390), .A2(G104), .ZN(new_n422));
  OAI21_X1  g236(.A(G101), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  XOR2_X1   g237(.A(KEYINPUT80), .B(G101), .Z(new_n424));
  OAI21_X1  g238(.A(new_n423), .B1(new_n394), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n404), .A2(KEYINPUT85), .ZN(new_n426));
  INV_X1    g240(.A(new_n405), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT85), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n428), .B1(new_n259), .B2(new_n403), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n425), .B1(new_n430), .B2(new_n262), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n412), .B(KEYINPUT8), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n262), .B1(new_n404), .B2(new_n405), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n432), .B1(new_n402), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n383), .A2(KEYINPUT7), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  OAI22_X1  g250(.A1(new_n431), .A2(new_n434), .B1(new_n382), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n420), .A2(new_n437), .ZN(new_n438));
  NOR3_X1   g252(.A1(new_n380), .A2(new_n381), .A3(new_n435), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(KEYINPUT86), .ZN(new_n440));
  AOI21_X1  g254(.A(G902), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G210), .B1(G237), .B2(G902), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n419), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n442), .B1(new_n419), .B2(new_n441), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n443), .B1(new_n444), .B2(KEYINPUT87), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT87), .ZN(new_n446));
  AOI211_X1 g260(.A(new_n446), .B(new_n442), .C1(new_n419), .C2(new_n441), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n378), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT20), .ZN(new_n449));
  XNOR2_X1  g263(.A(G113), .B(G122), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(new_n387), .ZN(new_n451));
  INV_X1    g265(.A(G237), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n452), .A2(new_n350), .A3(G143), .A4(G214), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT89), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT89), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n270), .A2(new_n455), .A3(G143), .A4(G214), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G214), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n458), .A2(G237), .A3(G953), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT88), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n459), .A2(new_n460), .A3(G143), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n270), .A2(G214), .ZN(new_n462));
  AOI21_X1  g276(.A(KEYINPUT88), .B1(new_n462), .B2(new_n208), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n457), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(KEYINPUT18), .A2(G131), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n464), .B(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n320), .A2(G146), .ZN(new_n467));
  XOR2_X1   g281(.A(new_n467), .B(KEYINPUT91), .Z(new_n468));
  AND2_X1   g282(.A1(new_n325), .A2(KEYINPUT90), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n468), .A2(new_n469), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n466), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n460), .B1(new_n459), .B2(G143), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n462), .A2(KEYINPUT88), .A3(new_n208), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n473), .A2(new_n474), .B1(new_n454), .B2(new_n456), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT92), .B1(new_n475), .B2(new_n235), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT92), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n464), .A2(new_n477), .A3(G131), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT95), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n480), .B1(new_n346), .B2(new_n322), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n323), .A2(KEYINPUT95), .A3(new_n345), .ZN(new_n482));
  AOI22_X1  g296(.A1(new_n479), .A2(KEYINPUT17), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT17), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n475), .A2(new_n235), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n476), .A2(new_n478), .A3(new_n484), .A4(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT96), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n486), .A2(new_n487), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n451), .B(new_n472), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n479), .B1(new_n235), .B2(new_n475), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT93), .ZN(new_n493));
  XOR2_X1   g307(.A(new_n493), .B(KEYINPUT19), .Z(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n210), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT94), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT94), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n494), .A2(new_n497), .A3(new_n210), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n496), .A2(new_n323), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n472), .B1(new_n492), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n451), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n491), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(G475), .A2(G902), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n449), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n504), .ZN(new_n506));
  AOI211_X1 g320(.A(KEYINPUT20), .B(new_n506), .C1(new_n491), .C2(new_n502), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n472), .B1(new_n489), .B2(new_n490), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n501), .ZN(new_n509));
  AOI21_X1  g323(.A(G902), .B1(new_n509), .B2(new_n491), .ZN(new_n510));
  INV_X1    g324(.A(G475), .ZN(new_n511));
  OAI22_X1  g325(.A1(new_n505), .A2(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(G116), .B(G122), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT14), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n257), .A2(KEYINPUT14), .A3(G122), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(G107), .A3(new_n516), .ZN(new_n517));
  XOR2_X1   g331(.A(new_n517), .B(KEYINPUT97), .Z(new_n518));
  NAND2_X1  g332(.A1(new_n513), .A2(new_n390), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n208), .A2(G128), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n204), .A2(G143), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(new_n243), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n518), .A2(new_n519), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n513), .B(new_n390), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT13), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n521), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n520), .A2(new_n526), .ZN(new_n529));
  OAI21_X1  g343(.A(G134), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n525), .B(new_n530), .C1(new_n243), .C2(new_n522), .ZN(new_n531));
  XOR2_X1   g345(.A(KEYINPUT9), .B(G234), .Z(new_n532));
  XNOR2_X1  g346(.A(new_n532), .B(KEYINPUT78), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(G217), .A3(new_n350), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n524), .A2(new_n531), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n536), .B1(new_n524), .B2(new_n531), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n366), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT15), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n541), .A3(G478), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(G478), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n366), .B(new_n543), .C1(new_n538), .C2(new_n539), .ZN(new_n544));
  AND2_X1   g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(G952), .ZN(new_n546));
  AOI211_X1 g360(.A(G953), .B(new_n546), .C1(G234), .C2(G237), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT21), .B(G898), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  OAI211_X1 g364(.A(G902), .B(G953), .C1(new_n369), .C2(new_n452), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n545), .A2(new_n552), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n448), .A2(new_n512), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT82), .B(G469), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n219), .B1(new_n395), .B2(new_n396), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT10), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n559));
  OAI21_X1  g373(.A(G128), .B1(new_n209), .B2(new_n224), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n561), .A2(new_n228), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n558), .B1(new_n562), .B2(new_n425), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n402), .A2(KEYINPUT10), .A3(new_n379), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n557), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n202), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n247), .A2(new_n557), .A3(new_n563), .A4(new_n564), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(G110), .B(G140), .ZN(new_n569));
  INV_X1    g383(.A(G227), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(G953), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n569), .B(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n572), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n567), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n425), .A2(new_n226), .A3(new_n228), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n576), .B1(new_n562), .B2(new_n425), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n202), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT12), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n202), .A2(new_n577), .A3(KEYINPUT12), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n575), .A2(new_n582), .ZN(new_n583));
  AOI211_X1 g397(.A(G902), .B(new_n556), .C1(new_n573), .C2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT81), .B1(new_n582), .B2(new_n567), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n202), .A2(new_n577), .A3(KEYINPUT12), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT12), .B1(new_n202), .B2(new_n577), .ZN(new_n587));
  OAI211_X1 g401(.A(KEYINPUT81), .B(new_n567), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n572), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n575), .A2(new_n566), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n366), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n584), .B1(new_n593), .B2(G469), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n534), .A2(new_n366), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(G221), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT79), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n312), .A2(new_n377), .A3(new_n554), .A4(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n424), .B(KEYINPUT98), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(G3));
  AOI21_X1  g415(.A(new_n297), .B1(new_n287), .B2(new_n366), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n603), .A2(new_n291), .A3(new_n293), .ZN(new_n604));
  INV_X1    g418(.A(new_n584), .ZN(new_n605));
  AOI21_X1  g419(.A(G902), .B1(new_n590), .B2(new_n591), .ZN(new_n606));
  INV_X1    g420(.A(G469), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n597), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n377), .A3(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n419), .A2(new_n441), .A3(new_n442), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n378), .B1(new_n612), .B2(new_n444), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(KEYINPUT99), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT99), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n615), .B(new_n378), .C1(new_n612), .C2(new_n444), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n552), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(KEYINPUT33), .B1(new_n538), .B2(new_n539), .ZN(new_n618));
  INV_X1    g432(.A(new_n539), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n619), .A2(new_n620), .A3(new_n537), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n618), .A2(new_n621), .A3(G478), .ZN(new_n622));
  NAND2_X1  g436(.A1(G478), .A2(G902), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n622), .B(new_n623), .C1(G478), .C2(new_n540), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n512), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n617), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n611), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT34), .B(G104), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  NAND2_X1  g444(.A1(new_n503), .A2(new_n504), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(KEYINPUT20), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n503), .A2(new_n449), .A3(new_n504), .ZN(new_n633));
  INV_X1    g447(.A(new_n490), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n634), .A2(new_n488), .A3(new_n483), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n451), .B1(new_n635), .B2(new_n472), .ZN(new_n636));
  INV_X1    g450(.A(new_n491), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n366), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  AOI22_X1  g452(.A1(new_n632), .A2(new_n633), .B1(new_n638), .B2(G475), .ZN(new_n639));
  INV_X1    g453(.A(new_n545), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n617), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n611), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(new_n390), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT100), .B(KEYINPUT35), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  AOI21_X1  g460(.A(KEYINPUT25), .B1(new_n365), .B2(new_n366), .ZN(new_n647));
  AOI211_X1 g461(.A(new_n313), .B(G902), .C1(new_n364), .C2(new_n353), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n372), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n359), .A2(KEYINPUT36), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n358), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n358), .A2(new_n650), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n649), .B1(new_n654), .B2(new_n375), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(new_n608), .A3(new_n609), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n287), .A2(KEYINPUT71), .A3(new_n288), .ZN(new_n658));
  AOI21_X1  g472(.A(KEYINPUT71), .B1(new_n287), .B2(new_n288), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n658), .A2(new_n659), .A3(new_n602), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n554), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT37), .B(G110), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  NAND2_X1  g477(.A1(new_n614), .A2(new_n616), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n656), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT101), .B(G900), .Z(new_n666));
  OAI21_X1  g480(.A(new_n548), .B1(new_n666), .B2(new_n551), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n639), .A2(new_n640), .A3(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n665), .A2(new_n669), .A3(new_n312), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G128), .ZN(G30));
  NOR2_X1   g485(.A1(new_n639), .A2(new_n545), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n667), .B(KEYINPUT39), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n598), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT40), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n378), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n676), .A2(new_n677), .A3(new_n655), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n366), .B1(new_n306), .B2(new_n274), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n282), .B1(new_n284), .B2(new_n269), .ZN(new_n680));
  OAI21_X1  g494(.A(G472), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT102), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OAI211_X1 g497(.A(KEYINPUT102), .B(G472), .C1(new_n679), .C2(new_n680), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n295), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n294), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n445), .A2(new_n447), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT38), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n674), .B2(new_n675), .ZN(new_n689));
  AND4_X1   g503(.A1(new_n672), .A2(new_n678), .A3(new_n686), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(new_n208), .ZN(G45));
  NAND3_X1  g505(.A1(new_n512), .A2(new_n625), .A3(new_n667), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n665), .A2(new_n312), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  INV_X1    g509(.A(new_n377), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n696), .B1(new_n294), .B2(new_n311), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n573), .A2(new_n583), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n607), .B1(new_n698), .B2(new_n366), .ZN(new_n699));
  INV_X1    g513(.A(new_n596), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n699), .A2(new_n584), .A3(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n697), .A2(new_n627), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT41), .B(G113), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G15));
  NAND3_X1  g518(.A1(new_n697), .A2(new_n642), .A3(new_n701), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT103), .B(G116), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G18));
  NAND3_X1  g521(.A1(new_n614), .A2(new_n616), .A3(new_n701), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  AOI22_X1  g523(.A1(new_n368), .A2(new_n372), .B1(new_n376), .B2(new_n653), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n512), .A2(new_n553), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n312), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  AND3_X1   g527(.A1(new_n614), .A2(new_n552), .A3(new_n616), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n276), .B(new_n286), .C1(new_n307), .C2(new_n274), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n715), .A2(KEYINPUT104), .A3(new_n288), .ZN(new_n716));
  AOI21_X1  g530(.A(KEYINPUT104), .B1(new_n715), .B2(new_n288), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n716), .A2(new_n717), .A3(new_n602), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n512), .A2(new_n701), .A3(new_n640), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n714), .A2(new_n718), .A3(new_n377), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G122), .ZN(G24));
  NOR2_X1   g535(.A1(new_n708), .A2(new_n692), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n715), .A2(new_n288), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT104), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n715), .A2(KEYINPUT104), .A3(new_n288), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n725), .A2(new_n603), .A3(new_n655), .A4(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n722), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT105), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT105), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n722), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  NAND4_X1  g548(.A1(new_n687), .A2(new_n378), .A3(new_n608), .A4(new_n596), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n692), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT42), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n697), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n632), .A2(new_n633), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n638), .A2(G475), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n624), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n567), .B1(new_n586), .B2(new_n587), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT81), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n588), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n745), .A2(new_n572), .B1(new_n575), .B2(new_n566), .ZN(new_n746));
  OAI21_X1  g560(.A(G469), .B1(new_n746), .B2(G902), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n700), .B1(new_n747), .B2(new_n605), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n445), .A2(new_n677), .A3(new_n447), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n741), .A2(new_n748), .A3(new_n667), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n289), .A2(new_n292), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n306), .A2(KEYINPUT28), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n279), .A3(new_n308), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n366), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT29), .B1(new_n298), .B2(new_n299), .ZN(new_n755));
  OAI21_X1  g569(.A(G472), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n751), .A2(new_n756), .A3(new_n295), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n377), .ZN(new_n758));
  OAI21_X1  g572(.A(KEYINPUT42), .B1(new_n750), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n738), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(new_n235), .ZN(G33));
  INV_X1    g575(.A(KEYINPUT106), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n658), .A2(new_n659), .A3(KEYINPUT32), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n756), .A2(new_n295), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n377), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n512), .A2(new_n545), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n766), .A2(new_n748), .A3(new_n667), .A4(new_n749), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n762), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n735), .A2(new_n668), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n697), .A2(new_n769), .A3(KEYINPUT106), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G134), .ZN(G36));
  NAND2_X1  g586(.A1(new_n639), .A2(new_n625), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT43), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n604), .A3(new_n655), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT44), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT107), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n778), .B(new_n779), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n776), .A2(new_n777), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n746), .A2(KEYINPUT45), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n746), .A2(KEYINPUT45), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(G469), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(G469), .A2(G902), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT46), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n584), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n784), .A2(KEYINPUT46), .A3(new_n785), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n789), .A2(new_n596), .A3(new_n673), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n780), .A2(new_n749), .A3(new_n781), .A4(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G137), .ZN(G39));
  OR3_X1    g606(.A1(new_n445), .A2(new_n677), .A3(new_n447), .ZN(new_n793));
  NOR4_X1   g607(.A1(new_n312), .A2(new_n377), .A3(new_n692), .A4(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT47), .B1(new_n789), .B2(new_n596), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT47), .ZN(new_n796));
  AOI211_X1 g610(.A(new_n796), .B(new_n700), .C1(new_n787), .C2(new_n788), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n794), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n798), .B(KEYINPUT108), .Z(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(new_n315), .ZN(G42));
  NAND2_X1  g614(.A1(new_n718), .A2(new_n377), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n775), .A2(new_n547), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n775), .A2(KEYINPUT114), .A3(new_n547), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n801), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n688), .A2(new_n677), .A3(new_n701), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(KEYINPUT50), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n801), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n775), .A2(KEYINPUT114), .A3(new_n547), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT114), .B1(new_n775), .B2(new_n547), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n809), .B(new_n807), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT50), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n808), .A2(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n749), .A2(new_n701), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n728), .B(new_n816), .C1(new_n810), .C2(new_n811), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT115), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n804), .A2(new_n805), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n819), .A2(new_n820), .A3(new_n728), .A4(new_n816), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n686), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n823), .A2(new_n377), .A3(new_n547), .A4(new_n816), .ZN(new_n824));
  OR3_X1    g638(.A1(new_n824), .A2(new_n512), .A3(new_n625), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n815), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n826), .A2(KEYINPUT116), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n809), .B(new_n749), .C1(new_n810), .C2(new_n811), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n795), .A2(new_n797), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n699), .A2(new_n584), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n597), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n826), .A2(KEYINPUT116), .B1(new_n829), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n827), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n815), .A2(new_n822), .A3(new_n825), .ZN(new_n838));
  INV_X1    g652(.A(new_n795), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n789), .A2(KEYINPUT47), .A3(new_n596), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n839), .A2(new_n840), .A3(new_n841), .A4(new_n832), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n842), .A2(new_n829), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n841), .B1(new_n830), .B2(new_n832), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n836), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n838), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n758), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n849), .B(new_n816), .C1(new_n810), .C2(new_n811), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT48), .ZN(new_n851));
  OR3_X1    g665(.A1(new_n850), .A2(KEYINPUT119), .A3(new_n851), .ZN(new_n852));
  XNOR2_X1  g666(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  OAI211_X1 g668(.A(G952), .B(new_n350), .C1(new_n824), .C2(new_n626), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(new_n806), .B2(new_n709), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n852), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(KEYINPUT120), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT120), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n852), .A2(new_n856), .A3(new_n859), .A4(new_n854), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n842), .A2(new_n829), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT51), .B1(new_n862), .B2(new_n844), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT118), .B1(new_n826), .B2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n837), .A2(new_n848), .A3(new_n861), .A4(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT110), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n626), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n512), .A2(new_n625), .A3(KEYINPUT110), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n868), .A2(new_n641), .A3(new_n869), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n378), .B(new_n552), .C1(new_n445), .C2(new_n447), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n870), .A2(new_n611), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n873), .A2(new_n702), .A3(new_n705), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n599), .A2(new_n712), .A3(new_n720), .A4(new_n661), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n874), .A2(new_n875), .A3(new_n760), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n542), .A2(new_n544), .A3(new_n667), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n739), .A2(new_n740), .A3(new_n877), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n656), .A2(new_n793), .A3(new_n878), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n879), .A2(new_n312), .B1(new_n736), .B2(new_n728), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n765), .A2(new_n767), .A3(new_n762), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT106), .B1(new_n697), .B2(new_n769), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT111), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n771), .A2(KEYINPUT111), .A3(new_n880), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n876), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n731), .B1(new_n722), .B2(new_n728), .ZN(new_n888));
  NOR4_X1   g702(.A1(new_n727), .A2(new_n708), .A3(new_n692), .A4(KEYINPUT105), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n670), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n664), .ZN(new_n891));
  AND4_X1   g705(.A1(new_n608), .A2(new_n710), .A3(new_n596), .A4(new_n667), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n686), .A2(new_n891), .A3(new_n892), .A4(new_n672), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n694), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT52), .B1(new_n890), .B2(new_n894), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n694), .A2(new_n893), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT52), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n733), .A2(new_n896), .A3(new_n897), .A4(new_n670), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n866), .B1(new_n887), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT113), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI211_X1 g716(.A(KEYINPUT113), .B(new_n866), .C1(new_n887), .C2(new_n899), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n665), .A2(new_n669), .A3(new_n312), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n730), .B2(new_n732), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n897), .B1(new_n905), .B2(new_n896), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n890), .A2(KEYINPUT52), .A3(new_n894), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT112), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT112), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n895), .A2(new_n898), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n887), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  AOI22_X1  g725(.A1(new_n902), .A2(new_n903), .B1(new_n911), .B2(KEYINPUT53), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT54), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OR2_X1    g728(.A1(new_n911), .A2(KEYINPUT53), .ZN(new_n915));
  OR3_X1    g729(.A1(new_n887), .A2(new_n899), .A3(new_n866), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n914), .B1(new_n917), .B2(new_n913), .ZN(new_n918));
  OAI22_X1  g732(.A1(new_n865), .A2(new_n918), .B1(G952), .B2(G953), .ZN(new_n919));
  INV_X1    g733(.A(new_n831), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n920), .A2(KEYINPUT49), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT109), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(KEYINPUT49), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n923), .A2(new_n377), .A3(new_n378), .A4(new_n609), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n922), .A2(new_n773), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n925), .A2(new_n823), .A3(new_n688), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n919), .A2(new_n926), .ZN(G75));
  OAI21_X1  g741(.A(new_n414), .B1(new_n417), .B2(new_n418), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT121), .Z(new_n929));
  XNOR2_X1  g743(.A(new_n385), .B(KEYINPUT55), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n929), .B(new_n930), .Z(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n912), .A2(new_n366), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(G210), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT122), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n935), .A2(KEYINPUT56), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n932), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n936), .ZN(new_n938));
  AOI211_X1 g752(.A(new_n931), .B(new_n938), .C1(new_n933), .C2(G210), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n350), .A2(G952), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(G51));
  XOR2_X1   g755(.A(new_n785), .B(KEYINPUT57), .Z(new_n942));
  INV_X1    g756(.A(new_n914), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n912), .A2(new_n913), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n698), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n902), .A2(new_n903), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n911), .A2(KEYINPUT53), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(G902), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n950), .A2(new_n784), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n940), .B1(new_n946), .B2(new_n951), .ZN(G54));
  INV_X1    g766(.A(new_n940), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n933), .A2(KEYINPUT58), .A3(G475), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n953), .B1(new_n954), .B2(new_n503), .ZN(new_n955));
  AND4_X1   g769(.A1(KEYINPUT58), .A2(new_n933), .A3(G475), .A4(new_n503), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n955), .A2(new_n956), .ZN(G60));
  NOR2_X1   g771(.A1(new_n943), .A2(new_n944), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n618), .A2(new_n621), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT123), .Z(new_n960));
  XNOR2_X1  g774(.A(new_n623), .B(KEYINPUT59), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n953), .B1(new_n958), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n960), .B1(new_n918), .B2(new_n961), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n963), .A2(new_n964), .ZN(G63));
  INV_X1    g779(.A(KEYINPUT61), .ZN(new_n966));
  NAND2_X1  g780(.A1(G217), .A2(G902), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT60), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n947), .B2(new_n948), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n966), .B1(new_n969), .B2(new_n653), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n970), .B(new_n953), .C1(new_n365), .C2(new_n969), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n953), .B1(new_n969), .B2(new_n365), .ZN(new_n972));
  AOI21_X1  g786(.A(KEYINPUT125), .B1(new_n969), .B2(new_n653), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT125), .ZN(new_n974));
  NOR4_X1   g788(.A1(new_n912), .A2(new_n974), .A3(new_n654), .A4(new_n968), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n972), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  XNOR2_X1  g790(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n971), .B1(new_n976), .B2(new_n977), .ZN(G66));
  AND2_X1   g792(.A1(new_n550), .A2(G224), .ZN(new_n979));
  OAI21_X1  g793(.A(KEYINPUT126), .B1(new_n979), .B2(new_n350), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n874), .A2(new_n875), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n981), .A2(G953), .ZN(new_n982));
  MUX2_X1   g796(.A(new_n980), .B(KEYINPUT126), .S(new_n982), .Z(new_n983));
  OAI21_X1  g797(.A(new_n929), .B1(G898), .B2(new_n350), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n983), .B(new_n984), .ZN(G69));
  NAND2_X1  g799(.A1(new_n234), .A2(new_n250), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(new_n494), .ZN(new_n987));
  NAND3_X1  g801(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n870), .A2(new_n674), .A3(new_n697), .A4(new_n749), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n791), .A2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n799), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n905), .A2(new_n694), .ZN(new_n992));
  OR3_X1    g806(.A1(new_n690), .A2(KEYINPUT62), .A3(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(KEYINPUT62), .B1(new_n690), .B2(new_n992), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n990), .A2(new_n991), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n987), .B(new_n988), .C1(new_n995), .C2(G953), .ZN(new_n996));
  INV_X1    g810(.A(new_n992), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n790), .A2(new_n891), .A3(new_n672), .A4(new_n849), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n760), .B1(new_n768), .B2(new_n770), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n791), .A2(new_n997), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT127), .ZN(new_n1001));
  OR3_X1    g815(.A1(new_n1000), .A2(new_n1001), .A3(new_n799), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1001), .B1(new_n1000), .B2(new_n799), .ZN(new_n1003));
  AOI21_X1  g817(.A(G953), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n570), .A2(G900), .A3(G953), .ZN(new_n1005));
  OR2_X1    g819(.A1(new_n987), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n996), .B1(new_n1004), .B2(new_n1006), .ZN(G72));
  NAND2_X1  g821(.A1(G472), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT63), .Z(new_n1009));
  INV_X1    g823(.A(new_n981), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1009), .B1(new_n995), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(new_n680), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n953), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1002), .A2(new_n1003), .A3(new_n981), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n299), .B1(new_n1014), .B2(new_n1009), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n299), .A2(new_n1009), .ZN(new_n1016));
  NOR3_X1   g830(.A1(new_n917), .A2(new_n680), .A3(new_n1016), .ZN(new_n1017));
  NOR3_X1   g831(.A1(new_n1013), .A2(new_n1015), .A3(new_n1017), .ZN(G57));
endmodule


