

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730;

  INV_X1 U375 ( .A(G953), .ZN(n714) );
  XNOR2_X2 U376 ( .A(n510), .B(KEYINPUT40), .ZN(n729) );
  AND2_X2 U377 ( .A1(n551), .A2(n624), .ZN(n510) );
  AND2_X2 U378 ( .A1(n415), .A2(n417), .ZN(n414) );
  NAND2_X2 U379 ( .A1(n360), .A2(n656), .ZN(n616) );
  OR2_X2 U380 ( .A1(n602), .A2(G902), .ZN(n419) );
  XNOR2_X2 U381 ( .A(n433), .B(n432), .ZN(n528) );
  XNOR2_X2 U382 ( .A(n500), .B(G469), .ZN(n389) );
  NOR2_X1 U383 ( .A1(n574), .A2(n559), .ZN(n561) );
  INV_X1 U384 ( .A(n585), .ZN(n582) );
  XNOR2_X1 U385 ( .A(KEYINPUT3), .B(G119), .ZN(n384) );
  AND2_X1 U386 ( .A1(n368), .A2(n365), .ZN(n376) );
  AND2_X1 U387 ( .A1(n366), .A2(n365), .ZN(n375) );
  XNOR2_X1 U388 ( .A(n561), .B(n560), .ZN(n565) );
  XNOR2_X1 U389 ( .A(n386), .B(n385), .ZN(n647) );
  INV_X1 U390 ( .A(n515), .ZN(n624) );
  NOR2_X1 U391 ( .A1(n680), .A2(n453), .ZN(n456) );
  OR2_X1 U392 ( .A1(n684), .A2(G902), .ZN(n500) );
  XNOR2_X1 U393 ( .A(n374), .B(n373), .ZN(n680) );
  XNOR2_X1 U394 ( .A(n462), .B(n407), .ZN(n373) );
  XNOR2_X1 U395 ( .A(n705), .B(n498), .ZN(n374) );
  XNOR2_X1 U396 ( .A(n410), .B(n408), .ZN(n407) );
  XNOR2_X1 U397 ( .A(n454), .B(KEYINPUT78), .ZN(n455) );
  XNOR2_X1 U398 ( .A(n704), .B(KEYINPUT69), .ZN(n498) );
  XNOR2_X1 U399 ( .A(n463), .B(G125), .ZN(n450) );
  XNOR2_X1 U400 ( .A(G110), .B(n447), .ZN(n704) );
  XNOR2_X1 U401 ( .A(n384), .B(G101), .ZN(n411) );
  INV_X1 U402 ( .A(G146), .ZN(n463) );
  NOR2_X2 U403 ( .A1(n556), .A2(n524), .ZN(n622) );
  XNOR2_X1 U404 ( .A(n530), .B(n387), .ZN(n642) );
  INV_X1 U405 ( .A(KEYINPUT38), .ZN(n387) );
  XNOR2_X1 U406 ( .A(KEYINPUT22), .B(KEYINPUT71), .ZN(n560) );
  INV_X1 U407 ( .A(KEYINPUT45), .ZN(n594) );
  NOR2_X1 U408 ( .A1(n728), .A2(n403), .ZN(n402) );
  XNOR2_X1 U409 ( .A(n450), .B(n395), .ZN(n479) );
  INV_X1 U410 ( .A(KEYINPUT10), .ZN(n395) );
  XOR2_X1 U411 ( .A(G140), .B(G122), .Z(n423) );
  XNOR2_X1 U412 ( .A(G143), .B(G131), .ZN(n422) );
  XNOR2_X1 U413 ( .A(KEYINPUT11), .B(KEYINPUT100), .ZN(n425) );
  XOR2_X1 U414 ( .A(KEYINPUT12), .B(KEYINPUT99), .Z(n426) );
  XNOR2_X1 U415 ( .A(n430), .B(KEYINPUT98), .ZN(n400) );
  XNOR2_X1 U416 ( .A(KEYINPUT87), .B(KEYINPUT48), .ZN(n542) );
  XNOR2_X1 U417 ( .A(n469), .B(n352), .ZN(n420) );
  XNOR2_X1 U418 ( .A(n482), .B(n481), .ZN(n483) );
  INV_X1 U419 ( .A(KEYINPUT24), .ZN(n481) );
  XOR2_X1 U420 ( .A(G128), .B(KEYINPUT23), .Z(n482) );
  XNOR2_X1 U421 ( .A(G119), .B(G110), .ZN(n485) );
  XNOR2_X1 U422 ( .A(n712), .B(n463), .ZN(n497) );
  XOR2_X1 U423 ( .A(G137), .B(G140), .Z(n496) );
  XNOR2_X1 U424 ( .A(n459), .B(n458), .ZN(n674) );
  INV_X1 U425 ( .A(KEYINPUT41), .ZN(n458) );
  NAND2_X1 U426 ( .A1(n361), .A2(n557), .ZN(n459) );
  INV_X1 U427 ( .A(n647), .ZN(n361) );
  XNOR2_X1 U428 ( .A(n380), .B(n379), .ZN(n551) );
  INV_X1 U429 ( .A(KEYINPUT39), .ZN(n379) );
  NOR2_X1 U430 ( .A1(n506), .A2(n377), .ZN(n380) );
  XNOR2_X1 U431 ( .A(n493), .B(n492), .ZN(n566) );
  NOR2_X1 U432 ( .A1(n696), .A2(G902), .ZN(n493) );
  NAND2_X1 U433 ( .A1(n413), .A2(n416), .ZN(n412) );
  BUF_X1 U434 ( .A(n690), .Z(n694) );
  XNOR2_X1 U435 ( .A(n497), .B(n391), .ZN(n684) );
  XNOR2_X1 U436 ( .A(n498), .B(n392), .ZN(n391) );
  XNOR2_X1 U437 ( .A(n393), .B(n496), .ZN(n392) );
  XNOR2_X1 U438 ( .A(n499), .B(n394), .ZN(n393) );
  NOR2_X1 U439 ( .A1(n639), .A2(n638), .ZN(n641) );
  INV_X1 U440 ( .A(KEYINPUT84), .ZN(n640) );
  NOR2_X1 U441 ( .A1(G237), .A2(G953), .ZN(n424) );
  XNOR2_X1 U442 ( .A(n471), .B(KEYINPUT20), .ZN(n487) );
  XNOR2_X1 U443 ( .A(n383), .B(n381), .ZN(n655) );
  XNOR2_X1 U444 ( .A(n382), .B(KEYINPUT21), .ZN(n381) );
  NAND2_X1 U445 ( .A1(n487), .A2(G221), .ZN(n383) );
  INV_X1 U446 ( .A(KEYINPUT93), .ZN(n382) );
  XNOR2_X1 U447 ( .A(n462), .B(n461), .ZN(n712) );
  XOR2_X1 U448 ( .A(KEYINPUT67), .B(G134), .Z(n460) );
  AND2_X1 U449 ( .A1(n713), .A2(n453), .ZN(n367) );
  INV_X1 U450 ( .A(KEYINPUT111), .ZN(n385) );
  NAND2_X1 U451 ( .A1(n642), .A2(n643), .ZN(n386) );
  AND2_X1 U452 ( .A1(n642), .A2(n508), .ZN(n390) );
  OR2_X1 U453 ( .A1(G237), .A2(G902), .ZN(n457) );
  XNOR2_X1 U454 ( .A(G116), .B(G134), .ZN(n435) );
  XOR2_X1 U455 ( .A(G107), .B(G122), .Z(n436) );
  XOR2_X1 U456 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n438) );
  XNOR2_X1 U457 ( .A(n401), .B(n399), .ZN(n686) );
  XNOR2_X1 U458 ( .A(n400), .B(n431), .ZN(n399) );
  XNOR2_X1 U459 ( .A(n428), .B(n429), .ZN(n401) );
  XOR2_X1 U460 ( .A(KEYINPUT91), .B(KEYINPUT17), .Z(n451) );
  XNOR2_X1 U461 ( .A(n452), .B(n409), .ZN(n408) );
  INV_X1 U462 ( .A(KEYINPUT18), .ZN(n409) );
  XNOR2_X1 U463 ( .A(G122), .B(KEYINPUT16), .ZN(n449) );
  NOR2_X1 U464 ( .A1(KEYINPUT2), .A2(n713), .ZN(n633) );
  NOR2_X1 U465 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U466 ( .A1(n544), .A2(n547), .ZN(n398) );
  XNOR2_X1 U467 ( .A(n358), .B(n504), .ZN(n505) );
  XNOR2_X1 U468 ( .A(KEYINPUT30), .B(KEYINPUT110), .ZN(n504) );
  NAND2_X1 U469 ( .A1(n582), .A2(n643), .ZN(n358) );
  XNOR2_X1 U470 ( .A(n362), .B(KEYINPUT95), .ZN(n586) );
  INV_X1 U471 ( .A(n566), .ZN(n656) );
  XNOR2_X1 U472 ( .A(n604), .B(n603), .ZN(n605) );
  XNOR2_X1 U473 ( .A(n484), .B(n364), .ZN(n486) );
  XNOR2_X1 U474 ( .A(n483), .B(n485), .ZN(n364) );
  XNOR2_X1 U475 ( .A(KEYINPUT112), .B(n517), .ZN(n723) );
  NAND2_X1 U476 ( .A1(n396), .A2(n652), .ZN(n517) );
  XNOR2_X1 U477 ( .A(n398), .B(n397), .ZN(n396) );
  XNOR2_X1 U478 ( .A(KEYINPUT36), .B(KEYINPUT88), .ZN(n397) );
  XNOR2_X1 U479 ( .A(n405), .B(KEYINPUT35), .ZN(n728) );
  XNOR2_X1 U480 ( .A(n569), .B(n404), .ZN(n726) );
  XNOR2_X1 U481 ( .A(KEYINPUT64), .B(KEYINPUT32), .ZN(n404) );
  XNOR2_X1 U482 ( .A(n682), .B(n369), .ZN(n685) );
  XNOR2_X1 U483 ( .A(n684), .B(n683), .ZN(n369) );
  AND2_X1 U484 ( .A1(n673), .A2(n370), .ZN(n676) );
  AND2_X1 U485 ( .A1(n672), .A2(n354), .ZN(n370) );
  XOR2_X1 U486 ( .A(n465), .B(n464), .Z(n352) );
  OR2_X1 U487 ( .A1(n536), .A2(n537), .ZN(n353) );
  INV_X1 U488 ( .A(G101), .ZN(n394) );
  OR2_X1 U489 ( .A1(n675), .A2(n674), .ZN(n354) );
  XOR2_X1 U490 ( .A(n688), .B(n687), .Z(n355) );
  XNOR2_X1 U491 ( .A(G902), .B(KEYINPUT15), .ZN(n596) );
  OR2_X1 U492 ( .A1(n635), .A2(n421), .ZN(n356) );
  XOR2_X1 U493 ( .A(n680), .B(n679), .Z(n357) );
  NOR2_X1 U494 ( .A1(G952), .A2(n714), .ZN(n698) );
  INV_X1 U495 ( .A(n698), .ZN(n365) );
  NAND2_X1 U496 ( .A1(n378), .A2(n390), .ZN(n377) );
  NOR2_X1 U497 ( .A1(n729), .A2(n730), .ZN(n511) );
  AND2_X2 U498 ( .A1(n371), .A2(n372), .ZN(n690) );
  XNOR2_X1 U499 ( .A(n359), .B(KEYINPUT44), .ZN(n593) );
  XNOR2_X1 U500 ( .A(n564), .B(KEYINPUT65), .ZN(n360) );
  NAND2_X1 U501 ( .A1(n616), .A2(n402), .ZN(n359) );
  NAND2_X1 U502 ( .A1(n690), .A2(G472), .ZN(n606) );
  INV_X1 U503 ( .A(n372), .ZN(n638) );
  NAND2_X1 U504 ( .A1(n651), .A2(n389), .ZN(n362) );
  NAND2_X1 U505 ( .A1(n363), .A2(n356), .ZN(n371) );
  NAND2_X1 U506 ( .A1(n367), .A2(n699), .ZN(n363) );
  NOR2_X1 U507 ( .A1(n353), .A2(n538), .ZN(n539) );
  INV_X1 U508 ( .A(n505), .ZN(n378) );
  NAND2_X1 U509 ( .A1(n601), .A2(n699), .ZN(n372) );
  XNOR2_X1 U510 ( .A(n681), .B(n357), .ZN(n366) );
  XNOR2_X1 U511 ( .A(n689), .B(n355), .ZN(n368) );
  NOR2_X2 U512 ( .A1(n607), .A2(n698), .ZN(n609) );
  XNOR2_X1 U513 ( .A(n375), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X2 U514 ( .A(n595), .B(n594), .ZN(n699) );
  XNOR2_X1 U515 ( .A(n376), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X1 U516 ( .A1(n506), .A2(n505), .ZN(n507) );
  XNOR2_X2 U517 ( .A(n468), .B(n449), .ZN(n705) );
  XNOR2_X1 U518 ( .A(n389), .B(n388), .ZN(n571) );
  INV_X1 U519 ( .A(KEYINPUT1), .ZN(n388) );
  NAND2_X1 U520 ( .A1(n501), .A2(n389), .ZN(n524) );
  NAND2_X1 U521 ( .A1(n507), .A2(n508), .ZN(n529) );
  XNOR2_X1 U522 ( .A(n573), .B(n572), .ZN(n675) );
  INV_X1 U523 ( .A(n726), .ZN(n403) );
  NAND2_X1 U524 ( .A1(n576), .A2(n406), .ZN(n405) );
  INV_X1 U525 ( .A(n577), .ZN(n406) );
  XNOR2_X1 U526 ( .A(n450), .B(n451), .ZN(n410) );
  XNOR2_X2 U527 ( .A(n411), .B(n448), .ZN(n468) );
  NAND2_X2 U528 ( .A1(n414), .A2(n412), .ZN(n574) );
  INV_X1 U529 ( .A(n556), .ZN(n413) );
  NAND2_X1 U530 ( .A1(n556), .A2(KEYINPUT0), .ZN(n415) );
  XNOR2_X2 U531 ( .A(n523), .B(n522), .ZN(n556) );
  NOR2_X1 U532 ( .A1(n555), .A2(KEYINPUT0), .ZN(n416) );
  NAND2_X1 U533 ( .A1(n555), .A2(KEYINPUT0), .ZN(n417) );
  XNOR2_X2 U534 ( .A(n446), .B(KEYINPUT4), .ZN(n462) );
  XNOR2_X2 U535 ( .A(n418), .B(n434), .ZN(n446) );
  XNOR2_X2 U536 ( .A(G143), .B(G128), .ZN(n418) );
  XNOR2_X2 U537 ( .A(n419), .B(n470), .ZN(n585) );
  XNOR2_X1 U538 ( .A(n497), .B(n420), .ZN(n602) );
  NOR2_X2 U539 ( .A1(n624), .A2(n550), .ZN(n646) );
  NAND2_X1 U540 ( .A1(n530), .A2(n643), .ZN(n523) );
  INV_X1 U541 ( .A(n530), .ZN(n547) );
  XNOR2_X1 U542 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U543 ( .A(n460), .B(G131), .ZN(n461) );
  INV_X1 U544 ( .A(KEYINPUT107), .ZN(n562) );
  XNOR2_X1 U545 ( .A(n491), .B(n490), .ZN(n492) );
  INV_X1 U546 ( .A(KEYINPUT77), .ZN(n434) );
  XNOR2_X1 U547 ( .A(n606), .B(n605), .ZN(n607) );
  XNOR2_X1 U548 ( .A(KEYINPUT89), .B(KEYINPUT63), .ZN(n608) );
  INV_X1 U549 ( .A(KEYINPUT2), .ZN(n635) );
  XOR2_X1 U550 ( .A(KEYINPUT85), .B(n596), .Z(n421) );
  XNOR2_X1 U551 ( .A(n423), .B(n422), .ZN(n431) );
  XNOR2_X1 U552 ( .A(n424), .B(KEYINPUT74), .ZN(n466) );
  NAND2_X1 U553 ( .A1(n466), .A2(G214), .ZN(n430) );
  XNOR2_X1 U554 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U555 ( .A(G113), .B(n427), .ZN(n429) );
  XNOR2_X1 U556 ( .A(G104), .B(n479), .ZN(n428) );
  NOR2_X1 U557 ( .A1(G902), .A2(n686), .ZN(n433) );
  XNOR2_X1 U558 ( .A(KEYINPUT13), .B(G475), .ZN(n432) );
  XNOR2_X1 U559 ( .A(n436), .B(n435), .ZN(n440) );
  XNOR2_X1 U560 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n437) );
  XNOR2_X1 U561 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U562 ( .A(n440), .B(n439), .Z(n443) );
  NAND2_X1 U563 ( .A1(n714), .A2(G234), .ZN(n441) );
  XOR2_X1 U564 ( .A(KEYINPUT8), .B(n441), .Z(n480) );
  NAND2_X1 U565 ( .A1(G217), .A2(n480), .ZN(n442) );
  XNOR2_X1 U566 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U567 ( .A(n446), .B(n444), .ZN(n692) );
  NOR2_X1 U568 ( .A1(G902), .A2(n692), .ZN(n445) );
  XNOR2_X1 U569 ( .A(G478), .B(n445), .ZN(n518) );
  INV_X1 U570 ( .A(n518), .ZN(n527) );
  NOR2_X1 U571 ( .A1(n528), .A2(n527), .ZN(n557) );
  INV_X1 U572 ( .A(n557), .ZN(n645) );
  INV_X1 U573 ( .A(n596), .ZN(n453) );
  XOR2_X1 U574 ( .A(G104), .B(G107), .Z(n447) );
  XNOR2_X1 U575 ( .A(G116), .B(G113), .ZN(n448) );
  NAND2_X1 U576 ( .A1(G224), .A2(n714), .ZN(n452) );
  NAND2_X1 U577 ( .A1(G210), .A2(n457), .ZN(n454) );
  XNOR2_X2 U578 ( .A(n456), .B(n455), .ZN(n530) );
  NAND2_X1 U579 ( .A1(G214), .A2(n457), .ZN(n643) );
  XOR2_X1 U580 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n465) );
  XNOR2_X1 U581 ( .A(G137), .B(KEYINPUT73), .ZN(n464) );
  NAND2_X1 U582 ( .A1(n466), .A2(G210), .ZN(n467) );
  XNOR2_X1 U583 ( .A(G472), .B(KEYINPUT97), .ZN(n470) );
  NAND2_X1 U584 ( .A1(G234), .A2(n596), .ZN(n471) );
  NAND2_X1 U585 ( .A1(G234), .A2(G237), .ZN(n472) );
  XNOR2_X1 U586 ( .A(n472), .B(KEYINPUT14), .ZN(n668) );
  NOR2_X1 U587 ( .A1(G902), .A2(n714), .ZN(n474) );
  NOR2_X1 U588 ( .A1(G953), .A2(G952), .ZN(n473) );
  NOR2_X1 U589 ( .A1(n474), .A2(n473), .ZN(n475) );
  AND2_X1 U590 ( .A1(n668), .A2(n475), .ZN(n554) );
  NAND2_X1 U591 ( .A1(G953), .A2(G900), .ZN(n476) );
  NAND2_X1 U592 ( .A1(n554), .A2(n476), .ZN(n477) );
  XOR2_X1 U593 ( .A(KEYINPUT79), .B(n477), .Z(n503) );
  NOR2_X1 U594 ( .A1(n655), .A2(n503), .ZN(n478) );
  XNOR2_X1 U595 ( .A(KEYINPUT68), .B(n478), .ZN(n494) );
  XOR2_X1 U596 ( .A(n479), .B(n496), .Z(n711) );
  NAND2_X1 U597 ( .A1(G221), .A2(n480), .ZN(n484) );
  XNOR2_X1 U598 ( .A(n711), .B(n486), .ZN(n696) );
  NAND2_X1 U599 ( .A1(G217), .A2(n487), .ZN(n491) );
  XOR2_X1 U600 ( .A(KEYINPUT75), .B(KEYINPUT92), .Z(n489) );
  XNOR2_X1 U601 ( .A(KEYINPUT25), .B(KEYINPUT76), .ZN(n488) );
  XNOR2_X1 U602 ( .A(n489), .B(n488), .ZN(n490) );
  NAND2_X1 U603 ( .A1(n494), .A2(n656), .ZN(n512) );
  NOR2_X1 U604 ( .A1(n585), .A2(n512), .ZN(n495) );
  XNOR2_X1 U605 ( .A(KEYINPUT28), .B(n495), .ZN(n501) );
  NAND2_X1 U606 ( .A1(G227), .A2(n714), .ZN(n499) );
  NOR2_X1 U607 ( .A1(n674), .A2(n524), .ZN(n502) );
  XNOR2_X1 U608 ( .A(n502), .B(KEYINPUT42), .ZN(n730) );
  INV_X1 U609 ( .A(n503), .ZN(n508) );
  XOR2_X1 U610 ( .A(KEYINPUT94), .B(n655), .Z(n558) );
  NAND2_X1 U611 ( .A1(n558), .A2(n566), .ZN(n570) );
  INV_X1 U612 ( .A(n570), .ZN(n651) );
  XNOR2_X1 U613 ( .A(n586), .B(KEYINPUT109), .ZN(n506) );
  NAND2_X1 U614 ( .A1(n518), .A2(n528), .ZN(n509) );
  XOR2_X1 U615 ( .A(n509), .B(KEYINPUT103), .Z(n515) );
  XNOR2_X1 U616 ( .A(n511), .B(KEYINPUT46), .ZN(n541) );
  XNOR2_X1 U617 ( .A(n585), .B(KEYINPUT6), .ZN(n578) );
  INV_X1 U618 ( .A(n512), .ZN(n513) );
  NAND2_X1 U619 ( .A1(n513), .A2(n643), .ZN(n514) );
  NOR2_X1 U620 ( .A1(n515), .A2(n514), .ZN(n516) );
  NAND2_X1 U621 ( .A1(n578), .A2(n516), .ZN(n544) );
  INV_X1 U622 ( .A(n571), .ZN(n652) );
  NOR2_X1 U623 ( .A1(n528), .A2(n518), .ZN(n626) );
  XNOR2_X1 U624 ( .A(KEYINPUT104), .B(n626), .ZN(n550) );
  XNOR2_X1 U625 ( .A(n646), .B(KEYINPUT82), .ZN(n589) );
  INV_X1 U626 ( .A(KEYINPUT47), .ZN(n534) );
  XOR2_X1 U627 ( .A(KEYINPUT66), .B(n534), .Z(n519) );
  NOR2_X1 U628 ( .A1(n589), .A2(n519), .ZN(n520) );
  XNOR2_X1 U629 ( .A(n520), .B(KEYINPUT72), .ZN(n521) );
  NOR2_X1 U630 ( .A1(KEYINPUT81), .A2(n521), .ZN(n526) );
  INV_X1 U631 ( .A(KEYINPUT19), .ZN(n522) );
  INV_X1 U632 ( .A(n622), .ZN(n525) );
  NOR2_X1 U633 ( .A1(n526), .A2(n525), .ZN(n538) );
  NAND2_X1 U634 ( .A1(KEYINPUT81), .A2(n534), .ZN(n532) );
  NAND2_X1 U635 ( .A1(n528), .A2(n527), .ZN(n577) );
  NOR2_X1 U636 ( .A1(n577), .A2(n529), .ZN(n531) );
  NAND2_X1 U637 ( .A1(n531), .A2(n530), .ZN(n621) );
  NAND2_X1 U638 ( .A1(n532), .A2(n621), .ZN(n537) );
  NOR2_X1 U639 ( .A1(n622), .A2(KEYINPUT81), .ZN(n533) );
  NOR2_X1 U640 ( .A1(n646), .A2(n533), .ZN(n535) );
  NOR2_X1 U641 ( .A1(n535), .A2(n534), .ZN(n536) );
  AND2_X1 U642 ( .A1(n723), .A2(n539), .ZN(n540) );
  NAND2_X1 U643 ( .A1(n541), .A2(n540), .ZN(n543) );
  XNOR2_X1 U644 ( .A(n543), .B(n542), .ZN(n549) );
  XOR2_X1 U645 ( .A(n544), .B(KEYINPUT108), .Z(n545) );
  NAND2_X1 U646 ( .A1(n545), .A2(n571), .ZN(n546) );
  XNOR2_X1 U647 ( .A(KEYINPUT43), .B(n546), .ZN(n548) );
  NAND2_X1 U648 ( .A1(n548), .A2(n547), .ZN(n631) );
  NAND2_X1 U649 ( .A1(n549), .A2(n631), .ZN(n599) );
  NAND2_X1 U650 ( .A1(n551), .A2(n550), .ZN(n629) );
  INV_X1 U651 ( .A(n629), .ZN(n552) );
  NOR2_X2 U652 ( .A1(n599), .A2(n552), .ZN(n713) );
  NAND2_X1 U653 ( .A1(G898), .A2(G953), .ZN(n553) );
  NAND2_X1 U654 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U655 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X2 U656 ( .A1(n565), .A2(n652), .ZN(n580) );
  XNOR2_X1 U657 ( .A(n580), .B(n562), .ZN(n563) );
  NAND2_X1 U658 ( .A1(n563), .A2(n585), .ZN(n564) );
  NOR2_X1 U659 ( .A1(n565), .A2(n571), .ZN(n568) );
  NOR2_X1 U660 ( .A1(n566), .A2(n578), .ZN(n567) );
  NAND2_X1 U661 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U662 ( .A(KEYINPUT33), .B(KEYINPUT70), .Z(n573) );
  NOR2_X1 U663 ( .A1(n571), .A2(n570), .ZN(n583) );
  NAND2_X1 U664 ( .A1(n583), .A2(n578), .ZN(n572) );
  NOR2_X1 U665 ( .A1(n675), .A2(n574), .ZN(n575) );
  XNOR2_X1 U666 ( .A(n575), .B(KEYINPUT34), .ZN(n576) );
  NOR2_X1 U667 ( .A1(n656), .A2(n578), .ZN(n579) );
  NAND2_X1 U668 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U669 ( .A(KEYINPUT105), .B(n581), .ZN(n727) );
  NAND2_X1 U670 ( .A1(n582), .A2(n583), .ZN(n661) );
  NOR2_X1 U671 ( .A1(n574), .A2(n661), .ZN(n584) );
  XOR2_X1 U672 ( .A(KEYINPUT31), .B(n584), .Z(n627) );
  NAND2_X1 U673 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U674 ( .A1(n574), .A2(n587), .ZN(n611) );
  NOR2_X1 U675 ( .A1(n627), .A2(n611), .ZN(n588) );
  NOR2_X1 U676 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U677 ( .A1(n727), .A2(n590), .ZN(n591) );
  XOR2_X1 U678 ( .A(KEYINPUT106), .B(n591), .Z(n592) );
  NOR2_X2 U679 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U680 ( .A1(KEYINPUT2), .A2(n629), .ZN(n597) );
  XNOR2_X1 U681 ( .A(KEYINPUT80), .B(n597), .ZN(n598) );
  XNOR2_X1 U682 ( .A(KEYINPUT86), .B(n600), .ZN(n601) );
  XNOR2_X1 U683 ( .A(n602), .B(KEYINPUT113), .ZN(n604) );
  XOR2_X1 U684 ( .A(KEYINPUT62), .B(KEYINPUT114), .Z(n603) );
  XNOR2_X1 U685 ( .A(n609), .B(n608), .ZN(G57) );
  NAND2_X1 U686 ( .A1(n611), .A2(n624), .ZN(n610) );
  XNOR2_X1 U687 ( .A(n610), .B(G104), .ZN(G6) );
  XOR2_X1 U688 ( .A(KEYINPUT115), .B(KEYINPUT27), .Z(n613) );
  NAND2_X1 U689 ( .A1(n611), .A2(n626), .ZN(n612) );
  XNOR2_X1 U690 ( .A(n613), .B(n612), .ZN(n615) );
  XOR2_X1 U691 ( .A(G107), .B(KEYINPUT26), .Z(n614) );
  XNOR2_X1 U692 ( .A(n615), .B(n614), .ZN(G9) );
  XNOR2_X1 U693 ( .A(G110), .B(KEYINPUT116), .ZN(n617) );
  XNOR2_X1 U694 ( .A(n617), .B(n616), .ZN(G12) );
  XOR2_X1 U695 ( .A(G128), .B(KEYINPUT29), .Z(n619) );
  NAND2_X1 U696 ( .A1(n622), .A2(n626), .ZN(n618) );
  XNOR2_X1 U697 ( .A(n619), .B(n618), .ZN(G30) );
  XOR2_X1 U698 ( .A(G143), .B(KEYINPUT117), .Z(n620) );
  XNOR2_X1 U699 ( .A(n621), .B(n620), .ZN(G45) );
  NAND2_X1 U700 ( .A1(n622), .A2(n624), .ZN(n623) );
  XNOR2_X1 U701 ( .A(n623), .B(G146), .ZN(G48) );
  NAND2_X1 U702 ( .A1(n627), .A2(n624), .ZN(n625) );
  XNOR2_X1 U703 ( .A(n625), .B(G113), .ZN(G15) );
  NAND2_X1 U704 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U705 ( .A(n628), .B(G116), .ZN(G18) );
  XOR2_X1 U706 ( .A(G134), .B(n629), .Z(n630) );
  XNOR2_X1 U707 ( .A(n630), .B(KEYINPUT119), .ZN(G36) );
  XNOR2_X1 U708 ( .A(G140), .B(KEYINPUT120), .ZN(n632) );
  XNOR2_X1 U709 ( .A(n632), .B(n631), .ZN(G42) );
  XNOR2_X1 U710 ( .A(n633), .B(KEYINPUT83), .ZN(n637) );
  INV_X1 U711 ( .A(n699), .ZN(n634) );
  NAND2_X1 U712 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n637), .A2(n636), .ZN(n639) );
  XNOR2_X1 U714 ( .A(n641), .B(n640), .ZN(n673) );
  NOR2_X1 U715 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U716 ( .A1(n645), .A2(n644), .ZN(n649) );
  NOR2_X1 U717 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U718 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U719 ( .A1(n675), .A2(n650), .ZN(n666) );
  NOR2_X1 U720 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U721 ( .A(n653), .B(KEYINPUT50), .ZN(n654) );
  XNOR2_X1 U722 ( .A(n654), .B(KEYINPUT121), .ZN(n660) );
  AND2_X1 U723 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U724 ( .A(KEYINPUT49), .B(n657), .Z(n658) );
  NOR2_X1 U725 ( .A1(n582), .A2(n658), .ZN(n659) );
  NAND2_X1 U726 ( .A1(n660), .A2(n659), .ZN(n662) );
  NAND2_X1 U727 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U728 ( .A(KEYINPUT51), .B(n663), .ZN(n664) );
  NOR2_X1 U729 ( .A1(n664), .A2(n674), .ZN(n665) );
  NOR2_X1 U730 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U731 ( .A(KEYINPUT52), .B(n667), .ZN(n670) );
  NAND2_X1 U732 ( .A1(G952), .A2(n668), .ZN(n669) );
  NOR2_X1 U733 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U734 ( .A1(G953), .A2(n671), .ZN(n672) );
  XNOR2_X1 U735 ( .A(KEYINPUT53), .B(n676), .ZN(G75) );
  NAND2_X1 U736 ( .A1(n690), .A2(G210), .ZN(n681) );
  XOR2_X1 U737 ( .A(KEYINPUT90), .B(KEYINPUT55), .Z(n678) );
  XNOR2_X1 U738 ( .A(KEYINPUT122), .B(KEYINPUT54), .ZN(n677) );
  XNOR2_X1 U739 ( .A(n678), .B(n677), .ZN(n679) );
  XOR2_X1 U740 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n683) );
  NAND2_X1 U741 ( .A1(n694), .A2(G469), .ZN(n682) );
  NOR2_X1 U742 ( .A1(n698), .A2(n685), .ZN(G54) );
  XNOR2_X1 U743 ( .A(KEYINPUT59), .B(KEYINPUT123), .ZN(n688) );
  XNOR2_X1 U744 ( .A(n686), .B(KEYINPUT124), .ZN(n687) );
  NAND2_X1 U745 ( .A1(n690), .A2(G475), .ZN(n689) );
  NAND2_X1 U746 ( .A1(G478), .A2(n694), .ZN(n691) );
  XNOR2_X1 U747 ( .A(n692), .B(n691), .ZN(n693) );
  NOR2_X1 U748 ( .A1(n698), .A2(n693), .ZN(G63) );
  NAND2_X1 U749 ( .A1(G217), .A2(n694), .ZN(n695) );
  XNOR2_X1 U750 ( .A(n696), .B(n695), .ZN(n697) );
  NOR2_X1 U751 ( .A1(n698), .A2(n697), .ZN(G66) );
  NAND2_X1 U752 ( .A1(n714), .A2(n699), .ZN(n703) );
  NAND2_X1 U753 ( .A1(G953), .A2(G224), .ZN(n700) );
  XNOR2_X1 U754 ( .A(KEYINPUT61), .B(n700), .ZN(n701) );
  NAND2_X1 U755 ( .A1(n701), .A2(G898), .ZN(n702) );
  NAND2_X1 U756 ( .A1(n703), .A2(n702), .ZN(n709) );
  XOR2_X1 U757 ( .A(n705), .B(n704), .Z(n707) );
  NOR2_X1 U758 ( .A1(G898), .A2(n714), .ZN(n706) );
  NOR2_X1 U759 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U760 ( .A(n709), .B(n708), .ZN(n710) );
  XOR2_X1 U761 ( .A(KEYINPUT125), .B(n710), .Z(G69) );
  XOR2_X1 U762 ( .A(n712), .B(n711), .Z(n717) );
  XOR2_X1 U763 ( .A(n717), .B(n713), .Z(n715) );
  NAND2_X1 U764 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U765 ( .A(n716), .B(KEYINPUT126), .ZN(n722) );
  XNOR2_X1 U766 ( .A(G227), .B(n717), .ZN(n718) );
  NAND2_X1 U767 ( .A1(n718), .A2(G900), .ZN(n719) );
  XOR2_X1 U768 ( .A(KEYINPUT127), .B(n719), .Z(n720) );
  NAND2_X1 U769 ( .A1(n720), .A2(G953), .ZN(n721) );
  NAND2_X1 U770 ( .A1(n722), .A2(n721), .ZN(G72) );
  XOR2_X1 U771 ( .A(KEYINPUT37), .B(KEYINPUT118), .Z(n725) );
  XNOR2_X1 U772 ( .A(G125), .B(n723), .ZN(n724) );
  XNOR2_X1 U773 ( .A(n725), .B(n724), .ZN(G27) );
  XNOR2_X1 U774 ( .A(G119), .B(n726), .ZN(G21) );
  XOR2_X1 U775 ( .A(G101), .B(n727), .Z(G3) );
  XOR2_X1 U776 ( .A(n728), .B(G122), .Z(G24) );
  XOR2_X1 U777 ( .A(n729), .B(G131), .Z(G33) );
  XOR2_X1 U778 ( .A(G137), .B(n730), .Z(G39) );
endmodule

