//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 1 0 0 0 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n823, new_n825, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G57gat), .ZN(new_n204));
  INV_X1    g003(.A(G85gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G225gat), .A2(G233gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G113gat), .B(G120gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n211));
  INV_X1    g010(.A(G134gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G127gat), .ZN(new_n213));
  INV_X1    g012(.A(G127gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G134gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  OR2_X1    g015(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n211), .A2(new_n218), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n216), .B(new_n217), .C1(new_n210), .C2(KEYINPUT1), .ZN(new_n220));
  NAND2_X1  g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221));
  INV_X1    g020(.A(G155gat), .ZN(new_n222));
  INV_X1    g021(.A(G162gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G141gat), .B(G148gat), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n221), .B(new_n224), .C1(new_n225), .C2(KEYINPUT2), .ZN(new_n226));
  XOR2_X1   g025(.A(G141gat), .B(G148gat), .Z(new_n227));
  NAND2_X1  g026(.A1(new_n224), .A2(new_n221), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n221), .A2(KEYINPUT2), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  AND4_X1   g029(.A1(new_n219), .A2(new_n220), .A3(new_n226), .A4(new_n230), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n219), .A2(new_n220), .B1(new_n230), .B2(new_n226), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n209), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT5), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n219), .A2(new_n220), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n230), .A2(new_n226), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT4), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n235), .A2(KEYINPUT76), .A3(new_n236), .A4(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT76), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n219), .A2(new_n220), .A3(new_n226), .A4(new_n230), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n240), .B2(KEYINPUT4), .ZN(new_n241));
  XOR2_X1   g040(.A(KEYINPUT75), .B(KEYINPUT4), .Z(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n238), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n230), .A2(new_n226), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n245), .B1(new_n230), .B2(new_n226), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n219), .A2(new_n220), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n209), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n234), .B1(new_n244), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n246), .ZN(new_n252));
  INV_X1    g051(.A(new_n247), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(new_n249), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n240), .A2(new_n237), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n231), .A2(new_n242), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n209), .A2(KEYINPUT5), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n254), .A2(new_n255), .A3(new_n256), .A4(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n207), .B1(new_n251), .B2(new_n259), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n244), .A2(new_n250), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n206), .B(new_n258), .C1(new_n261), .C2(new_n234), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT6), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n260), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT79), .ZN(new_n265));
  OR2_X1    g064(.A1(new_n260), .A2(new_n263), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT79), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n260), .A2(new_n262), .A3(new_n267), .A4(new_n263), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n265), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G226gat), .ZN(new_n270));
  INV_X1    g069(.A(G233gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n272), .A2(KEYINPUT29), .ZN(new_n273));
  INV_X1    g072(.A(G169gat), .ZN(new_n274));
  INV_X1    g073(.A(G176gat), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT67), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT67), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n277), .A2(G169gat), .A3(G176gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n274), .A2(new_n275), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT23), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT25), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT66), .B(G176gat), .ZN(new_n284));
  NOR3_X1   g083(.A1(new_n284), .A2(new_n281), .A3(G169gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(G183gat), .A2(G190gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT24), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G183gat), .ZN(new_n290));
  INV_X1    g089(.A(G190gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n291), .A3(KEYINPUT65), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT65), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(G183gat), .B2(G190gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n289), .A2(new_n292), .A3(new_n294), .A4(new_n295), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n289), .B(new_n295), .C1(G183gat), .C2(G190gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(G169gat), .A2(G176gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT23), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n280), .A2(new_n281), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n297), .A2(new_n279), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  AOI22_X1  g100(.A1(new_n286), .A2(new_n296), .B1(KEYINPUT25), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n280), .A2(KEYINPUT26), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT26), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT68), .B1(new_n298), .B2(new_n304), .ZN(new_n305));
  AND4_X1   g104(.A1(KEYINPUT68), .A2(new_n304), .A3(new_n274), .A4(new_n275), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n279), .B(new_n303), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT27), .B(G183gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(new_n291), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT28), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT28), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n308), .A2(new_n311), .A3(new_n291), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n307), .A2(new_n287), .A3(new_n310), .A4(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT73), .B1(new_n302), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n301), .A2(KEYINPUT25), .ZN(new_n315));
  INV_X1    g114(.A(new_n284), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n316), .A2(KEYINPUT23), .A3(new_n274), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n317), .A2(new_n279), .A3(new_n296), .A4(new_n282), .ZN(new_n318));
  AND4_X1   g117(.A1(KEYINPUT73), .A2(new_n313), .A3(new_n315), .A4(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n273), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G197gat), .B(G204gat), .ZN(new_n321));
  INV_X1    g120(.A(G211gat), .ZN(new_n322));
  INV_X1    g121(.A(G218gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n321), .B1(KEYINPUT22), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G211gat), .B(G218gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n313), .A2(new_n315), .A3(new_n318), .ZN(new_n328));
  NOR3_X1   g127(.A1(new_n328), .A2(new_n270), .A3(new_n271), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n320), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT74), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT37), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT73), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n328), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n302), .A2(KEYINPUT73), .A3(new_n313), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(new_n337), .A3(new_n272), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n328), .A2(new_n273), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n327), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n320), .A2(new_n330), .A3(KEYINPUT74), .A4(new_n327), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n333), .A2(new_n334), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT38), .ZN(new_n345));
  XNOR2_X1  g144(.A(G8gat), .B(G36gat), .ZN(new_n346));
  INV_X1    g145(.A(G64gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(G92gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n340), .A2(new_n327), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n320), .A2(new_n330), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n351), .B(KEYINPUT37), .C1(new_n327), .C2(new_n352), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n344), .A2(new_n345), .A3(new_n350), .A4(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT80), .ZN(new_n355));
  INV_X1    g154(.A(new_n350), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n333), .A2(new_n342), .A3(new_n343), .A4(new_n356), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n269), .A2(new_n354), .A3(new_n355), .A4(new_n357), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n265), .A2(new_n266), .A3(new_n357), .A4(new_n268), .ZN(new_n359));
  INV_X1    g158(.A(new_n354), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT80), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n333), .A2(new_n342), .A3(new_n343), .ZN(new_n362));
  AND2_X1   g161(.A1(new_n362), .A2(KEYINPUT37), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n344), .A2(new_n350), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT38), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n358), .A2(new_n361), .A3(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n327), .B1(new_n246), .B2(KEYINPUT29), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT3), .B1(new_n341), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n367), .B1(new_n369), .B2(new_n236), .ZN(new_n370));
  NAND2_X1  g169(.A1(G228gat), .A2(G233gat), .ZN(new_n371));
  XOR2_X1   g170(.A(new_n370), .B(new_n371), .Z(new_n372));
  XNOR2_X1  g171(.A(G78gat), .B(G106gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT31), .B(G50gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT77), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n376), .A3(G22gat), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n377), .B1(G22gat), .B2(new_n375), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n372), .B(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n350), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(KEYINPUT30), .A3(new_n357), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n333), .A2(new_n343), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT30), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n382), .A2(new_n383), .A3(new_n342), .A4(new_n356), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(new_n209), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT78), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT39), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n387), .B(KEYINPUT78), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n231), .A2(new_n232), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n390), .B1(new_n393), .B2(new_n208), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n391), .A2(new_n395), .A3(new_n206), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT40), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n396), .A2(new_n397), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n385), .A2(new_n399), .A3(new_n260), .A4(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n366), .A2(new_n379), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT72), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT34), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT32), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n313), .A2(new_n235), .A3(new_n315), .A4(new_n318), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT70), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n302), .A2(KEYINPUT70), .A3(new_n235), .A4(new_n313), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n328), .A2(new_n249), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G227gat), .A2(G233gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT64), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n406), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT33), .B1(new_n412), .B2(new_n414), .ZN(new_n416));
  XOR2_X1   g215(.A(G15gat), .B(G43gat), .Z(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(KEYINPUT71), .ZN(new_n418));
  XOR2_X1   g217(.A(G71gat), .B(G99gat), .Z(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NOR3_X1   g220(.A1(new_n415), .A2(new_n416), .A3(new_n421), .ZN(new_n422));
  AOI221_X4 g221(.A(new_n406), .B1(KEYINPUT33), .B2(new_n420), .C1(new_n412), .C2(new_n414), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n405), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  OAI22_X1  g223(.A1(new_n412), .A2(new_n414), .B1(new_n403), .B2(KEYINPUT34), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n412), .A2(new_n414), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT33), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n421), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n415), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n423), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n432), .A3(new_n404), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n424), .A2(new_n426), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n426), .B1(new_n424), .B2(new_n433), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT36), .ZN(new_n436));
  NOR3_X1   g235(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n381), .A2(new_n384), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n266), .A2(new_n264), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n379), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n422), .A2(new_n405), .A3(new_n423), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n404), .B1(new_n431), .B2(new_n432), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n425), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n424), .A2(new_n426), .A3(new_n433), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT36), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n437), .A2(new_n440), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n443), .A2(new_n444), .ZN(new_n447));
  INV_X1    g246(.A(new_n439), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n448), .B1(new_n381), .B2(new_n384), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n449), .A3(new_n379), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT35), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT81), .B(KEYINPUT35), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n452), .B1(new_n381), .B2(new_n384), .ZN(new_n453));
  INV_X1    g252(.A(new_n269), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n447), .A2(new_n379), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n402), .A2(new_n446), .B1(new_n451), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(G43gat), .B(G50gat), .ZN(new_n457));
  NOR2_X1   g256(.A1(G29gat), .A2(G36gat), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n458), .A2(KEYINPUT14), .ZN(new_n459));
  INV_X1    g258(.A(new_n458), .ZN(new_n460));
  INV_X1    g259(.A(G29gat), .ZN(new_n461));
  INV_X1    g260(.A(G36gat), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT14), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n459), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n464), .A2(KEYINPUT15), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n464), .A2(KEYINPUT15), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n457), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n464), .A2(KEYINPUT15), .ZN(new_n468));
  INV_X1    g267(.A(new_n457), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT17), .ZN(new_n472));
  XNOR2_X1  g271(.A(G15gat), .B(G22gat), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT16), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n473), .B1(new_n474), .B2(G1gat), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n475), .B1(G1gat), .B2(new_n473), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n476), .B(G8gat), .ZN(new_n477));
  OR2_X1    g276(.A1(new_n477), .A2(KEYINPUT83), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(KEYINPUT83), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT17), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n467), .A2(new_n480), .A3(new_n470), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n472), .A2(new_n478), .A3(new_n479), .A4(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(G8gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n476), .B(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT85), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT85), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n477), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n485), .A2(new_n487), .A3(new_n467), .A4(new_n470), .ZN(new_n488));
  NAND2_X1  g287(.A1(G229gat), .A2(G233gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(KEYINPUT84), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n482), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT18), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n485), .A2(new_n487), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n471), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n488), .ZN(new_n497));
  XOR2_X1   g296(.A(new_n490), .B(KEYINPUT13), .Z(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n482), .A2(KEYINPUT18), .A3(new_n488), .A4(new_n491), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n494), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(G169gat), .B(G197gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(G113gat), .B(G141gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n507), .B(KEYINPUT12), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n502), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n494), .A2(new_n500), .A3(new_n508), .A4(new_n501), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n456), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(G57gat), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n515), .A2(KEYINPUT89), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n515), .A2(KEYINPUT89), .ZN(new_n517));
  OAI21_X1  g316(.A(G64gat), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n515), .A2(G64gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT90), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n520), .B(G64gat), .C1(new_n516), .C2(new_n517), .ZN(new_n523));
  INV_X1    g322(.A(G71gat), .ZN(new_n524));
  INV_X1    g323(.A(G78gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(new_n525), .A3(KEYINPUT9), .ZN(new_n526));
  NAND2_X1  g325(.A1(G71gat), .A2(G78gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n522), .A2(new_n523), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n347), .A2(G57gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n515), .A2(G64gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OR2_X1    g331(.A1(KEYINPUT86), .A2(KEYINPUT9), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT87), .B1(G71gat), .B2(G78gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT87), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n535), .A2(new_n524), .A3(new_n525), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n532), .A2(new_n533), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT86), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n527), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(KEYINPUT86), .A2(G71gat), .A3(G78gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT88), .B1(new_n537), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n347), .A2(G57gat), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n533), .B1(new_n519), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n536), .A2(new_n534), .ZN(new_n545));
  AND4_X1   g344(.A1(KEYINPUT88), .A2(new_n544), .A3(new_n541), .A4(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n529), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n547), .A2(KEYINPUT91), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n544), .A2(new_n541), .A3(new_n545), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT88), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n537), .A2(KEYINPUT88), .A3(new_n541), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n518), .A2(new_n521), .B1(new_n527), .B2(new_n526), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n551), .A2(new_n552), .B1(new_n553), .B2(new_n523), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT91), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT21), .B1(new_n548), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n495), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n554), .A2(KEYINPUT21), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(new_n214), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n558), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n562));
  XNOR2_X1  g361(.A(G155gat), .B(G183gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n561), .B(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(new_n322), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n565), .B(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G85gat), .A2(G92gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT7), .ZN(new_n571));
  NAND2_X1  g370(.A1(G99gat), .A2(G106gat), .ZN(new_n572));
  AOI22_X1  g371(.A1(KEYINPUT8), .A2(new_n572), .B1(new_n205), .B2(new_n349), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G99gat), .B(G106gat), .Z(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n575), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n577), .A2(new_n573), .A3(new_n571), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n472), .A2(new_n481), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT41), .ZN(new_n581));
  NAND2_X1  g380(.A1(G232gat), .A2(G233gat), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n582), .B(KEYINPUT92), .Z(new_n583));
  OAI221_X1 g382(.A(new_n580), .B1(new_n581), .B2(new_n583), .C1(new_n471), .C2(new_n579), .ZN(new_n584));
  XOR2_X1   g383(.A(KEYINPUT93), .B(G134gat), .Z(new_n585));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n584), .B(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n583), .A2(new_n581), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(new_n223), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n588), .B(new_n590), .Z(new_n591));
  INV_X1    g390(.A(KEYINPUT10), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n578), .A2(KEYINPUT95), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(new_n576), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n574), .A2(KEYINPUT95), .A3(new_n575), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n554), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n576), .A2(new_n578), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT94), .ZN(new_n598));
  NOR3_X1   g397(.A1(new_n554), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT94), .B1(new_n547), .B2(new_n579), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n592), .B(new_n596), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  OAI211_X1 g400(.A(KEYINPUT10), .B(new_n597), .C1(new_n548), .C2(new_n556), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G230gat), .A2(G233gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G120gat), .B(G148gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(new_n275), .ZN(new_n607));
  INV_X1    g406(.A(G204gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n596), .B1(new_n599), .B2(new_n600), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n611), .A2(G230gat), .A3(G233gat), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n605), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT96), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n605), .A2(KEYINPUT96), .A3(new_n610), .A4(new_n612), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n604), .B(KEYINPUT97), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n619), .B1(new_n601), .B2(new_n602), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(new_n612), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(new_n609), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n617), .A2(new_n623), .ZN(new_n624));
  NOR3_X1   g423(.A1(new_n569), .A2(new_n591), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n514), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n626), .A2(new_n439), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT98), .B(G1gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(G1324gat));
  INV_X1    g428(.A(new_n626), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n483), .B1(new_n630), .B2(new_n385), .ZN(new_n631));
  NOR2_X1   g430(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n474), .A2(new_n483), .ZN(new_n633));
  NOR4_X1   g432(.A1(new_n626), .A2(new_n438), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(KEYINPUT42), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n635), .B1(KEYINPUT42), .B2(new_n634), .ZN(G1325gat));
  INV_X1    g435(.A(G15gat), .ZN(new_n637));
  INV_X1    g436(.A(new_n447), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n637), .B1(new_n626), .B2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT99), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n437), .A2(new_n445), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n626), .A2(new_n637), .A3(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n640), .A2(new_n642), .ZN(G1326gat));
  INV_X1    g442(.A(new_n379), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n630), .A2(KEYINPUT100), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT100), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(new_n626), .B2(new_n379), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT43), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G22gat), .ZN(G1327gat));
  NOR2_X1   g449(.A1(new_n568), .A2(new_n624), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n514), .A2(new_n591), .A3(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n652), .A2(G29gat), .A3(new_n439), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n653), .B(KEYINPUT45), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n588), .B(new_n590), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n402), .A2(new_n446), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n451), .A2(new_n455), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT44), .B1(new_n658), .B2(KEYINPUT102), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT44), .ZN(new_n661));
  NOR4_X1   g460(.A1(new_n456), .A2(new_n660), .A3(new_n661), .A4(new_n655), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT101), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n512), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n510), .A2(KEYINPUT101), .A3(new_n511), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n663), .A2(new_n668), .A3(new_n651), .ZN(new_n669));
  OAI21_X1  g468(.A(G29gat), .B1(new_n669), .B2(new_n439), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n670), .ZN(G1328gat));
  NOR3_X1   g470(.A1(new_n652), .A2(G36gat), .A3(new_n438), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT46), .ZN(new_n673));
  OAI21_X1  g472(.A(G36gat), .B1(new_n669), .B2(new_n438), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n675), .B(KEYINPUT103), .Z(G1329gat));
  OR3_X1    g475(.A1(new_n669), .A2(KEYINPUT105), .A3(new_n641), .ZN(new_n677));
  OAI21_X1  g476(.A(KEYINPUT105), .B1(new_n669), .B2(new_n641), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n677), .A2(G43gat), .A3(new_n678), .ZN(new_n679));
  OR3_X1    g478(.A1(new_n652), .A2(G43gat), .A3(new_n638), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(KEYINPUT47), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(G43gat), .B1(new_n669), .B2(new_n641), .ZN(new_n682));
  AOI21_X1  g481(.A(KEYINPUT47), .B1(new_n682), .B2(new_n680), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(KEYINPUT104), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n685));
  AOI211_X1 g484(.A(new_n685), .B(KEYINPUT47), .C1(new_n682), .C2(new_n680), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n681), .B1(new_n684), .B2(new_n686), .ZN(G1330gat));
  NAND2_X1  g486(.A1(new_n644), .A2(G50gat), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n652), .A2(new_n379), .ZN(new_n689));
  OAI22_X1  g488(.A1(new_n669), .A2(new_n688), .B1(G50gat), .B2(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g490(.A(new_n624), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n568), .A2(new_n655), .A3(new_n667), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n456), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n448), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n516), .A2(new_n517), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1332gat));
  INV_X1    g496(.A(new_n694), .ZN(new_n698));
  AOI211_X1 g497(.A(new_n438), .B(new_n698), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n699));
  NOR2_X1   g498(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT108), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n699), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(KEYINPUT106), .B(KEYINPUT107), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1333gat));
  OAI21_X1  g503(.A(G71gat), .B1(new_n698), .B2(new_n641), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n694), .A2(new_n524), .A3(new_n447), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g507(.A1(new_n694), .A2(new_n644), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(G78gat), .ZN(G1335gat));
  OAI21_X1  g509(.A(new_n436), .B1(new_n434), .B2(new_n435), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n443), .A2(KEYINPUT36), .A3(new_n444), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n711), .B(new_n712), .C1(new_n449), .C2(new_n379), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n400), .A2(new_n260), .A3(new_n381), .A4(new_n384), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(new_n398), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(new_n644), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n713), .B1(new_n716), .B2(new_n366), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n638), .A2(new_n644), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n453), .A2(new_n454), .ZN(new_n719));
  AOI22_X1  g518(.A1(new_n718), .A2(new_n719), .B1(new_n450), .B2(KEYINPUT35), .ZN(new_n720));
  OAI211_X1 g519(.A(KEYINPUT102), .B(new_n591), .C1(new_n717), .C2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n661), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n658), .A2(KEYINPUT102), .A3(KEYINPUT44), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n668), .A2(new_n568), .A3(new_n692), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(KEYINPUT109), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n722), .A2(new_n723), .A3(new_n727), .A4(new_n724), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n439), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(KEYINPUT110), .B1(new_n456), .B2(new_n655), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT110), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n731), .B(new_n591), .C1(new_n717), .C2(new_n720), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n668), .A2(new_n568), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n730), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT51), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n730), .A2(new_n732), .A3(KEYINPUT51), .A4(new_n733), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n624), .A2(new_n205), .A3(new_n448), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT111), .ZN(new_n741));
  OAI22_X1  g540(.A1(new_n729), .A2(new_n205), .B1(new_n739), .B2(new_n741), .ZN(G1336gat));
  AOI21_X1  g541(.A(new_n727), .B1(new_n663), .B2(new_n724), .ZN(new_n743));
  INV_X1    g542(.A(new_n728), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n385), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n745), .A2(KEYINPUT112), .A3(G92gat), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n692), .B1(new_n736), .B2(new_n737), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n747), .A2(new_n349), .A3(new_n385), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT112), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n438), .B1(new_n726), .B2(new_n728), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n750), .B2(new_n349), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n746), .A2(new_n748), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT52), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754));
  OAI21_X1  g553(.A(G92gat), .B1(new_n725), .B2(new_n438), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n748), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n753), .A2(new_n756), .ZN(G1337gat));
  AOI21_X1  g556(.A(G99gat), .B1(new_n747), .B2(new_n447), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n641), .B1(new_n726), .B2(new_n728), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n758), .B1(G99gat), .B2(new_n759), .ZN(G1338gat));
  INV_X1    g559(.A(G106gat), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n738), .A2(new_n761), .A3(new_n644), .A4(new_n624), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n379), .B1(new_n726), .B2(new_n728), .ZN(new_n763));
  XNOR2_X1  g562(.A(KEYINPUT113), .B(G106gat), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n762), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(KEYINPUT53), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT114), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XOR2_X1   g568(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n770));
  NAND3_X1  g569(.A1(new_n663), .A2(new_n644), .A3(new_n724), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(new_n764), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n762), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n772), .A2(new_n762), .A3(KEYINPUT116), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n766), .A2(KEYINPUT114), .A3(KEYINPUT53), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n769), .A2(new_n777), .A3(new_n778), .ZN(G1339gat));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n610), .B1(new_n620), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n601), .A2(new_n602), .A3(new_n619), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n605), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n782), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT54), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n781), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI211_X1 g588(.A(KEYINPUT55), .B(new_n781), .C1(new_n784), .C2(new_n786), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(new_n617), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n789), .A2(KEYINPUT118), .A3(new_n617), .A4(new_n790), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n667), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n497), .A2(new_n499), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n491), .B1(new_n482), .B2(new_n488), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n507), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n511), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n624), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n624), .A2(KEYINPUT119), .A3(new_n800), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n655), .B1(new_n795), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n793), .A2(new_n794), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n807), .A2(new_n591), .A3(new_n800), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n569), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n693), .A2(new_n624), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n813), .A2(new_n718), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n385), .A2(new_n439), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(G113gat), .B1(new_n816), .B2(new_n513), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n816), .A2(G113gat), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n817), .B1(new_n818), .B2(new_n667), .ZN(G1340gat));
  INV_X1    g618(.A(new_n816), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n624), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(G120gat), .ZN(G1341gat));
  NOR2_X1   g621(.A1(new_n816), .A2(new_n569), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(new_n214), .ZN(G1342gat));
  NOR2_X1   g623(.A1(new_n816), .A2(new_n655), .ZN(new_n825));
  NOR2_X1   g624(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n826));
  AND2_X1   g625(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n828), .B1(new_n825), .B2(new_n826), .ZN(G1343gat));
  AND2_X1   g628(.A1(new_n641), .A2(new_n815), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n813), .A2(new_n644), .A3(new_n830), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n831), .A2(G141gat), .A3(new_n513), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n832), .A2(KEYINPUT58), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT57), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n813), .A2(new_n834), .A3(new_n644), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n789), .A2(new_n512), .A3(new_n617), .A4(new_n790), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n591), .B1(new_n801), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n808), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n811), .B1(new_n839), .B2(new_n569), .ZN(new_n840));
  OAI21_X1  g639(.A(KEYINPUT57), .B1(new_n840), .B2(new_n379), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n835), .A2(new_n830), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(G141gat), .B1(new_n842), .B2(new_n513), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n833), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n835), .A2(new_n668), .A3(new_n830), .A4(new_n841), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n845), .A2(KEYINPUT120), .A3(G141gat), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT120), .B1(new_n845), .B2(G141gat), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n846), .A2(new_n847), .A3(new_n832), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT58), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n844), .B1(new_n848), .B2(new_n849), .ZN(G1344gat));
  INV_X1    g649(.A(new_n831), .ZN(new_n851));
  INV_X1    g650(.A(G148gat), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n852), .A3(new_n624), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n854), .B1(new_n842), .B2(new_n692), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n852), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n655), .A2(new_n791), .A3(new_n799), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n569), .B1(new_n837), .B2(new_n857), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n568), .A2(new_n513), .A3(new_n655), .A4(new_n692), .ZN(new_n859));
  AOI211_X1 g658(.A(KEYINPUT57), .B(new_n379), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n568), .B1(new_n806), .B2(new_n808), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n644), .B1(new_n861), .B2(new_n811), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n860), .B1(new_n862), .B2(KEYINPUT57), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(new_n624), .A3(new_n830), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n854), .B1(new_n864), .B2(G148gat), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n853), .B1(new_n856), .B2(new_n865), .ZN(G1345gat));
  OAI21_X1  g665(.A(G155gat), .B1(new_n842), .B2(new_n569), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n851), .A2(new_n222), .A3(new_n568), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(G1346gat));
  OAI21_X1  g668(.A(G162gat), .B1(new_n842), .B2(new_n655), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n851), .A2(new_n223), .A3(new_n591), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1347gat));
  AOI21_X1  g671(.A(new_n448), .B1(new_n810), .B2(new_n812), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(new_n385), .A3(new_n718), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n274), .A3(new_n668), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(KEYINPUT121), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n875), .A2(new_n512), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n879), .B2(G169gat), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n877), .B1(new_n876), .B2(new_n880), .ZN(G1348gat));
  NOR2_X1   g680(.A1(new_n874), .A2(new_n692), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n316), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n883), .B1(new_n275), .B2(new_n882), .ZN(G1349gat));
  NAND3_X1  g683(.A1(new_n875), .A2(new_n308), .A3(new_n568), .ZN(new_n885));
  OAI21_X1  g684(.A(G183gat), .B1(new_n874), .B2(new_n569), .ZN(new_n886));
  XOR2_X1   g685(.A(KEYINPUT122), .B(KEYINPUT60), .Z(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n885), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT60), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n890), .B1(new_n885), .B2(new_n886), .ZN(new_n891));
  OAI21_X1  g690(.A(KEYINPUT123), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n885), .A2(new_n886), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n894), .B2(new_n887), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n892), .A2(new_n895), .ZN(G1350gat));
  NAND3_X1  g695(.A1(new_n875), .A2(new_n291), .A3(new_n591), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT124), .ZN(new_n898));
  OAI21_X1  g697(.A(G190gat), .B1(new_n874), .B2(new_n655), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT61), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(new_n900), .ZN(G1351gat));
  INV_X1    g700(.A(G197gat), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT126), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n862), .A2(KEYINPUT57), .ZN(new_n904));
  INV_X1    g703(.A(new_n860), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI211_X1 g705(.A(KEYINPUT126), .B(new_n860), .C1(new_n862), .C2(KEYINPUT57), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n437), .A2(new_n445), .A3(new_n438), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n439), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n902), .B1(new_n910), .B2(new_n512), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n908), .A2(new_n644), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n873), .B1(KEYINPUT125), .B2(new_n912), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n912), .A2(KEYINPUT125), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(new_n902), .A3(new_n668), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT127), .B1(new_n911), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n904), .A2(new_n905), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT126), .ZN(new_n920));
  INV_X1    g719(.A(new_n909), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n863), .A2(new_n903), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(G197gat), .B1(new_n923), .B2(new_n513), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT127), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n924), .A2(new_n925), .A3(new_n916), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n918), .A2(new_n926), .ZN(G1352gat));
  NOR4_X1   g726(.A1(new_n913), .A2(G204gat), .A3(new_n692), .A4(new_n914), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT62), .ZN(new_n929));
  OAI21_X1  g728(.A(G204gat), .B1(new_n923), .B2(new_n692), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1353gat));
  NAND3_X1  g730(.A1(new_n915), .A2(new_n322), .A3(new_n568), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n863), .A2(new_n568), .A3(new_n921), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n933), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n934));
  AOI21_X1  g733(.A(KEYINPUT63), .B1(new_n933), .B2(G211gat), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(G1354gat));
  AOI21_X1  g735(.A(G218gat), .B1(new_n915), .B2(new_n591), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n655), .A2(new_n323), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n937), .B1(new_n910), .B2(new_n938), .ZN(G1355gat));
endmodule


