//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0 1 1 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n597, new_n598, new_n599, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n649, new_n650, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1214,
    new_n1215, new_n1216, new_n1217;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G221), .A3(G219), .A4(G218), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT68), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n454), .ZN(new_n461));
  AOI22_X1  g036(.A1(new_n458), .A2(new_n459), .B1(G567), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n468), .A2(KEYINPUT69), .ZN(new_n476));
  NOR3_X1   g051(.A1(new_n475), .A2(new_n476), .A3(G2105), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n477), .A2(new_n478), .A3(G101), .ZN(new_n479));
  XNOR2_X1  g054(.A(KEYINPUT69), .B(G2104), .ZN(new_n480));
  INV_X1    g055(.A(G2105), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n480), .A2(G101), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT70), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n473), .A2(new_n479), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g059(.A(KEYINPUT3), .B1(new_n475), .B2(new_n476), .ZN(new_n485));
  AND4_X1   g060(.A1(G137), .A2(new_n485), .A3(new_n481), .A4(new_n467), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n484), .A2(new_n486), .ZN(G160));
  NAND2_X1  g062(.A1(new_n468), .A2(KEYINPUT69), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n474), .A2(G2104), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n466), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n491));
  NOR3_X1   g066(.A1(new_n490), .A2(G2105), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G136), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT72), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n494), .A2(G100), .A3(G2105), .ZN(new_n495));
  OR2_X1    g070(.A1(new_n481), .A2(G112), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n494), .B1(G100), .B2(G2105), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n496), .A2(G2104), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n493), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n500));
  OAI211_X1 g075(.A(G2105), .B(new_n467), .C1(new_n480), .C2(new_n466), .ZN(new_n501));
  INV_X1    g076(.A(G124), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  NOR3_X1   g079(.A1(new_n501), .A2(new_n500), .A3(new_n502), .ZN(new_n505));
  OR3_X1    g080(.A1(new_n499), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G162));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(new_n481), .A3(G138), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n470), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G138), .ZN(new_n512));
  NOR4_X1   g087(.A1(new_n490), .A2(new_n512), .A3(G2105), .A4(new_n491), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n511), .B1(new_n513), .B2(new_n508), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n481), .A2(G114), .ZN(new_n516));
  OAI21_X1  g091(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NOR3_X1   g093(.A1(new_n490), .A2(new_n481), .A3(new_n491), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n518), .B1(new_n519), .B2(G126), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n514), .A2(new_n515), .A3(new_n520), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n485), .A2(G138), .A3(new_n481), .A4(new_n467), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n510), .B1(new_n522), .B2(KEYINPUT4), .ZN(new_n523));
  INV_X1    g098(.A(G126), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n501), .A2(new_n524), .B1(new_n516), .B2(new_n517), .ZN(new_n525));
  OAI21_X1  g100(.A(KEYINPUT73), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n521), .A2(new_n526), .ZN(G164));
  XOR2_X1   g102(.A(KEYINPUT74), .B(G651), .Z(new_n528));
  INV_X1    g103(.A(KEYINPUT5), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(G543), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G543), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n529), .A2(KEYINPUT76), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT5), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n532), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT77), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n531), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n534), .A2(KEYINPUT5), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n529), .A2(KEYINPUT76), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n537), .B(G543), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G62), .ZN(new_n544));
  NAND2_X1  g119(.A1(G75), .A2(G543), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n528), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  XNOR2_X1  g121(.A(KEYINPUT76), .B(KEYINPUT5), .ZN(new_n547));
  OAI21_X1  g122(.A(KEYINPUT77), .B1(new_n547), .B2(new_n532), .ZN(new_n548));
  NAND2_X1  g123(.A1(KEYINPUT75), .A2(G651), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(KEYINPUT6), .ZN(new_n550));
  OAI21_X1  g125(.A(KEYINPUT6), .B1(KEYINPUT74), .B2(G651), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g127(.A1(KEYINPUT74), .A2(KEYINPUT75), .A3(G651), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n548), .A2(new_n554), .A3(new_n541), .A4(new_n531), .ZN(new_n555));
  INV_X1    g130(.A(G88), .ZN(new_n556));
  INV_X1    g131(.A(G50), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(G543), .ZN(new_n558));
  OAI22_X1  g133(.A1(new_n555), .A2(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n546), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT78), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT78), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n562), .B1(new_n546), .B2(new_n559), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(G166));
  NAND3_X1  g139(.A1(new_n543), .A2(G63), .A3(G651), .ZN(new_n565));
  NAND3_X1  g140(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n566));
  XOR2_X1   g141(.A(new_n566), .B(KEYINPUT7), .Z(new_n567));
  INV_X1    g142(.A(new_n558), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n567), .B1(new_n568), .B2(G51), .ZN(new_n569));
  INV_X1    g144(.A(G89), .ZN(new_n570));
  OAI211_X1 g145(.A(new_n565), .B(new_n569), .C1(new_n570), .C2(new_n555), .ZN(G286));
  INV_X1    g146(.A(G286), .ZN(G168));
  NAND2_X1  g147(.A1(G77), .A2(G543), .ZN(new_n573));
  OAI21_X1  g148(.A(G543), .B1(new_n539), .B2(new_n540), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n530), .B1(new_n574), .B2(KEYINPUT77), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(new_n541), .ZN(new_n576));
  INV_X1    g151(.A(G64), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n573), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n528), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT79), .ZN(new_n581));
  INV_X1    g156(.A(new_n555), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G90), .B1(G52), .B2(new_n568), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n580), .A2(KEYINPUT79), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n584), .A2(new_n585), .ZN(G171));
  NAND2_X1  g161(.A1(G68), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G56), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n576), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(new_n579), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n582), .A2(G81), .B1(G43), .B2(new_n568), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G860), .ZN(G153));
  AND3_X1   g169(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G36), .ZN(G176));
  NAND2_X1  g171(.A1(G1), .A2(G3), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT80), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT8), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(G188));
  OAI21_X1  g175(.A(KEYINPUT83), .B1(new_n538), .B2(new_n542), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT83), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n575), .A2(new_n602), .A3(new_n541), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n601), .A2(new_n603), .A3(G65), .ZN(new_n604));
  NAND2_X1  g179(.A1(G78), .A2(G543), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G651), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT82), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n555), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n575), .A2(KEYINPUT82), .A3(new_n541), .A4(new_n554), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(KEYINPUT81), .A2(G53), .ZN(new_n612));
  OR3_X1    g187(.A1(new_n558), .A2(KEYINPUT9), .A3(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(KEYINPUT9), .B1(new_n558), .B2(new_n612), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n611), .A2(G91), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n607), .A2(new_n615), .ZN(G299));
  INV_X1    g191(.A(G171), .ZN(G301));
  INV_X1    g192(.A(G166), .ZN(G303));
  INV_X1    g193(.A(G651), .ZN(new_n619));
  INV_X1    g194(.A(G74), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n619), .B1(new_n576), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(G49), .B2(new_n568), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n611), .A2(G87), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(G288));
  NAND3_X1  g199(.A1(new_n575), .A2(G61), .A3(new_n541), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT84), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n625), .A2(new_n626), .B1(G73), .B2(G543), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n543), .A2(KEYINPUT84), .A3(G61), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n528), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AND2_X1   g204(.A1(new_n568), .A2(G48), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n611), .A2(G86), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(new_n632), .ZN(G305));
  AOI22_X1  g208(.A1(new_n543), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n634), .A2(new_n528), .ZN(new_n635));
  AOI22_X1  g210(.A1(new_n582), .A2(G85), .B1(G47), .B2(new_n568), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(G290));
  NAND3_X1  g212(.A1(new_n601), .A2(new_n603), .A3(G66), .ZN(new_n638));
  INV_X1    g213(.A(G79), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n638), .B1(new_n639), .B2(new_n532), .ZN(new_n640));
  AOI22_X1  g215(.A1(new_n640), .A2(G651), .B1(G54), .B2(new_n568), .ZN(new_n641));
  AOI21_X1  g216(.A(KEYINPUT10), .B1(new_n611), .B2(G92), .ZN(new_n642));
  AND3_X1   g217(.A1(new_n611), .A2(KEYINPUT10), .A3(G92), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(G868), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(G171), .ZN(G284));
  OAI21_X1  g222(.A(new_n646), .B1(new_n645), .B2(G171), .ZN(G321));
  NAND2_X1  g223(.A1(G286), .A2(G868), .ZN(new_n649));
  XNOR2_X1  g224(.A(G299), .B(KEYINPUT85), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n649), .B1(new_n650), .B2(G868), .ZN(G297));
  OAI21_X1  g226(.A(new_n649), .B1(new_n650), .B2(G868), .ZN(G280));
  INV_X1    g227(.A(new_n644), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT86), .B(G559), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n653), .B1(G860), .B2(new_n654), .ZN(G148));
  NAND2_X1  g230(.A1(new_n592), .A2(new_n645), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n653), .A2(new_n654), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(KEYINPUT87), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT87), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n653), .A2(new_n659), .A3(new_n654), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n656), .B1(new_n662), .B2(new_n645), .ZN(G323));
  XNOR2_X1  g238(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g239(.A1(new_n492), .A2(G135), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n481), .A2(G111), .ZN(new_n666));
  OAI21_X1  g241(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(G123), .B2(new_n519), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT89), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(G2096), .Z(new_n671));
  NAND3_X1  g246(.A1(new_n477), .A2(new_n467), .A3(new_n469), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT12), .Z(new_n673));
  INV_X1    g248(.A(G2100), .ZN(new_n674));
  OAI22_X1  g249(.A1(new_n673), .A2(KEYINPUT13), .B1(KEYINPUT88), .B2(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(KEYINPUT13), .B2(new_n673), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(KEYINPUT88), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n671), .A2(new_n678), .ZN(G156));
  XOR2_X1   g254(.A(KEYINPUT15), .B(G2435), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G2438), .ZN(new_n681));
  XOR2_X1   g256(.A(G2427), .B(G2430), .Z(new_n682));
  OAI21_X1  g257(.A(KEYINPUT14), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT90), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n682), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G2451), .B(G2454), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT16), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G2443), .B(G2446), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1341), .B(G1348), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g269(.A(G14), .B1(new_n691), .B2(new_n693), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(G401));
  XOR2_X1   g271(.A(G2084), .B(G2090), .Z(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G2067), .B(G2678), .Z(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(G2072), .B(G2078), .Z(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n700), .A2(KEYINPUT17), .A3(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n698), .A2(new_n699), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n700), .A2(KEYINPUT17), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n703), .B(new_n705), .C1(new_n706), .C2(new_n702), .ZN(new_n707));
  OR3_X1    g282(.A1(new_n705), .A2(KEYINPUT18), .A3(new_n701), .ZN(new_n708));
  OAI21_X1  g283(.A(KEYINPUT18), .B1(new_n705), .B2(new_n701), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(new_n674), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT91), .B(G2096), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(G227));
  XNOR2_X1  g288(.A(G1971), .B(G1976), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT19), .ZN(new_n715));
  XOR2_X1   g290(.A(G1956), .B(G2474), .Z(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  XOR2_X1   g292(.A(G1961), .B(G1966), .Z(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  NOR3_X1   g294(.A1(new_n715), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT92), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n721), .A2(KEYINPUT20), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(KEYINPUT20), .ZN(new_n723));
  NOR3_X1   g298(.A1(new_n715), .A2(new_n716), .A3(new_n718), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n716), .B(new_n718), .Z(new_n725));
  AOI21_X1  g300(.A(new_n724), .B1(new_n715), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n722), .A2(new_n723), .A3(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(G1991), .B(G1996), .Z(new_n728));
  XNOR2_X1  g303(.A(G1981), .B(G1986), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT93), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n730), .B(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n727), .B(new_n733), .ZN(G229));
  NOR2_X1   g309(.A1(G16), .A2(G22), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G166), .B2(G16), .ZN(new_n736));
  INV_X1    g311(.A(G1971), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G6), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(G16), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G305), .B2(G16), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT32), .B(G1981), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G16), .A2(G23), .ZN(new_n744));
  INV_X1    g319(.A(G288), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(G16), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT33), .B(G1976), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n738), .A2(new_n743), .A3(new_n748), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT34), .Z(new_n750));
  MUX2_X1   g325(.A(G24), .B(G290), .S(G16), .Z(new_n751));
  OR2_X1    g326(.A1(new_n751), .A2(G1986), .ZN(new_n752));
  INV_X1    g327(.A(G29), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(G25), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n519), .A2(G119), .ZN(new_n755));
  OR2_X1    g330(.A1(G95), .A2(G2105), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n756), .B(G2104), .C1(G107), .C2(new_n481), .ZN(new_n757));
  INV_X1    g332(.A(new_n492), .ZN(new_n758));
  INV_X1    g333(.A(G131), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n755), .B(new_n757), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n754), .B1(new_n761), .B2(new_n753), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT35), .B(G1991), .Z(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n752), .A2(KEYINPUT94), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G1986), .B2(new_n751), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n750), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(KEYINPUT36), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT36), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n750), .A2(new_n769), .A3(new_n766), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n753), .A2(G35), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G162), .B2(new_n753), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT29), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n774), .A2(G2090), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n753), .A2(G27), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G164), .B2(new_n753), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n775), .B1(G2078), .B2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT98), .ZN(new_n779));
  NOR2_X1   g354(.A1(G5), .A2(G16), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G171), .B2(G16), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G1961), .ZN(new_n782));
  OAI221_X1 g357(.A(new_n778), .B1(G2078), .B2(new_n777), .C1(new_n779), .C2(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n779), .B2(new_n782), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n753), .A2(G33), .ZN(new_n785));
  NAND2_X1  g360(.A1(G115), .A2(G2104), .ZN(new_n786));
  INV_X1    g361(.A(G127), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n470), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(G2105), .B1(new_n788), .B2(KEYINPUT96), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(KEYINPUT96), .B2(new_n788), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n481), .A2(G103), .A3(G2104), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT25), .Z(new_n792));
  INV_X1    g367(.A(G139), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n792), .B1(new_n758), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n790), .A2(new_n794), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT97), .Z(new_n796));
  OAI21_X1  g371(.A(new_n785), .B1(new_n796), .B2(new_n753), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(G2072), .Z(new_n798));
  INV_X1    g373(.A(G28), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n799), .A2(KEYINPUT30), .ZN(new_n800));
  AOI21_X1  g375(.A(G29), .B1(new_n799), .B2(KEYINPUT30), .ZN(new_n801));
  OR2_X1    g376(.A1(KEYINPUT31), .A2(G11), .ZN(new_n802));
  NAND2_X1  g377(.A1(KEYINPUT31), .A2(G11), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n800), .A2(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n670), .B2(new_n753), .ZN(new_n805));
  NOR2_X1   g380(.A1(G16), .A2(G21), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G168), .B2(G16), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n807), .A2(G1966), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n807), .A2(G1966), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n805), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  AND2_X1   g385(.A1(KEYINPUT24), .A2(G34), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n753), .B1(KEYINPUT24), .B2(G34), .ZN(new_n812));
  OAI22_X1  g387(.A1(G160), .A2(new_n753), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(G2084), .ZN(new_n814));
  NOR2_X1   g389(.A1(G29), .A2(G32), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n492), .A2(G141), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n519), .A2(G129), .ZN(new_n817));
  NAND3_X1  g392(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT26), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n477), .A2(G105), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n816), .A2(new_n817), .A3(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n815), .B1(new_n824), .B2(G29), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT27), .B(G1996), .Z(new_n826));
  OAI21_X1  g401(.A(new_n814), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G2084), .B2(new_n813), .ZN(new_n829));
  INV_X1    g404(.A(G2067), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n753), .A2(G26), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n519), .A2(G128), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n492), .A2(G140), .ZN(new_n833));
  NOR3_X1   g408(.A1(KEYINPUT95), .A2(G104), .A3(G2105), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n481), .A2(G116), .ZN(new_n835));
  OAI21_X1  g410(.A(KEYINPUT95), .B1(G104), .B2(G2105), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n835), .A2(G2104), .A3(new_n836), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n832), .B(new_n833), .C1(new_n834), .C2(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n831), .B1(new_n838), .B2(G29), .ZN(new_n839));
  MUX2_X1   g414(.A(new_n831), .B(new_n839), .S(KEYINPUT28), .Z(new_n840));
  AOI211_X1 g415(.A(new_n827), .B(new_n829), .C1(new_n830), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n774), .A2(G2090), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n798), .A2(new_n810), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT23), .ZN(new_n844));
  INV_X1    g419(.A(G20), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n845), .A2(G16), .ZN(new_n846));
  AOI211_X1 g421(.A(new_n844), .B(new_n846), .C1(G299), .C2(G16), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(new_n844), .B2(new_n846), .ZN(new_n848));
  XNOR2_X1  g423(.A(KEYINPUT99), .B(G1956), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n848), .B(new_n849), .Z(new_n850));
  INV_X1    g425(.A(G4), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n851), .A2(G16), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(new_n644), .B2(G16), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(G1348), .Z(new_n854));
  INV_X1    g429(.A(new_n840), .ZN(new_n855));
  INV_X1    g430(.A(G1341), .ZN(new_n856));
  INV_X1    g431(.A(G19), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n857), .A2(G16), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n858), .B1(new_n592), .B2(G16), .ZN(new_n859));
  AOI22_X1  g434(.A1(new_n855), .A2(G2067), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  OAI221_X1 g435(.A(new_n860), .B1(new_n856), .B2(new_n859), .C1(new_n781), .C2(G1961), .ZN(new_n861));
  NOR4_X1   g436(.A1(new_n843), .A2(new_n850), .A3(new_n854), .A4(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n771), .A2(new_n784), .A3(new_n862), .ZN(G150));
  INV_X1    g438(.A(G150), .ZN(G311));
  INV_X1    g439(.A(G93), .ZN(new_n865));
  INV_X1    g440(.A(G55), .ZN(new_n866));
  OAI22_X1  g441(.A1(new_n555), .A2(new_n865), .B1(new_n866), .B2(new_n558), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n543), .A2(G67), .ZN(new_n868));
  NAND2_X1  g443(.A1(G80), .A2(G543), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n867), .B1(new_n870), .B2(new_n579), .ZN(new_n871));
  INV_X1    g446(.A(G860), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT37), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n653), .A2(G559), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT38), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n592), .A2(new_n871), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n528), .B1(new_n868), .B2(new_n869), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n591), .B(new_n590), .C1(new_n878), .C2(new_n867), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n876), .B(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT39), .ZN(new_n883));
  OR3_X1    g458(.A1(new_n882), .A2(KEYINPUT101), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(KEYINPUT101), .B1(new_n882), .B2(new_n883), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n883), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n884), .B(new_n885), .C1(KEYINPUT100), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(KEYINPUT100), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(new_n872), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n874), .B1(new_n887), .B2(new_n889), .ZN(G145));
  NAND2_X1  g465(.A1(new_n514), .A2(new_n520), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n838), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n796), .B(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(new_n823), .ZN(new_n894));
  OAI21_X1  g469(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n895));
  INV_X1    g470(.A(G118), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n895), .B1(new_n896), .B2(G2105), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n897), .B1(new_n492), .B2(G142), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n519), .A2(KEYINPUT102), .A3(G130), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT102), .ZN(new_n900));
  INV_X1    g475(.A(G130), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n900), .B1(new_n501), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n898), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(new_n760), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT103), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n905), .B(new_n673), .Z(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n908));
  OR3_X1    g483(.A1(new_n894), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n894), .B1(new_n907), .B2(new_n908), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n670), .B(new_n506), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(G160), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n909), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n894), .B2(new_n906), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n894), .A2(new_n906), .ZN(new_n915));
  AOI21_X1  g490(.A(G37), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g493(.A1(new_n662), .A2(new_n880), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n661), .A2(new_n881), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G299), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n644), .A2(new_n922), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n643), .A2(new_n642), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n924), .A2(G299), .A3(new_n641), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n921), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT41), .ZN(new_n928));
  INV_X1    g503(.A(new_n925), .ZN(new_n929));
  AOI21_X1  g504(.A(G299), .B1(new_n924), .B2(new_n641), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n923), .A2(new_n925), .A3(KEYINPUT41), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n919), .A2(new_n933), .A3(new_n920), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n927), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(G303), .A2(G305), .ZN(new_n936));
  NAND3_X1  g511(.A1(G166), .A2(new_n632), .A3(new_n631), .ZN(new_n937));
  XNOR2_X1  g512(.A(G290), .B(G288), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n938), .B1(new_n936), .B2(new_n937), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT42), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT105), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT105), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT42), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n942), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n941), .A2(KEYINPUT105), .A3(new_n943), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT106), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n935), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n927), .A2(new_n947), .A3(new_n934), .A4(new_n948), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n950), .B1(new_n935), .B2(new_n949), .ZN(new_n954));
  OAI21_X1  g529(.A(G868), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n645), .B1(new_n878), .B2(new_n867), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(G295));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n956), .ZN(G331));
  NAND3_X1  g533(.A1(new_n877), .A2(new_n879), .A3(G286), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(G286), .B1(new_n877), .B2(new_n879), .ZN(new_n961));
  OAI21_X1  g536(.A(G301), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n880), .A2(G168), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n963), .A2(G171), .A3(new_n959), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n962), .A2(new_n926), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n931), .A2(new_n967), .A3(new_n932), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n962), .A2(new_n964), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n926), .A2(KEYINPUT108), .A3(new_n928), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n966), .B1(new_n971), .B2(KEYINPUT109), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n968), .A2(new_n973), .A3(new_n969), .A4(new_n970), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n942), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT43), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n933), .A2(new_n969), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n965), .A2(KEYINPUT107), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT107), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n962), .A2(new_n926), .A3(new_n964), .A4(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n979), .A2(new_n941), .A3(new_n980), .A4(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G37), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n976), .A2(new_n977), .A3(new_n978), .A4(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n941), .B1(new_n972), .B2(new_n974), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n989), .A2(KEYINPUT43), .A3(new_n985), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n933), .A2(new_n969), .B1(new_n965), .B2(KEYINPUT107), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n941), .B1(new_n991), .B2(new_n982), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT43), .B1(new_n985), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT110), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n987), .B(new_n988), .C1(new_n990), .C2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n985), .A2(new_n992), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n988), .B1(new_n996), .B2(new_n978), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT43), .B1(new_n989), .B2(new_n985), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n997), .A2(new_n998), .A3(KEYINPUT111), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT111), .B1(new_n997), .B2(new_n998), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n995), .B1(new_n999), .B2(new_n1000), .ZN(G397));
  INV_X1    g576(.A(KEYINPUT57), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n611), .A2(G91), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n613), .A2(new_n614), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n619), .B1(new_n604), .B2(new_n605), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1002), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n607), .A2(KEYINPUT57), .A3(new_n615), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n1010));
  INV_X1    g585(.A(G1384), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n521), .A2(new_n526), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n472), .A2(G2105), .B1(new_n482), .B2(KEYINPUT70), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n492), .A2(G137), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1013), .A2(new_n1014), .A3(G40), .A4(new_n479), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1011), .B1(new_n523), .B2(new_n525), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1015), .B1(new_n1016), .B2(KEYINPUT50), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1012), .A2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g593(.A(KEYINPUT121), .B(G1956), .Z(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g595(.A(KEYINPUT45), .B(new_n1011), .C1(new_n523), .C2(new_n525), .ZN(new_n1021));
  INV_X1    g596(.A(G40), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n484), .A2(new_n1022), .A3(new_n486), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n521), .A2(new_n526), .A3(new_n1011), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1024), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g602(.A(KEYINPUT56), .B(G2072), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n1028), .B(KEYINPUT122), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1009), .B1(new_n1020), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1023), .B1(new_n1016), .B2(KEYINPUT50), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1032), .B1(KEYINPUT50), .B2(new_n1025), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1016), .A2(new_n1015), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  OAI22_X1  g610(.A1(new_n1033), .A2(G1348), .B1(G2067), .B2(new_n1035), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1036), .A2(new_n653), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n1027), .A2(new_n1029), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n1009), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1031), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n1036), .A2(KEYINPUT60), .A3(new_n644), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1036), .B(new_n653), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1041), .B1(new_n1042), .B2(KEYINPUT60), .ZN(new_n1043));
  XOR2_X1   g618(.A(KEYINPUT58), .B(G1341), .Z(new_n1044));
  NAND2_X1  g619(.A1(new_n1035), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1046), .A2(new_n1023), .A3(new_n1021), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1045), .B1(new_n1047), .B2(G1996), .ZN(new_n1048));
  XNOR2_X1  g623(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(new_n593), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n1051));
  INV_X1    g626(.A(G1996), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1027), .A2(new_n1052), .B1(new_n1035), .B2(new_n1044), .ZN(new_n1053));
  OAI211_X1 g628(.A(KEYINPUT123), .B(new_n1051), .C1(new_n1053), .C2(new_n592), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1050), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT124), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(new_n1038), .B2(new_n1009), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1009), .A2(new_n1030), .A3(new_n1020), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1057), .B(KEYINPUT61), .C1(new_n1058), .C2(new_n1031), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1030), .A2(new_n1020), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1009), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT61), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1062), .B(new_n1039), .C1(new_n1056), .C2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1055), .B1(new_n1059), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT125), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1043), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  AOI211_X1 g642(.A(KEYINPUT125), .B(new_n1055), .C1(new_n1059), .C2(new_n1064), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1040), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT49), .ZN(new_n1070));
  INV_X1    g645(.A(G86), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n555), .A2(new_n1071), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n629), .A2(new_n630), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1981), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n632), .ZN(new_n1076));
  NOR4_X1   g651(.A1(new_n629), .A2(new_n1076), .A3(G1981), .A4(new_n630), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1070), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n631), .A2(new_n1074), .A3(new_n632), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1079), .B(KEYINPUT49), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1080));
  INV_X1    g655(.A(G8), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1034), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1078), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G1976), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT52), .B1(G288), .B2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1085), .B(new_n1082), .C1(new_n1084), .C2(G288), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1082), .B1(G288), .B2(new_n1084), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT52), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1083), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT55), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1091), .B1(G166), .B2(new_n1081), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n561), .A2(KEYINPUT55), .A3(G8), .A4(new_n563), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1047), .A2(new_n737), .ZN(new_n1095));
  INV_X1    g670(.A(G2090), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1033), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1081), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT115), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1094), .A2(new_n1098), .A3(KEYINPUT115), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1090), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(G2090), .B1(new_n1018), .B2(KEYINPUT116), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(KEYINPUT116), .B2(new_n1018), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(new_n1106), .A3(new_n1095), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(G8), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1106), .B1(new_n1105), .B2(new_n1095), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1092), .B(new_n1093), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1103), .A2(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(G171), .B(KEYINPUT54), .ZN(new_n1112));
  INV_X1    g687(.A(G2078), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT53), .B1(new_n1027), .B2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1033), .A2(G1961), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1113), .A2(KEYINPUT53), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT127), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1118), .B1(new_n1023), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1016), .A2(new_n1026), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1015), .A2(KEYINPUT127), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1120), .A2(new_n1121), .A3(new_n1021), .A4(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1112), .A2(new_n1116), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT118), .ZN(new_n1125));
  AOI21_X1  g700(.A(G1384), .B1(new_n514), .B2(new_n520), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1125), .B1(new_n1126), .B2(KEYINPUT45), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n521), .A2(new_n526), .A3(KEYINPUT45), .A4(new_n1011), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1023), .B1(new_n1128), .B2(KEYINPUT118), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1129), .A2(new_n1130), .A3(new_n1118), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1131), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1124), .B1(new_n1132), .B2(new_n1112), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1111), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(G1966), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1135), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT119), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT119), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1138), .B(new_n1135), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1139));
  AOI211_X1 g714(.A(G2084), .B(new_n1032), .C1(KEYINPUT50), .C2(new_n1025), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1137), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(G168), .A2(new_n1081), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1140), .B1(new_n1136), .B2(KEYINPUT119), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1081), .B1(new_n1145), .B2(new_n1139), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT51), .B1(new_n1146), .B2(KEYINPUT126), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1146), .A2(new_n1143), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI221_X4 g724(.A(new_n1143), .B1(KEYINPUT126), .B2(KEYINPUT51), .C1(new_n1142), .C2(G8), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1144), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1069), .A2(new_n1134), .A3(new_n1151), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1083), .A2(new_n1084), .A3(new_n745), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1082), .B1(new_n1153), .B2(new_n1077), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1154), .B1(new_n1155), .B2(new_n1090), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1142), .A2(G8), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1157), .A2(G286), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1103), .A2(new_n1110), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT63), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1162));
  OR3_X1    g737(.A1(new_n1090), .A2(KEYINPUT120), .A3(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(KEYINPUT120), .B1(new_n1090), .B2(new_n1162), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1160), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1163), .A2(new_n1158), .A3(new_n1164), .A4(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1156), .B1(new_n1161), .B2(new_n1166), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n1132), .A2(G301), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1111), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1144), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1157), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1143), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1157), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1172), .A2(new_n1174), .A3(KEYINPUT51), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1170), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1169), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  AOI211_X1 g754(.A(KEYINPUT62), .B(new_n1170), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1152), .B(new_n1167), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1121), .A2(new_n1015), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(new_n1052), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1183), .A2(new_n823), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1182), .B(KEYINPUT113), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n838), .B(new_n830), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT114), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1184), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1185), .A2(G1996), .A3(new_n823), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n760), .B(new_n763), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1185), .ZN(new_n1191));
  OAI211_X1 g766(.A(new_n1188), .B(new_n1189), .C1(new_n1190), .C2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(G290), .ZN(new_n1193));
  INV_X1    g768(.A(G1986), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  XOR2_X1   g770(.A(new_n1195), .B(KEYINPUT112), .Z(new_n1196));
  INV_X1    g771(.A(new_n1196), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1197), .B1(new_n1194), .B2(new_n1193), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1192), .B1(new_n1198), .B2(new_n1182), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1181), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1196), .A2(new_n1182), .ZN(new_n1201));
  XOR2_X1   g776(.A(new_n1201), .B(KEYINPUT48), .Z(new_n1202));
  NOR2_X1   g777(.A1(new_n1202), .A2(new_n1192), .ZN(new_n1203));
  NAND4_X1  g778(.A1(new_n1188), .A2(new_n763), .A3(new_n1189), .A4(new_n761), .ZN(new_n1204));
  OR2_X1    g779(.A1(new_n838), .A2(G2067), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1191), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g781(.A(new_n1183), .B(KEYINPUT46), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1207), .B1(new_n1191), .B2(new_n824), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1208), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n1209), .B(KEYINPUT47), .ZN(new_n1210));
  NOR3_X1   g785(.A1(new_n1203), .A2(new_n1206), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1200), .A2(new_n1211), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g787(.A1(new_n976), .A2(new_n978), .A3(new_n986), .ZN(new_n1214));
  NAND3_X1  g788(.A1(new_n1214), .A2(KEYINPUT110), .A3(new_n993), .ZN(new_n1215));
  NOR4_X1   g789(.A1(G401), .A2(new_n463), .A3(G227), .A4(G229), .ZN(new_n1216));
  AND2_X1   g790(.A1(new_n917), .A2(new_n1216), .ZN(new_n1217));
  AND3_X1   g791(.A1(new_n1215), .A2(new_n1217), .A3(new_n987), .ZN(G308));
  NAND3_X1  g792(.A1(new_n1215), .A2(new_n1217), .A3(new_n987), .ZN(G225));
endmodule


