

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741;

  NAND2_X1 U377 ( .A1(n379), .A2(n606), .ZN(n610) );
  OR2_X1 U378 ( .A1(n632), .A2(n631), .ZN(n628) );
  XNOR2_X1 U379 ( .A(n563), .B(KEYINPUT1), .ZN(n523) );
  XNOR2_X1 U380 ( .A(KEYINPUT90), .B(G110), .ZN(n409) );
  XNOR2_X1 U381 ( .A(n417), .B(G125), .ZN(n449) );
  XNOR2_X1 U382 ( .A(n414), .B(G143), .ZN(n465) );
  INV_X2 U383 ( .A(G953), .ZN(n469) );
  AND2_X1 U384 ( .A1(n368), .A2(n367), .ZN(n665) );
  AND2_X1 U385 ( .A1(n370), .A2(n367), .ZN(n687) );
  XNOR2_X1 U386 ( .A(n528), .B(KEYINPUT35), .ZN(n682) );
  NAND2_X2 U387 ( .A1(n375), .A2(n372), .ZN(n381) );
  AND2_X2 U388 ( .A1(n543), .A2(n355), .ZN(n375) );
  AND2_X2 U389 ( .A1(n369), .A2(n367), .ZN(n693) );
  XNOR2_X2 U390 ( .A(G128), .B(KEYINPUT80), .ZN(n414) );
  NAND2_X2 U391 ( .A1(n390), .A2(n388), .ZN(n563) );
  XNOR2_X2 U392 ( .A(n483), .B(KEYINPUT22), .ZN(n541) );
  AND2_X2 U393 ( .A1(n669), .A2(n380), .ZN(n655) );
  NAND2_X1 U394 ( .A1(n374), .A2(n373), .ZN(n372) );
  NAND2_X1 U395 ( .A1(n357), .A2(n522), .ZN(n374) );
  OR2_X1 U396 ( .A1(n682), .A2(KEYINPUT44), .ZN(n357) );
  INV_X1 U397 ( .A(KEYINPUT71), .ZN(n387) );
  XNOR2_X1 U398 ( .A(n371), .B(n360), .ZN(n683) );
  NOR2_X1 U399 ( .A1(n597), .A2(n578), .ZN(n558) );
  XNOR2_X1 U400 ( .A(n545), .B(n386), .ZN(n580) );
  XNOR2_X1 U401 ( .A(n387), .B(G131), .ZN(n485) );
  NAND2_X1 U402 ( .A1(n411), .A2(n632), .ZN(n681) );
  XNOR2_X1 U403 ( .A(n412), .B(KEYINPUT67), .ZN(n411) );
  NAND2_X1 U404 ( .A1(n504), .A2(n503), .ZN(n412) );
  OR2_X1 U405 ( .A1(n580), .A2(n559), .ZN(n518) );
  NAND2_X1 U406 ( .A1(n592), .A2(n591), .ZN(n398) );
  NAND2_X1 U407 ( .A1(n681), .A2(n683), .ZN(n544) );
  INV_X1 U408 ( .A(G146), .ZN(n417) );
  XNOR2_X1 U409 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U410 ( .A(KEYINPUT103), .B(KEYINPUT12), .ZN(n451) );
  XOR2_X1 U411 ( .A(G122), .B(G104), .Z(n457) );
  XNOR2_X1 U412 ( .A(n730), .B(n487), .ZN(n502) );
  INV_X1 U413 ( .A(G146), .ZN(n487) );
  XNOR2_X1 U414 ( .A(n401), .B(n400), .ZN(n399) );
  NOR2_X1 U415 ( .A1(n523), .A2(n628), .ZN(n529) );
  XNOR2_X1 U416 ( .A(n410), .B(n409), .ZN(n496) );
  XNOR2_X1 U417 ( .A(G107), .B(G104), .ZN(n410) );
  XNOR2_X1 U418 ( .A(n424), .B(n423), .ZN(n492) );
  XNOR2_X1 U419 ( .A(n467), .B(n405), .ZN(n404) );
  XNOR2_X1 U420 ( .A(G107), .B(KEYINPUT9), .ZN(n467) );
  XNOR2_X1 U421 ( .A(KEYINPUT106), .B(KEYINPUT7), .ZN(n405) );
  XNOR2_X1 U422 ( .A(G116), .B(G134), .ZN(n466) );
  NOR2_X2 U423 ( .A1(n408), .A2(n554), .ZN(n587) );
  XNOR2_X1 U424 ( .A(n462), .B(G475), .ZN(n463) );
  INV_X1 U425 ( .A(KEYINPUT6), .ZN(n386) );
  XOR2_X1 U426 ( .A(KEYINPUT102), .B(KEYINPUT11), .Z(n452) );
  INV_X1 U427 ( .A(KEYINPUT85), .ZN(n400) );
  NOR2_X1 U428 ( .A1(n396), .A2(n593), .ZN(n395) );
  XNOR2_X1 U429 ( .A(n398), .B(n397), .ZN(n396) );
  INV_X1 U430 ( .A(KEYINPUT81), .ZN(n397) );
  NOR2_X1 U431 ( .A1(n682), .A2(n378), .ZN(n377) );
  INV_X1 U432 ( .A(n544), .ZN(n373) );
  XNOR2_X1 U433 ( .A(n465), .B(n415), .ZN(n484) );
  XNOR2_X1 U434 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n418) );
  XNOR2_X1 U435 ( .A(KEYINPUT15), .B(G902), .ZN(n656) );
  AND2_X1 U436 ( .A1(n392), .A2(n391), .ZN(n390) );
  NAND2_X1 U437 ( .A1(n393), .A2(G902), .ZN(n391) );
  XNOR2_X1 U438 ( .A(G128), .B(G110), .ZN(n506) );
  XNOR2_X1 U439 ( .A(n731), .B(n455), .ZN(n461) );
  XNOR2_X1 U440 ( .A(n596), .B(n595), .ZN(n379) );
  NAND2_X1 U441 ( .A1(n529), .A2(n580), .ZN(n524) );
  XNOR2_X1 U442 ( .A(n407), .B(n406), .ZN(n597) );
  INV_X1 U443 ( .A(KEYINPUT39), .ZN(n406) );
  NAND2_X1 U444 ( .A1(n403), .A2(n535), .ZN(n578) );
  XNOR2_X1 U445 ( .A(n515), .B(KEYINPUT25), .ZN(n516) );
  BUF_X1 U446 ( .A(n523), .Z(n629) );
  XNOR2_X1 U447 ( .A(n496), .B(n426), .ZN(n384) );
  XNOR2_X1 U448 ( .A(KEYINPUT74), .B(KEYINPUT16), .ZN(n425) );
  XNOR2_X1 U449 ( .A(n468), .B(n404), .ZN(n472) );
  BUF_X1 U450 ( .A(n714), .Z(n725) );
  OR2_X1 U451 ( .A1(n585), .A2(n586), .ZN(n401) );
  NOR2_X1 U452 ( .A1(n541), .A2(n519), .ZN(n371) );
  XNOR2_X1 U453 ( .A(n578), .B(n402), .ZN(n705) );
  INV_X1 U454 ( .A(KEYINPUT109), .ZN(n402) );
  INV_X1 U455 ( .A(n592), .ZN(n667) );
  OR2_X1 U456 ( .A1(n727), .A2(G902), .ZN(n354) );
  XNOR2_X1 U457 ( .A(n464), .B(n463), .ZN(n536) );
  INV_X1 U458 ( .A(n536), .ZN(n403) );
  AND2_X1 U459 ( .A1(n542), .A2(n668), .ZN(n355) );
  AND2_X1 U460 ( .A1(n399), .A2(n395), .ZN(n356) );
  AND2_X1 U461 ( .A1(n589), .A2(n588), .ZN(n358) );
  XOR2_X1 U462 ( .A(KEYINPUT53), .B(n654), .Z(G75) );
  XOR2_X1 U463 ( .A(n521), .B(n520), .Z(n360) );
  XOR2_X1 U464 ( .A(KEYINPUT68), .B(KEYINPUT19), .Z(n361) );
  INV_X1 U465 ( .A(G469), .ZN(n393) );
  XNOR2_X1 U466 ( .A(n502), .B(n501), .ZN(n715) );
  XNOR2_X1 U467 ( .A(n502), .B(n493), .ZN(n658) );
  XOR2_X1 U468 ( .A(n658), .B(n661), .Z(n362) );
  XOR2_X1 U469 ( .A(n688), .B(n691), .Z(n363) );
  XNOR2_X1 U470 ( .A(KEYINPUT59), .B(n684), .ZN(n364) );
  XNOR2_X1 U471 ( .A(n492), .B(n384), .ZN(n676) );
  OR2_X1 U472 ( .A1(KEYINPUT65), .A2(KEYINPUT44), .ZN(n365) );
  XNOR2_X1 U473 ( .A(n394), .B(n484), .ZN(n730) );
  INV_X1 U474 ( .A(n729), .ZN(n367) );
  INV_X1 U475 ( .A(n688), .ZN(n427) );
  XNOR2_X1 U476 ( .A(n382), .B(n676), .ZN(n688) );
  NAND2_X1 U477 ( .A1(n366), .A2(n365), .ZN(n543) );
  NAND2_X1 U478 ( .A1(n376), .A2(n377), .ZN(n366) );
  XNOR2_X1 U479 ( .A(n662), .B(n362), .ZN(n368) );
  XNOR2_X1 U480 ( .A(n692), .B(n363), .ZN(n369) );
  XNOR2_X1 U481 ( .A(n685), .B(n364), .ZN(n370) );
  NAND2_X1 U482 ( .A1(n544), .A2(n522), .ZN(n376) );
  INV_X1 U483 ( .A(KEYINPUT44), .ZN(n378) );
  INV_X1 U484 ( .A(n610), .ZN(n380) );
  XNOR2_X2 U485 ( .A(n381), .B(KEYINPUT45), .ZN(n669) );
  XNOR2_X1 U486 ( .A(n582), .B(n361), .ZN(n569) );
  XNOR2_X2 U487 ( .A(n436), .B(KEYINPUT86), .ZN(n582) );
  XNOR2_X1 U488 ( .A(n383), .B(n484), .ZN(n382) );
  XNOR2_X1 U489 ( .A(n419), .B(n420), .ZN(n383) );
  NAND2_X1 U490 ( .A1(n385), .A2(n648), .ZN(n526) );
  NAND2_X1 U491 ( .A1(n385), .A2(n534), .ZN(n695) );
  XNOR2_X1 U492 ( .A(n530), .B(KEYINPUT96), .ZN(n385) );
  INV_X1 U493 ( .A(n545), .ZN(n561) );
  XNOR2_X2 U494 ( .A(n495), .B(G472), .ZN(n545) );
  NAND2_X1 U495 ( .A1(n587), .A2(n358), .ZN(n592) );
  OR2_X1 U496 ( .A1(n715), .A2(n389), .ZN(n388) );
  NAND2_X1 U497 ( .A1(G469), .A2(n494), .ZN(n389) );
  NAND2_X1 U498 ( .A1(n715), .A2(n393), .ZN(n392) );
  XNOR2_X1 U499 ( .A(n486), .B(G137), .ZN(n394) );
  INV_X1 U500 ( .A(n401), .ZN(n712) );
  INV_X1 U501 ( .A(n535), .ZN(n537) );
  NOR2_X1 U502 ( .A1(n705), .A2(n579), .ZN(n581) );
  NAND2_X1 U503 ( .A1(n587), .A2(n617), .ZN(n407) );
  XNOR2_X2 U504 ( .A(n533), .B(KEYINPUT100), .ZN(n554) );
  NAND2_X1 U505 ( .A1(n553), .A2(n599), .ZN(n408) );
  AND2_X1 U506 ( .A1(n669), .A2(n609), .ZN(n607) );
  BUF_X1 U507 ( .A(n555), .Z(n604) );
  NOR2_X2 U508 ( .A1(n657), .A2(n656), .ZN(n714) );
  XOR2_X1 U509 ( .A(n447), .B(KEYINPUT0), .Z(n413) );
  XNOR2_X1 U510 ( .A(n449), .B(n418), .ZN(n419) );
  XNOR2_X1 U511 ( .A(n655), .B(KEYINPUT2), .ZN(n657) );
  INV_X1 U512 ( .A(KEYINPUT40), .ZN(n557) );
  INV_X1 U513 ( .A(KEYINPUT63), .ZN(n664) );
  INV_X1 U514 ( .A(KEYINPUT4), .ZN(n415) );
  NAND2_X1 U515 ( .A1(n469), .A2(G224), .ZN(n416) );
  XNOR2_X1 U516 ( .A(n416), .B(KEYINPUT78), .ZN(n420) );
  XNOR2_X1 U517 ( .A(G116), .B(G113), .ZN(n422) );
  XNOR2_X1 U518 ( .A(G101), .B(KEYINPUT72), .ZN(n421) );
  XNOR2_X1 U519 ( .A(n422), .B(n421), .ZN(n424) );
  XNOR2_X1 U520 ( .A(KEYINPUT3), .B(G119), .ZN(n423) );
  XNOR2_X1 U521 ( .A(n425), .B(G122), .ZN(n426) );
  NAND2_X1 U522 ( .A1(n427), .A2(n656), .ZN(n432) );
  INV_X1 U523 ( .A(G902), .ZN(n494) );
  INV_X1 U524 ( .A(G237), .ZN(n428) );
  NAND2_X1 U525 ( .A1(n494), .A2(n428), .ZN(n433) );
  NAND2_X1 U526 ( .A1(n433), .A2(G210), .ZN(n430) );
  INV_X1 U527 ( .A(KEYINPUT91), .ZN(n429) );
  XNOR2_X1 U528 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U529 ( .A(n432), .B(n431), .ZN(n555) );
  NAND2_X1 U530 ( .A1(n433), .A2(G214), .ZN(n434) );
  XNOR2_X1 U531 ( .A(n434), .B(KEYINPUT92), .ZN(n616) );
  INV_X1 U532 ( .A(n616), .ZN(n435) );
  NOR2_X2 U533 ( .A1(n555), .A2(n435), .ZN(n436) );
  XOR2_X1 U534 ( .A(KEYINPUT93), .B(KEYINPUT14), .Z(n438) );
  NAND2_X1 U535 ( .A1(G234), .A2(G237), .ZN(n437) );
  XNOR2_X1 U536 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U537 ( .A(KEYINPUT76), .B(n439), .ZN(n443) );
  NAND2_X1 U538 ( .A1(G952), .A2(n443), .ZN(n441) );
  INV_X1 U539 ( .A(KEYINPUT94), .ZN(n440) );
  XNOR2_X1 U540 ( .A(n441), .B(n440), .ZN(n645) );
  NAND2_X1 U541 ( .A1(n645), .A2(n469), .ZN(n442) );
  XNOR2_X1 U542 ( .A(n442), .B(KEYINPUT95), .ZN(n548) );
  NAND2_X1 U543 ( .A1(G902), .A2(n443), .ZN(n549) );
  NOR2_X1 U544 ( .A1(G898), .A2(n469), .ZN(n677) );
  INV_X1 U545 ( .A(n677), .ZN(n444) );
  NOR2_X1 U546 ( .A1(n549), .A2(n444), .ZN(n445) );
  OR2_X1 U547 ( .A1(n548), .A2(n445), .ZN(n446) );
  NAND2_X1 U548 ( .A1(n569), .A2(n446), .ZN(n448) );
  INV_X1 U549 ( .A(KEYINPUT69), .ZN(n447) );
  XNOR2_X2 U550 ( .A(n448), .B(n413), .ZN(n530) );
  XNOR2_X1 U551 ( .A(n449), .B(G140), .ZN(n450) );
  XNOR2_X1 U552 ( .A(n450), .B(KEYINPUT10), .ZN(n731) );
  XOR2_X1 U553 ( .A(n452), .B(n451), .Z(n454) );
  NOR2_X1 U554 ( .A1(G953), .A2(G237), .ZN(n488) );
  NAND2_X1 U555 ( .A1(G214), .A2(n488), .ZN(n453) );
  XNOR2_X1 U556 ( .A(n485), .B(KEYINPUT104), .ZN(n459) );
  XNOR2_X1 U557 ( .A(G113), .B(G143), .ZN(n456) );
  XNOR2_X1 U558 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U559 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U560 ( .A(n461), .B(n460), .ZN(n684) );
  NOR2_X1 U561 ( .A1(G902), .A2(n684), .ZN(n464) );
  XNOR2_X1 U562 ( .A(KEYINPUT13), .B(KEYINPUT105), .ZN(n462) );
  XNOR2_X1 U563 ( .A(n466), .B(G122), .ZN(n468) );
  NAND2_X1 U564 ( .A1(G234), .A2(n469), .ZN(n470) );
  XOR2_X1 U565 ( .A(KEYINPUT8), .B(n470), .Z(n510) );
  NAND2_X1 U566 ( .A1(G217), .A2(n510), .ZN(n471) );
  XNOR2_X1 U567 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U568 ( .A(n465), .B(n473), .ZN(n721) );
  NOR2_X1 U569 ( .A1(G902), .A2(n721), .ZN(n475) );
  XOR2_X1 U570 ( .A(KEYINPUT107), .B(G478), .Z(n474) );
  XNOR2_X1 U571 ( .A(n475), .B(n474), .ZN(n535) );
  AND2_X1 U572 ( .A1(n536), .A2(n535), .ZN(n615) );
  XOR2_X1 U573 ( .A(KEYINPUT99), .B(KEYINPUT21), .Z(n478) );
  NAND2_X1 U574 ( .A1(G234), .A2(n656), .ZN(n476) );
  XNOR2_X1 U575 ( .A(KEYINPUT20), .B(n476), .ZN(n514) );
  NAND2_X1 U576 ( .A1(G221), .A2(n514), .ZN(n477) );
  XNOR2_X1 U577 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U578 ( .A(KEYINPUT98), .B(n479), .ZN(n631) );
  INV_X1 U579 ( .A(n631), .ZN(n480) );
  AND2_X1 U580 ( .A1(n615), .A2(n480), .ZN(n481) );
  XNOR2_X1 U581 ( .A(n481), .B(KEYINPUT108), .ZN(n482) );
  NAND2_X1 U582 ( .A1(n530), .A2(n482), .ZN(n483) );
  INV_X1 U583 ( .A(n541), .ZN(n504) );
  XOR2_X1 U584 ( .A(n485), .B(G134), .Z(n486) );
  XOR2_X1 U585 ( .A(KEYINPUT5), .B(KEYINPUT101), .Z(n490) );
  NAND2_X1 U586 ( .A1(n488), .A2(G210), .ZN(n489) );
  XNOR2_X1 U587 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U588 ( .A(n492), .B(n491), .ZN(n493) );
  NAND2_X1 U589 ( .A1(n658), .A2(n494), .ZN(n495) );
  INV_X1 U590 ( .A(n496), .ZN(n500) );
  XOR2_X1 U591 ( .A(G101), .B(G140), .Z(n498) );
  NAND2_X1 U592 ( .A1(G227), .A2(n469), .ZN(n497) );
  XNOR2_X1 U593 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U594 ( .A(n500), .B(n499), .ZN(n501) );
  AND2_X1 U595 ( .A1(n561), .A2(n629), .ZN(n503) );
  XNOR2_X1 U596 ( .A(G119), .B(G137), .ZN(n505) );
  XNOR2_X1 U597 ( .A(n505), .B(KEYINPUT97), .ZN(n509) );
  XOR2_X1 U598 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n507) );
  XNOR2_X1 U599 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U600 ( .A(n509), .B(n508), .Z(n512) );
  NAND2_X1 U601 ( .A1(G221), .A2(n510), .ZN(n511) );
  XNOR2_X1 U602 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U603 ( .A(n731), .B(n513), .ZN(n727) );
  NAND2_X1 U604 ( .A1(n514), .A2(G217), .ZN(n515) );
  XNOR2_X2 U605 ( .A(n354), .B(n516), .ZN(n632) );
  INV_X1 U606 ( .A(n632), .ZN(n559) );
  INV_X1 U607 ( .A(KEYINPUT89), .ZN(n517) );
  XNOR2_X1 U608 ( .A(n523), .B(n517), .ZN(n586) );
  OR2_X1 U609 ( .A1(n586), .A2(n518), .ZN(n519) );
  XNOR2_X1 U610 ( .A(KEYINPUT79), .B(KEYINPUT32), .ZN(n521) );
  INV_X1 U611 ( .A(KEYINPUT66), .ZN(n520) );
  INV_X1 U612 ( .A(KEYINPUT65), .ZN(n522) );
  XNOR2_X2 U613 ( .A(n524), .B(KEYINPUT33), .ZN(n648) );
  XNOR2_X1 U614 ( .A(KEYINPUT73), .B(KEYINPUT34), .ZN(n525) );
  XNOR2_X1 U615 ( .A(n526), .B(n525), .ZN(n527) );
  NOR2_X1 U616 ( .A1(n536), .A2(n535), .ZN(n589) );
  NAND2_X1 U617 ( .A1(n527), .A2(n589), .ZN(n528) );
  BUF_X1 U618 ( .A(n545), .Z(n635) );
  NAND2_X1 U619 ( .A1(n529), .A2(n635), .ZN(n638) );
  INV_X1 U620 ( .A(n530), .ZN(n531) );
  NOR2_X1 U621 ( .A1(n638), .A2(n531), .ZN(n532) );
  XNOR2_X1 U622 ( .A(n532), .B(KEYINPUT31), .ZN(n708) );
  OR2_X2 U623 ( .A1(n628), .A2(n563), .ZN(n533) );
  NOR2_X1 U624 ( .A1(n554), .A2(n635), .ZN(n534) );
  NAND2_X1 U625 ( .A1(n708), .A2(n695), .ZN(n538) );
  NAND2_X1 U626 ( .A1(n536), .A2(n537), .ZN(n709) );
  NAND2_X1 U627 ( .A1(n578), .A2(n709), .ZN(n622) );
  NAND2_X1 U628 ( .A1(n538), .A2(n622), .ZN(n542) );
  NOR2_X1 U629 ( .A1(n580), .A2(n632), .ZN(n539) );
  NAND2_X1 U630 ( .A1(n539), .A2(n629), .ZN(n540) );
  OR2_X1 U631 ( .A1(n541), .A2(n540), .ZN(n668) );
  NAND2_X1 U632 ( .A1(n545), .A2(n616), .ZN(n547) );
  XOR2_X1 U633 ( .A(KEYINPUT110), .B(KEYINPUT30), .Z(n546) );
  XNOR2_X1 U634 ( .A(n547), .B(n546), .ZN(n553) );
  INV_X1 U635 ( .A(n548), .ZN(n552) );
  NOR2_X1 U636 ( .A1(G900), .A2(n549), .ZN(n550) );
  NAND2_X1 U637 ( .A1(G953), .A2(n550), .ZN(n551) );
  NAND2_X1 U638 ( .A1(n552), .A2(n551), .ZN(n599) );
  XOR2_X1 U639 ( .A(KEYINPUT77), .B(KEYINPUT38), .Z(n556) );
  XNOR2_X1 U640 ( .A(n604), .B(n556), .ZN(n617) );
  XNOR2_X1 U641 ( .A(n558), .B(n557), .ZN(n740) );
  NOR2_X1 U642 ( .A1(n631), .A2(n559), .ZN(n577) );
  NAND2_X1 U643 ( .A1(n577), .A2(n599), .ZN(n560) );
  NOR2_X1 U644 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U645 ( .A(KEYINPUT28), .B(n562), .Z(n564) );
  NOR2_X1 U646 ( .A1(n564), .A2(n563), .ZN(n570) );
  AND2_X1 U647 ( .A1(n617), .A2(n616), .ZN(n623) );
  NAND2_X1 U648 ( .A1(n615), .A2(n623), .ZN(n565) );
  XNOR2_X1 U649 ( .A(n565), .B(KEYINPUT41), .ZN(n647) );
  NAND2_X1 U650 ( .A1(n570), .A2(n647), .ZN(n566) );
  XNOR2_X1 U651 ( .A(n566), .B(KEYINPUT42), .ZN(n741) );
  NAND2_X1 U652 ( .A1(n740), .A2(n741), .ZN(n568) );
  XOR2_X1 U653 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n567) );
  XNOR2_X1 U654 ( .A(n568), .B(n567), .ZN(n594) );
  AND2_X1 U655 ( .A1(n569), .A2(n570), .ZN(n574) );
  XOR2_X1 U656 ( .A(KEYINPUT47), .B(KEYINPUT70), .Z(n571) );
  NAND2_X1 U657 ( .A1(n571), .A2(n622), .ZN(n572) );
  XNOR2_X1 U658 ( .A(n572), .B(KEYINPUT75), .ZN(n573) );
  NAND2_X1 U659 ( .A1(n574), .A2(n573), .ZN(n576) );
  INV_X1 U660 ( .A(n574), .ZN(n703) );
  NAND2_X1 U661 ( .A1(n703), .A2(KEYINPUT47), .ZN(n575) );
  NAND2_X1 U662 ( .A1(n576), .A2(n575), .ZN(n593) );
  INV_X1 U663 ( .A(n577), .ZN(n579) );
  NAND2_X1 U664 ( .A1(n581), .A2(n580), .ZN(n601) );
  NAND2_X1 U665 ( .A1(n582), .A2(n599), .ZN(n583) );
  NOR2_X1 U666 ( .A1(n601), .A2(n583), .ZN(n584) );
  XOR2_X1 U667 ( .A(KEYINPUT36), .B(n584), .Z(n585) );
  INV_X1 U668 ( .A(n604), .ZN(n588) );
  INV_X1 U669 ( .A(n622), .ZN(n590) );
  NAND2_X1 U670 ( .A1(n590), .A2(KEYINPUT47), .ZN(n591) );
  NAND2_X1 U671 ( .A1(n594), .A2(n356), .ZN(n596) );
  XOR2_X1 U672 ( .A(KEYINPUT48), .B(KEYINPUT84), .Z(n595) );
  NOR2_X1 U673 ( .A1(n597), .A2(n709), .ZN(n598) );
  XOR2_X1 U674 ( .A(KEYINPUT111), .B(n598), .Z(n739) );
  NAND2_X1 U675 ( .A1(n616), .A2(n599), .ZN(n600) );
  NOR2_X1 U676 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U677 ( .A1(n629), .A2(n602), .ZN(n603) );
  XNOR2_X1 U678 ( .A(n603), .B(KEYINPUT43), .ZN(n605) );
  AND2_X1 U679 ( .A1(n605), .A2(n604), .ZN(n680) );
  NOR2_X1 U680 ( .A1(n739), .A2(n680), .ZN(n606) );
  INV_X1 U681 ( .A(KEYINPUT2), .ZN(n609) );
  NOR2_X1 U682 ( .A1(n655), .A2(n609), .ZN(n608) );
  NOR2_X1 U683 ( .A1(n608), .A2(n607), .ZN(n613) );
  NAND2_X1 U684 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U685 ( .A(KEYINPUT82), .B(n611), .Z(n612) );
  NOR2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U687 ( .A(n614), .B(KEYINPUT83), .ZN(n653) );
  INV_X1 U688 ( .A(n615), .ZN(n620) );
  NOR2_X1 U689 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U690 ( .A(n618), .B(KEYINPUT118), .ZN(n619) );
  NOR2_X1 U691 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U692 ( .A(n621), .B(KEYINPUT119), .ZN(n625) );
  NAND2_X1 U693 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U694 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U695 ( .A1(n648), .A2(n626), .ZN(n627) );
  XNOR2_X1 U696 ( .A(n627), .B(KEYINPUT120), .ZN(n643) );
  NAND2_X1 U697 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U698 ( .A(n630), .B(KEYINPUT50), .ZN(n637) );
  NAND2_X1 U699 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U700 ( .A(KEYINPUT49), .B(n633), .ZN(n634) );
  NOR2_X1 U701 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U702 ( .A1(n637), .A2(n636), .ZN(n639) );
  NAND2_X1 U703 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U704 ( .A(KEYINPUT51), .B(n640), .Z(n641) );
  NAND2_X1 U705 ( .A1(n647), .A2(n641), .ZN(n642) );
  NAND2_X1 U706 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U707 ( .A(n644), .B(KEYINPUT52), .ZN(n646) );
  AND2_X1 U708 ( .A1(n646), .A2(n645), .ZN(n651) );
  NAND2_X1 U709 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U710 ( .A1(n649), .A2(n469), .ZN(n650) );
  NOR2_X1 U711 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U712 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U713 ( .A1(n714), .A2(G472), .ZN(n662) );
  XNOR2_X1 U714 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n660) );
  XNOR2_X1 U715 ( .A(KEYINPUT62), .B(KEYINPUT88), .ZN(n659) );
  XNOR2_X1 U716 ( .A(n660), .B(n659), .ZN(n661) );
  INV_X1 U717 ( .A(G952), .ZN(n663) );
  AND2_X1 U718 ( .A1(n663), .A2(G953), .ZN(n729) );
  XNOR2_X1 U719 ( .A(n665), .B(n664), .ZN(G57) );
  INV_X1 U720 ( .A(G143), .ZN(n666) );
  XNOR2_X1 U721 ( .A(n667), .B(n666), .ZN(G45) );
  XNOR2_X1 U722 ( .A(n668), .B(G101), .ZN(G3) );
  NAND2_X1 U723 ( .A1(n669), .A2(n469), .ZN(n675) );
  XOR2_X1 U724 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n671) );
  NAND2_X1 U725 ( .A1(G224), .A2(G953), .ZN(n670) );
  XNOR2_X1 U726 ( .A(n671), .B(n670), .ZN(n672) );
  NAND2_X1 U727 ( .A1(G898), .A2(n672), .ZN(n673) );
  XNOR2_X1 U728 ( .A(n673), .B(KEYINPUT126), .ZN(n674) );
  NAND2_X1 U729 ( .A1(n675), .A2(n674), .ZN(n679) );
  NOR2_X1 U730 ( .A1(n676), .A2(n677), .ZN(n678) );
  XNOR2_X1 U731 ( .A(n679), .B(n678), .ZN(G69) );
  XOR2_X1 U732 ( .A(n680), .B(G140), .Z(G42) );
  XNOR2_X1 U733 ( .A(n681), .B(G110), .ZN(G12) );
  XOR2_X1 U734 ( .A(n682), .B(G122), .Z(G24) );
  XNOR2_X1 U735 ( .A(n683), .B(G119), .ZN(G21) );
  NAND2_X1 U736 ( .A1(n714), .A2(G475), .ZN(n685) );
  XOR2_X1 U737 ( .A(KEYINPUT123), .B(KEYINPUT60), .Z(n686) );
  XNOR2_X1 U738 ( .A(n687), .B(n686), .ZN(G60) );
  NAND2_X1 U739 ( .A1(n714), .A2(G210), .ZN(n692) );
  XOR2_X1 U740 ( .A(KEYINPUT55), .B(KEYINPUT87), .Z(n690) );
  XNOR2_X1 U741 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n689) );
  XNOR2_X1 U742 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U743 ( .A(n693), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X1 U744 ( .A1(n705), .A2(n695), .ZN(n694) );
  XOR2_X1 U745 ( .A(G104), .B(n694), .Z(G6) );
  NOR2_X1 U746 ( .A1(n709), .A2(n695), .ZN(n700) );
  XOR2_X1 U747 ( .A(KEYINPUT27), .B(KEYINPUT115), .Z(n697) );
  XNOR2_X1 U748 ( .A(G107), .B(KEYINPUT114), .ZN(n696) );
  XNOR2_X1 U749 ( .A(n697), .B(n696), .ZN(n698) );
  XNOR2_X1 U750 ( .A(KEYINPUT26), .B(n698), .ZN(n699) );
  XNOR2_X1 U751 ( .A(n700), .B(n699), .ZN(G9) );
  NOR2_X1 U752 ( .A1(n703), .A2(n709), .ZN(n702) );
  XNOR2_X1 U753 ( .A(G128), .B(KEYINPUT29), .ZN(n701) );
  XNOR2_X1 U754 ( .A(n702), .B(n701), .ZN(G30) );
  NOR2_X1 U755 ( .A1(n703), .A2(n705), .ZN(n704) );
  XOR2_X1 U756 ( .A(G146), .B(n704), .Z(G48) );
  NOR2_X1 U757 ( .A1(n705), .A2(n708), .ZN(n706) );
  XOR2_X1 U758 ( .A(KEYINPUT116), .B(n706), .Z(n707) );
  XNOR2_X1 U759 ( .A(G113), .B(n707), .ZN(G15) );
  NOR2_X1 U760 ( .A1(n709), .A2(n708), .ZN(n711) );
  XNOR2_X1 U761 ( .A(G116), .B(KEYINPUT117), .ZN(n710) );
  XNOR2_X1 U762 ( .A(n711), .B(n710), .ZN(G18) );
  XNOR2_X1 U763 ( .A(G125), .B(n712), .ZN(n713) );
  XNOR2_X1 U764 ( .A(n713), .B(KEYINPUT37), .ZN(G27) );
  NAND2_X1 U765 ( .A1(n725), .A2(G469), .ZN(n719) );
  XOR2_X1 U766 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n717) );
  XNOR2_X1 U767 ( .A(n715), .B(KEYINPUT122), .ZN(n716) );
  XNOR2_X1 U768 ( .A(n717), .B(n716), .ZN(n718) );
  XNOR2_X1 U769 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U770 ( .A1(n729), .A2(n720), .ZN(G54) );
  NAND2_X1 U771 ( .A1(n725), .A2(G478), .ZN(n723) );
  XNOR2_X1 U772 ( .A(n721), .B(KEYINPUT124), .ZN(n722) );
  XNOR2_X1 U773 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U774 ( .A1(n729), .A2(n724), .ZN(G63) );
  NAND2_X1 U775 ( .A1(n725), .A2(G217), .ZN(n726) );
  XNOR2_X1 U776 ( .A(n727), .B(n726), .ZN(n728) );
  NOR2_X1 U777 ( .A1(n729), .A2(n728), .ZN(G66) );
  XNOR2_X1 U778 ( .A(n730), .B(n731), .ZN(n734) );
  XNOR2_X1 U779 ( .A(G227), .B(n734), .ZN(n732) );
  NAND2_X1 U780 ( .A1(n732), .A2(G900), .ZN(n733) );
  NAND2_X1 U781 ( .A1(n733), .A2(G953), .ZN(n738) );
  XOR2_X1 U782 ( .A(n734), .B(n610), .Z(n735) );
  XNOR2_X1 U783 ( .A(n735), .B(KEYINPUT127), .ZN(n736) );
  NAND2_X1 U784 ( .A1(n736), .A2(n469), .ZN(n737) );
  NAND2_X1 U785 ( .A1(n738), .A2(n737), .ZN(G72) );
  XOR2_X1 U786 ( .A(G134), .B(n739), .Z(G36) );
  XNOR2_X1 U787 ( .A(n740), .B(G131), .ZN(G33) );
  XNOR2_X1 U788 ( .A(G137), .B(n741), .ZN(G39) );
endmodule

