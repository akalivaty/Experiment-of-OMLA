

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U553 ( .A1(G2104), .A2(n556), .ZN(n902) );
  AND2_X1 U554 ( .A1(n556), .A2(G2104), .ZN(n906) );
  INV_X1 U555 ( .A(n762), .ZN(n738) );
  XNOR2_X1 U556 ( .A(n565), .B(n564), .ZN(G164) );
  NOR2_X1 U557 ( .A1(n725), .A2(n942), .ZN(n734) );
  NAND2_X1 U558 ( .A1(n553), .A2(n552), .ZN(n724) );
  NOR2_X1 U559 ( .A1(G164), .A2(n554), .ZN(n553) );
  NAND2_X1 U560 ( .A1(n532), .A2(n521), .ZN(n531) );
  NAND2_X1 U561 ( .A1(n533), .A2(KEYINPUT29), .ZN(n532) );
  INV_X1 U562 ( .A(G8), .ZN(n550) );
  OR2_X1 U563 ( .A1(n768), .A2(n544), .ZN(n543) );
  AND2_X1 U564 ( .A1(n546), .A2(n545), .ZN(n544) );
  NAND2_X1 U565 ( .A1(n525), .A2(n547), .ZN(n546) );
  NAND2_X1 U566 ( .A1(n769), .A2(KEYINPUT98), .ZN(n545) );
  NAND2_X1 U567 ( .A1(n542), .A2(n541), .ZN(n540) );
  NAND2_X1 U568 ( .A1(n525), .A2(KEYINPUT98), .ZN(n542) );
  NAND2_X1 U569 ( .A1(n769), .A2(n547), .ZN(n541) );
  NOR2_X1 U570 ( .A1(n683), .A2(n573), .ZN(n669) );
  NAND2_X1 U571 ( .A1(G1996), .A2(n555), .ZN(n554) );
  INV_X1 U572 ( .A(G1384), .ZN(n555) );
  INV_X1 U573 ( .A(KEYINPUT96), .ZN(n727) );
  AND2_X1 U574 ( .A1(n726), .A2(n734), .ZN(n728) );
  AND2_X1 U575 ( .A1(n749), .A2(n536), .ZN(n528) );
  INV_X1 U576 ( .A(KEYINPUT98), .ZN(n547) );
  NOR2_X1 U577 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U578 ( .A1(n534), .A2(n531), .ZN(n760) );
  INV_X1 U579 ( .A(n804), .ZN(n552) );
  NAND2_X1 U580 ( .A1(n520), .A2(n549), .ZN(n548) );
  NAND2_X1 U581 ( .A1(n543), .A2(n539), .ZN(n551) );
  NAND2_X1 U582 ( .A1(n769), .A2(n550), .ZN(n549) );
  AND2_X1 U583 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U584 ( .A1(G164), .A2(G1384), .ZN(n805) );
  NAND2_X1 U585 ( .A1(n527), .A2(n556), .ZN(n526) );
  INV_X1 U586 ( .A(G2104), .ZN(n527) );
  NAND2_X1 U587 ( .A1(G2105), .A2(G2104), .ZN(n559) );
  XNOR2_X1 U588 ( .A(n627), .B(KEYINPUT15), .ZN(n940) );
  NOR2_X1 U589 ( .A1(G651), .A2(n683), .ZN(n677) );
  NOR2_X1 U590 ( .A1(G651), .A2(G543), .ZN(n667) );
  AND2_X1 U591 ( .A1(n744), .A2(KEYINPUT29), .ZN(n519) );
  OR2_X1 U592 ( .A1(n774), .A2(n773), .ZN(n520) );
  NAND2_X1 U593 ( .A1(n805), .A2(n552), .ZN(n762) );
  OR2_X1 U594 ( .A1(G301), .A2(n755), .ZN(n521) );
  OR2_X1 U595 ( .A1(n794), .A2(n961), .ZN(n522) );
  NOR2_X1 U596 ( .A1(n551), .A2(n548), .ZN(n794) );
  AND2_X1 U597 ( .A1(n946), .A2(n846), .ZN(n523) );
  NOR2_X1 U598 ( .A1(n833), .A2(n523), .ZN(n524) );
  AND2_X1 U599 ( .A1(KEYINPUT32), .A2(G8), .ZN(n525) );
  INV_X1 U600 ( .A(KEYINPUT29), .ZN(n536) );
  INV_X1 U601 ( .A(KEYINPUT32), .ZN(n769) );
  XNOR2_X2 U602 ( .A(n526), .B(KEYINPUT17), .ZN(n907) );
  NAND2_X1 U603 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U604 ( .A1(n745), .A2(n744), .ZN(n529) );
  NAND2_X1 U605 ( .A1(n530), .A2(n535), .ZN(n534) );
  NAND2_X1 U606 ( .A1(n745), .A2(n519), .ZN(n535) );
  INV_X1 U607 ( .A(n749), .ZN(n533) );
  NAND2_X1 U608 ( .A1(n537), .A2(n848), .ZN(n850) );
  NAND2_X1 U609 ( .A1(n538), .A2(n524), .ZN(n537) );
  NAND2_X1 U610 ( .A1(n802), .A2(n803), .ZN(n538) );
  NAND2_X1 U611 ( .A1(n768), .A2(n540), .ZN(n539) );
  XOR2_X2 U612 ( .A(KEYINPUT64), .B(n559), .Z(n903) );
  INV_X1 U613 ( .A(KEYINPUT95), .ZN(n739) );
  XNOR2_X1 U614 ( .A(n739), .B(KEYINPUT27), .ZN(n740) );
  XNOR2_X1 U615 ( .A(n741), .B(n740), .ZN(n743) );
  INV_X1 U616 ( .A(n798), .ZN(n782) );
  XNOR2_X1 U617 ( .A(KEYINPUT72), .B(KEYINPUT12), .ZN(n611) );
  XNOR2_X1 U618 ( .A(n612), .B(n611), .ZN(n614) );
  AND2_X1 U619 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U620 ( .A1(n722), .A2(n721), .ZN(n804) );
  INV_X1 U621 ( .A(KEYINPUT89), .ZN(n565) );
  INV_X1 U622 ( .A(G2105), .ZN(n556) );
  NAND2_X1 U623 ( .A1(G126), .A2(n902), .ZN(n558) );
  NAND2_X1 U624 ( .A1(G102), .A2(n906), .ZN(n557) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n563) );
  NAND2_X1 U626 ( .A1(G138), .A2(n907), .ZN(n561) );
  NAND2_X1 U627 ( .A1(G114), .A2(n903), .ZN(n560) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  INV_X1 U630 ( .A(G651), .ZN(n573) );
  NOR2_X1 U631 ( .A1(G543), .A2(n573), .ZN(n567) );
  XNOR2_X1 U632 ( .A(KEYINPUT69), .B(KEYINPUT1), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n681) );
  NAND2_X1 U634 ( .A1(G63), .A2(n681), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G543), .B(KEYINPUT0), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n568), .B(KEYINPUT67), .ZN(n683) );
  NAND2_X1 U637 ( .A1(G51), .A2(n677), .ZN(n569) );
  NAND2_X1 U638 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U639 ( .A(KEYINPUT6), .B(n571), .ZN(n579) );
  NAND2_X1 U640 ( .A1(n667), .A2(G89), .ZN(n572) );
  XNOR2_X1 U641 ( .A(n572), .B(KEYINPUT4), .ZN(n575) );
  NAND2_X1 U642 ( .A1(G76), .A2(n669), .ZN(n574) );
  NAND2_X1 U643 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U644 ( .A(KEYINPUT5), .B(n576), .ZN(n577) );
  XNOR2_X1 U645 ( .A(KEYINPUT73), .B(n577), .ZN(n578) );
  NOR2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n581) );
  XOR2_X1 U647 ( .A(KEYINPUT74), .B(KEYINPUT7), .Z(n580) );
  XNOR2_X1 U648 ( .A(n581), .B(n580), .ZN(G168) );
  XOR2_X1 U649 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U650 ( .A1(G137), .A2(n907), .ZN(n583) );
  NAND2_X1 U651 ( .A1(G113), .A2(n903), .ZN(n582) );
  NAND2_X1 U652 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U653 ( .A(n584), .B(KEYINPUT65), .ZN(n722) );
  NAND2_X1 U654 ( .A1(G125), .A2(n902), .ZN(n719) );
  AND2_X1 U655 ( .A1(n722), .A2(n719), .ZN(n586) );
  NAND2_X1 U656 ( .A1(G101), .A2(n906), .ZN(n585) );
  XOR2_X1 U657 ( .A(KEYINPUT23), .B(n585), .Z(n718) );
  AND2_X1 U658 ( .A1(n586), .A2(n718), .ZN(G160) );
  AND2_X1 U659 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U660 ( .A1(G65), .A2(n681), .ZN(n588) );
  NAND2_X1 U661 ( .A1(G53), .A2(n677), .ZN(n587) );
  NAND2_X1 U662 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U663 ( .A1(G91), .A2(n667), .ZN(n590) );
  NAND2_X1 U664 ( .A1(G78), .A2(n669), .ZN(n589) );
  NAND2_X1 U665 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U666 ( .A1(n592), .A2(n591), .ZN(n746) );
  INV_X1 U667 ( .A(n746), .ZN(G299) );
  INV_X1 U668 ( .A(G57), .ZN(G237) );
  NAND2_X1 U669 ( .A1(G88), .A2(n667), .ZN(n594) );
  NAND2_X1 U670 ( .A1(G75), .A2(n669), .ZN(n593) );
  NAND2_X1 U671 ( .A1(n594), .A2(n593), .ZN(n598) );
  NAND2_X1 U672 ( .A1(G62), .A2(n681), .ZN(n596) );
  NAND2_X1 U673 ( .A1(G50), .A2(n677), .ZN(n595) );
  NAND2_X1 U674 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U675 ( .A1(n598), .A2(n597), .ZN(G166) );
  NAND2_X1 U676 ( .A1(G64), .A2(n681), .ZN(n599) );
  XOR2_X1 U677 ( .A(KEYINPUT70), .B(n599), .Z(n606) );
  NAND2_X1 U678 ( .A1(G90), .A2(n667), .ZN(n601) );
  NAND2_X1 U679 ( .A1(G77), .A2(n669), .ZN(n600) );
  NAND2_X1 U680 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U681 ( .A(n602), .B(KEYINPUT9), .ZN(n604) );
  NAND2_X1 U682 ( .A1(G52), .A2(n677), .ZN(n603) );
  NAND2_X1 U683 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U684 ( .A1(n606), .A2(n605), .ZN(G171) );
  NAND2_X1 U685 ( .A1(G7), .A2(G661), .ZN(n607) );
  XNOR2_X1 U686 ( .A(n607), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U687 ( .A(G223), .ZN(n851) );
  NAND2_X1 U688 ( .A1(n851), .A2(G567), .ZN(n608) );
  XNOR2_X1 U689 ( .A(n608), .B(KEYINPUT11), .ZN(n609) );
  XNOR2_X1 U690 ( .A(KEYINPUT71), .B(n609), .ZN(G234) );
  NAND2_X1 U691 ( .A1(G56), .A2(n681), .ZN(n610) );
  XOR2_X1 U692 ( .A(KEYINPUT14), .B(n610), .Z(n617) );
  NAND2_X1 U693 ( .A1(G81), .A2(n667), .ZN(n612) );
  NAND2_X1 U694 ( .A1(G68), .A2(n669), .ZN(n613) );
  NAND2_X1 U695 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U696 ( .A(KEYINPUT13), .B(n615), .Z(n616) );
  NOR2_X1 U697 ( .A1(n617), .A2(n616), .ZN(n619) );
  NAND2_X1 U698 ( .A1(n677), .A2(G43), .ZN(n618) );
  NAND2_X1 U699 ( .A1(n619), .A2(n618), .ZN(n942) );
  INV_X1 U700 ( .A(n942), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n620), .A2(G860), .ZN(G153) );
  INV_X1 U702 ( .A(G171), .ZN(G301) );
  NAND2_X1 U703 ( .A1(G868), .A2(G301), .ZN(n629) );
  NAND2_X1 U704 ( .A1(G79), .A2(n669), .ZN(n622) );
  NAND2_X1 U705 ( .A1(G54), .A2(n677), .ZN(n621) );
  NAND2_X1 U706 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U707 ( .A1(G92), .A2(n667), .ZN(n624) );
  NAND2_X1 U708 ( .A1(G66), .A2(n681), .ZN(n623) );
  NAND2_X1 U709 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U710 ( .A1(n626), .A2(n625), .ZN(n627) );
  INV_X1 U711 ( .A(G868), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n940), .A2(n630), .ZN(n628) );
  NAND2_X1 U713 ( .A1(n629), .A2(n628), .ZN(G284) );
  NAND2_X1 U714 ( .A1(G868), .A2(G286), .ZN(n632) );
  NAND2_X1 U715 ( .A1(G299), .A2(n630), .ZN(n631) );
  NAND2_X1 U716 ( .A1(n632), .A2(n631), .ZN(G297) );
  INV_X1 U717 ( .A(G559), .ZN(n633) );
  NOR2_X1 U718 ( .A1(G860), .A2(n633), .ZN(n634) );
  XNOR2_X1 U719 ( .A(KEYINPUT75), .B(n634), .ZN(n635) );
  INV_X1 U720 ( .A(n940), .ZN(n723) );
  NAND2_X1 U721 ( .A1(n635), .A2(n723), .ZN(n636) );
  XNOR2_X1 U722 ( .A(n636), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U723 ( .A1(G868), .A2(n942), .ZN(n639) );
  NAND2_X1 U724 ( .A1(n723), .A2(G868), .ZN(n637) );
  NOR2_X1 U725 ( .A1(G559), .A2(n637), .ZN(n638) );
  NOR2_X1 U726 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U727 ( .A(KEYINPUT76), .B(n640), .ZN(G282) );
  NAND2_X1 U728 ( .A1(G123), .A2(n902), .ZN(n641) );
  XNOR2_X1 U729 ( .A(n641), .B(KEYINPUT18), .ZN(n644) );
  NAND2_X1 U730 ( .A1(G99), .A2(n906), .ZN(n642) );
  XOR2_X1 U731 ( .A(KEYINPUT77), .B(n642), .Z(n643) );
  NAND2_X1 U732 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U733 ( .A1(G135), .A2(n907), .ZN(n646) );
  NAND2_X1 U734 ( .A1(G111), .A2(n903), .ZN(n645) );
  NAND2_X1 U735 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U736 ( .A1(n648), .A2(n647), .ZN(n1017) );
  XNOR2_X1 U737 ( .A(G2096), .B(n1017), .ZN(n650) );
  INV_X1 U738 ( .A(G2100), .ZN(n649) );
  NAND2_X1 U739 ( .A1(n650), .A2(n649), .ZN(G156) );
  NAND2_X1 U740 ( .A1(G559), .A2(n723), .ZN(n651) );
  XNOR2_X1 U741 ( .A(n651), .B(n942), .ZN(n695) );
  NOR2_X1 U742 ( .A1(n695), .A2(G860), .ZN(n658) );
  NAND2_X1 U743 ( .A1(G67), .A2(n681), .ZN(n653) );
  NAND2_X1 U744 ( .A1(G55), .A2(n677), .ZN(n652) );
  NAND2_X1 U745 ( .A1(n653), .A2(n652), .ZN(n657) );
  NAND2_X1 U746 ( .A1(G93), .A2(n667), .ZN(n655) );
  NAND2_X1 U747 ( .A1(G80), .A2(n669), .ZN(n654) );
  NAND2_X1 U748 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U749 ( .A1(n657), .A2(n656), .ZN(n689) );
  XNOR2_X1 U750 ( .A(n658), .B(n689), .ZN(G145) );
  NAND2_X1 U751 ( .A1(G86), .A2(n667), .ZN(n660) );
  NAND2_X1 U752 ( .A1(G61), .A2(n681), .ZN(n659) );
  NAND2_X1 U753 ( .A1(n660), .A2(n659), .ZN(n664) );
  NAND2_X1 U754 ( .A1(G73), .A2(n669), .ZN(n661) );
  XNOR2_X1 U755 ( .A(n661), .B(KEYINPUT2), .ZN(n662) );
  XNOR2_X1 U756 ( .A(n662), .B(KEYINPUT79), .ZN(n663) );
  NOR2_X1 U757 ( .A1(n664), .A2(n663), .ZN(n666) );
  NAND2_X1 U758 ( .A1(n677), .A2(G48), .ZN(n665) );
  NAND2_X1 U759 ( .A1(n666), .A2(n665), .ZN(G305) );
  NAND2_X1 U760 ( .A1(n667), .A2(G85), .ZN(n668) );
  XNOR2_X1 U761 ( .A(n668), .B(KEYINPUT66), .ZN(n671) );
  NAND2_X1 U762 ( .A1(G72), .A2(n669), .ZN(n670) );
  NAND2_X1 U763 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U764 ( .A(KEYINPUT68), .B(n672), .Z(n676) );
  NAND2_X1 U765 ( .A1(G60), .A2(n681), .ZN(n674) );
  NAND2_X1 U766 ( .A1(G47), .A2(n677), .ZN(n673) );
  AND2_X1 U767 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U768 ( .A1(n676), .A2(n675), .ZN(G290) );
  NAND2_X1 U769 ( .A1(G49), .A2(n677), .ZN(n679) );
  NAND2_X1 U770 ( .A1(G74), .A2(G651), .ZN(n678) );
  NAND2_X1 U771 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U772 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U773 ( .A(n682), .B(KEYINPUT78), .ZN(n685) );
  NAND2_X1 U774 ( .A1(G87), .A2(n683), .ZN(n684) );
  NAND2_X1 U775 ( .A1(n685), .A2(n684), .ZN(G288) );
  NOR2_X1 U776 ( .A1(G868), .A2(n689), .ZN(n686) );
  XNOR2_X1 U777 ( .A(n686), .B(KEYINPUT83), .ZN(n699) );
  XNOR2_X1 U778 ( .A(KEYINPUT81), .B(KEYINPUT19), .ZN(n688) );
  XNOR2_X1 U779 ( .A(G305), .B(KEYINPUT80), .ZN(n687) );
  XNOR2_X1 U780 ( .A(n688), .B(n687), .ZN(n690) );
  XOR2_X1 U781 ( .A(n690), .B(n689), .Z(n692) );
  XNOR2_X1 U782 ( .A(n746), .B(G166), .ZN(n691) );
  XNOR2_X1 U783 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X1 U784 ( .A(n693), .B(G290), .ZN(n694) );
  XNOR2_X1 U785 ( .A(n694), .B(G288), .ZN(n918) );
  XNOR2_X1 U786 ( .A(n918), .B(KEYINPUT82), .ZN(n696) );
  XNOR2_X1 U787 ( .A(n696), .B(n695), .ZN(n697) );
  NAND2_X1 U788 ( .A1(G868), .A2(n697), .ZN(n698) );
  NAND2_X1 U789 ( .A1(n699), .A2(n698), .ZN(G295) );
  XOR2_X1 U790 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n701) );
  NAND2_X1 U791 ( .A1(G2084), .A2(G2078), .ZN(n700) );
  XNOR2_X1 U792 ( .A(n701), .B(n700), .ZN(n702) );
  NAND2_X1 U793 ( .A1(n702), .A2(G2090), .ZN(n703) );
  XOR2_X1 U794 ( .A(KEYINPUT21), .B(n703), .Z(n704) );
  XNOR2_X1 U795 ( .A(KEYINPUT85), .B(n704), .ZN(n705) );
  NAND2_X1 U796 ( .A1(n705), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U797 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U798 ( .A1(G132), .A2(G82), .ZN(n706) );
  XNOR2_X1 U799 ( .A(n706), .B(KEYINPUT86), .ZN(n707) );
  XNOR2_X1 U800 ( .A(n707), .B(KEYINPUT22), .ZN(n708) );
  NOR2_X1 U801 ( .A1(G218), .A2(n708), .ZN(n709) );
  NAND2_X1 U802 ( .A1(G96), .A2(n709), .ZN(n855) );
  NAND2_X1 U803 ( .A1(G2106), .A2(n855), .ZN(n713) );
  NAND2_X1 U804 ( .A1(G108), .A2(G120), .ZN(n710) );
  NOR2_X1 U805 ( .A1(G237), .A2(n710), .ZN(n711) );
  NAND2_X1 U806 ( .A1(G69), .A2(n711), .ZN(n856) );
  NAND2_X1 U807 ( .A1(G567), .A2(n856), .ZN(n712) );
  NAND2_X1 U808 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U809 ( .A(KEYINPUT87), .B(n714), .ZN(G319) );
  INV_X1 U810 ( .A(G319), .ZN(n716) );
  NAND2_X1 U811 ( .A1(G661), .A2(G483), .ZN(n715) );
  NOR2_X1 U812 ( .A1(n716), .A2(n715), .ZN(n854) );
  NAND2_X1 U813 ( .A1(n854), .A2(G36), .ZN(n717) );
  XNOR2_X1 U814 ( .A(KEYINPUT88), .B(n717), .ZN(G176) );
  INV_X1 U815 ( .A(G166), .ZN(G303) );
  AND2_X1 U816 ( .A1(G40), .A2(n718), .ZN(n720) );
  NAND2_X1 U817 ( .A1(G1341), .A2(n762), .ZN(n733) );
  AND2_X1 U818 ( .A1(n723), .A2(n733), .ZN(n726) );
  XOR2_X1 U819 ( .A(KEYINPUT26), .B(n724), .Z(n725) );
  XNOR2_X1 U820 ( .A(n728), .B(n727), .ZN(n732) );
  NOR2_X1 U821 ( .A1(n738), .A2(G1348), .ZN(n730) );
  NOR2_X1 U822 ( .A1(G2067), .A2(n762), .ZN(n729) );
  NOR2_X1 U823 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U824 ( .A1(n732), .A2(n731), .ZN(n737) );
  NAND2_X1 U825 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U826 ( .A1(n940), .A2(n735), .ZN(n736) );
  NAND2_X1 U827 ( .A1(n737), .A2(n736), .ZN(n745) );
  NAND2_X1 U828 ( .A1(G2072), .A2(n738), .ZN(n741) );
  INV_X1 U829 ( .A(G1956), .ZN(n969) );
  NOR2_X1 U830 ( .A1(n738), .A2(n969), .ZN(n742) );
  NOR2_X1 U831 ( .A1(n743), .A2(n742), .ZN(n747) );
  NAND2_X1 U832 ( .A1(n746), .A2(n747), .ZN(n744) );
  NOR2_X1 U833 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U834 ( .A(n748), .B(KEYINPUT28), .Z(n749) );
  XOR2_X1 U835 ( .A(G2078), .B(KEYINPUT25), .Z(n999) );
  NOR2_X1 U836 ( .A1(n999), .A2(n762), .ZN(n751) );
  XNOR2_X1 U837 ( .A(KEYINPUT94), .B(G1961), .ZN(n966) );
  NOR2_X1 U838 ( .A1(n738), .A2(n966), .ZN(n750) );
  NOR2_X1 U839 ( .A1(n751), .A2(n750), .ZN(n755) );
  NAND2_X1 U840 ( .A1(G8), .A2(n762), .ZN(n798) );
  NOR2_X1 U841 ( .A1(G1966), .A2(n798), .ZN(n774) );
  NOR2_X1 U842 ( .A1(G2084), .A2(n762), .ZN(n770) );
  NOR2_X1 U843 ( .A1(n774), .A2(n770), .ZN(n752) );
  NAND2_X1 U844 ( .A1(G8), .A2(n752), .ZN(n753) );
  XNOR2_X1 U845 ( .A(KEYINPUT30), .B(n753), .ZN(n754) );
  NOR2_X1 U846 ( .A1(G168), .A2(n754), .ZN(n757) );
  AND2_X1 U847 ( .A1(G301), .A2(n755), .ZN(n756) );
  NOR2_X1 U848 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U849 ( .A(n758), .B(KEYINPUT31), .ZN(n759) );
  XNOR2_X1 U850 ( .A(n761), .B(KEYINPUT97), .ZN(n772) );
  NAND2_X1 U851 ( .A1(n772), .A2(G286), .ZN(n767) );
  NOR2_X1 U852 ( .A1(G1971), .A2(n798), .ZN(n764) );
  NOR2_X1 U853 ( .A1(G2090), .A2(n762), .ZN(n763) );
  NOR2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U855 ( .A1(n765), .A2(G303), .ZN(n766) );
  NAND2_X1 U856 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U857 ( .A1(G8), .A2(n770), .ZN(n771) );
  NAND2_X1 U858 ( .A1(n772), .A2(n771), .ZN(n773) );
  OR2_X1 U859 ( .A1(G1976), .A2(G288), .ZN(n776) );
  INV_X1 U860 ( .A(G1971), .ZN(n978) );
  NAND2_X1 U861 ( .A1(G166), .A2(n978), .ZN(n775) );
  NAND2_X1 U862 ( .A1(n776), .A2(n775), .ZN(n961) );
  NAND2_X1 U863 ( .A1(G1976), .A2(G288), .ZN(n958) );
  INV_X1 U864 ( .A(KEYINPUT33), .ZN(n786) );
  OR2_X1 U865 ( .A1(n798), .A2(n776), .ZN(n777) );
  NOR2_X1 U866 ( .A1(n786), .A2(n777), .ZN(n778) );
  XNOR2_X1 U867 ( .A(n778), .B(KEYINPUT99), .ZN(n785) );
  AND2_X1 U868 ( .A1(n958), .A2(n785), .ZN(n781) );
  XNOR2_X1 U869 ( .A(G1981), .B(KEYINPUT100), .ZN(n779) );
  XNOR2_X1 U870 ( .A(n779), .B(G305), .ZN(n951) );
  INV_X1 U871 ( .A(n951), .ZN(n780) );
  AND2_X1 U872 ( .A1(n781), .A2(n780), .ZN(n783) );
  NAND2_X1 U873 ( .A1(n522), .A2(n784), .ZN(n790) );
  INV_X1 U874 ( .A(n785), .ZN(n787) );
  OR2_X1 U875 ( .A1(n787), .A2(n786), .ZN(n788) );
  OR2_X1 U876 ( .A1(n951), .A2(n788), .ZN(n789) );
  NAND2_X1 U877 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U878 ( .A(n791), .B(KEYINPUT101), .ZN(n803) );
  NOR2_X1 U879 ( .A1(G1981), .A2(G305), .ZN(n792) );
  XOR2_X1 U880 ( .A(n792), .B(KEYINPUT24), .Z(n793) );
  NOR2_X1 U881 ( .A1(n798), .A2(n793), .ZN(n801) );
  INV_X1 U882 ( .A(n794), .ZN(n797) );
  NOR2_X1 U883 ( .A1(G2090), .A2(G303), .ZN(n795) );
  NAND2_X1 U884 ( .A1(G8), .A2(n795), .ZN(n796) );
  NAND2_X1 U885 ( .A1(n797), .A2(n796), .ZN(n799) );
  AND2_X1 U886 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U887 ( .A1(n801), .A2(n800), .ZN(n802) );
  NOR2_X1 U888 ( .A1(n805), .A2(n804), .ZN(n846) );
  XNOR2_X1 U889 ( .A(KEYINPUT34), .B(KEYINPUT90), .ZN(n809) );
  NAND2_X1 U890 ( .A1(G104), .A2(n906), .ZN(n807) );
  NAND2_X1 U891 ( .A1(G140), .A2(n907), .ZN(n806) );
  NAND2_X1 U892 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U893 ( .A(n809), .B(n808), .ZN(n815) );
  NAND2_X1 U894 ( .A1(n902), .A2(G128), .ZN(n810) );
  XOR2_X1 U895 ( .A(KEYINPUT91), .B(n810), .Z(n812) );
  NAND2_X1 U896 ( .A1(G116), .A2(n903), .ZN(n811) );
  NAND2_X1 U897 ( .A1(n812), .A2(n811), .ZN(n813) );
  XOR2_X1 U898 ( .A(KEYINPUT35), .B(n813), .Z(n814) );
  NOR2_X1 U899 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U900 ( .A(n816), .B(KEYINPUT36), .ZN(n817) );
  XOR2_X1 U901 ( .A(n817), .B(KEYINPUT92), .Z(n887) );
  XOR2_X1 U902 ( .A(KEYINPUT37), .B(G2067), .Z(n843) );
  AND2_X1 U903 ( .A1(n887), .A2(n843), .ZN(n1024) );
  NAND2_X1 U904 ( .A1(n846), .A2(n1024), .ZN(n840) );
  NAND2_X1 U905 ( .A1(G105), .A2(n906), .ZN(n818) );
  XNOR2_X1 U906 ( .A(n818), .B(KEYINPUT38), .ZN(n825) );
  NAND2_X1 U907 ( .A1(G129), .A2(n902), .ZN(n820) );
  NAND2_X1 U908 ( .A1(G141), .A2(n907), .ZN(n819) );
  NAND2_X1 U909 ( .A1(n820), .A2(n819), .ZN(n823) );
  NAND2_X1 U910 ( .A1(G117), .A2(n903), .ZN(n821) );
  XNOR2_X1 U911 ( .A(KEYINPUT93), .B(n821), .ZN(n822) );
  NOR2_X1 U912 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U913 ( .A1(n825), .A2(n824), .ZN(n897) );
  AND2_X1 U914 ( .A1(n897), .A2(G1996), .ZN(n1020) );
  NAND2_X1 U915 ( .A1(G95), .A2(n906), .ZN(n827) );
  NAND2_X1 U916 ( .A1(G131), .A2(n907), .ZN(n826) );
  NAND2_X1 U917 ( .A1(n827), .A2(n826), .ZN(n831) );
  NAND2_X1 U918 ( .A1(G119), .A2(n902), .ZN(n829) );
  NAND2_X1 U919 ( .A1(G107), .A2(n903), .ZN(n828) );
  NAND2_X1 U920 ( .A1(n829), .A2(n828), .ZN(n830) );
  OR2_X1 U921 ( .A1(n831), .A2(n830), .ZN(n896) );
  AND2_X1 U922 ( .A1(n896), .A2(G1991), .ZN(n1018) );
  OR2_X1 U923 ( .A1(n1020), .A2(n1018), .ZN(n832) );
  NAND2_X1 U924 ( .A1(n846), .A2(n832), .ZN(n834) );
  NAND2_X1 U925 ( .A1(n840), .A2(n834), .ZN(n833) );
  XNOR2_X1 U926 ( .A(G1986), .B(G290), .ZN(n946) );
  NOR2_X1 U927 ( .A1(G1996), .A2(n897), .ZN(n1028) );
  INV_X1 U928 ( .A(n834), .ZN(n837) );
  NOR2_X1 U929 ( .A1(G1991), .A2(n896), .ZN(n1019) );
  NOR2_X1 U930 ( .A1(G1986), .A2(G290), .ZN(n835) );
  NOR2_X1 U931 ( .A1(n1019), .A2(n835), .ZN(n836) );
  NOR2_X1 U932 ( .A1(n837), .A2(n836), .ZN(n838) );
  NOR2_X1 U933 ( .A1(n1028), .A2(n838), .ZN(n839) );
  XNOR2_X1 U934 ( .A(n839), .B(KEYINPUT39), .ZN(n841) );
  NAND2_X1 U935 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U936 ( .A(n842), .B(KEYINPUT102), .ZN(n845) );
  NOR2_X1 U937 ( .A1(n887), .A2(n843), .ZN(n844) );
  XNOR2_X1 U938 ( .A(n844), .B(KEYINPUT103), .ZN(n1041) );
  NAND2_X1 U939 ( .A1(n845), .A2(n1041), .ZN(n847) );
  NAND2_X1 U940 ( .A1(n847), .A2(n846), .ZN(n848) );
  XNOR2_X1 U941 ( .A(KEYINPUT40), .B(KEYINPUT104), .ZN(n849) );
  XNOR2_X1 U942 ( .A(n850), .B(n849), .ZN(G329) );
  NAND2_X1 U943 ( .A1(G2106), .A2(n851), .ZN(G217) );
  AND2_X1 U944 ( .A1(G15), .A2(G2), .ZN(n852) );
  NAND2_X1 U945 ( .A1(G661), .A2(n852), .ZN(G259) );
  NAND2_X1 U946 ( .A1(G3), .A2(G1), .ZN(n853) );
  NAND2_X1 U947 ( .A1(n854), .A2(n853), .ZN(G188) );
  XOR2_X1 U948 ( .A(G120), .B(KEYINPUT106), .Z(G236) );
  INV_X1 U950 ( .A(G132), .ZN(G219) );
  INV_X1 U951 ( .A(G108), .ZN(G238) );
  INV_X1 U952 ( .A(G82), .ZN(G220) );
  NOR2_X1 U953 ( .A1(n856), .A2(n855), .ZN(G325) );
  INV_X1 U954 ( .A(G325), .ZN(G261) );
  XOR2_X1 U955 ( .A(KEYINPUT42), .B(G2090), .Z(n858) );
  XNOR2_X1 U956 ( .A(G2078), .B(G2084), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U958 ( .A(n859), .B(G2096), .Z(n861) );
  XNOR2_X1 U959 ( .A(G2067), .B(G2072), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U961 ( .A(KEYINPUT43), .B(KEYINPUT107), .Z(n863) );
  XNOR2_X1 U962 ( .A(G2678), .B(G2100), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U964 ( .A(n865), .B(n864), .Z(G227) );
  XNOR2_X1 U965 ( .A(G1981), .B(KEYINPUT41), .ZN(n875) );
  XOR2_X1 U966 ( .A(G1976), .B(G1971), .Z(n867) );
  XNOR2_X1 U967 ( .A(G1986), .B(G1956), .ZN(n866) );
  XNOR2_X1 U968 ( .A(n867), .B(n866), .ZN(n871) );
  XOR2_X1 U969 ( .A(G1961), .B(G1966), .Z(n869) );
  XNOR2_X1 U970 ( .A(G1996), .B(G1991), .ZN(n868) );
  XNOR2_X1 U971 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U972 ( .A(n871), .B(n870), .Z(n873) );
  XNOR2_X1 U973 ( .A(KEYINPUT108), .B(G2474), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n875), .B(n874), .ZN(G229) );
  NAND2_X1 U976 ( .A1(G100), .A2(n906), .ZN(n877) );
  NAND2_X1 U977 ( .A1(G112), .A2(n903), .ZN(n876) );
  NAND2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U979 ( .A(n878), .B(KEYINPUT109), .ZN(n880) );
  NAND2_X1 U980 ( .A1(G136), .A2(n907), .ZN(n879) );
  NAND2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n883) );
  NAND2_X1 U982 ( .A1(n902), .A2(G124), .ZN(n881) );
  XOR2_X1 U983 ( .A(KEYINPUT44), .B(n881), .Z(n882) );
  NOR2_X1 U984 ( .A1(n883), .A2(n882), .ZN(G162) );
  XOR2_X1 U985 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n885) );
  XNOR2_X1 U986 ( .A(G162), .B(n1017), .ZN(n884) );
  XNOR2_X1 U987 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U988 ( .A(n887), .B(n886), .Z(n901) );
  NAND2_X1 U989 ( .A1(G103), .A2(n906), .ZN(n889) );
  NAND2_X1 U990 ( .A1(G139), .A2(n907), .ZN(n888) );
  NAND2_X1 U991 ( .A1(n889), .A2(n888), .ZN(n895) );
  NAND2_X1 U992 ( .A1(G127), .A2(n902), .ZN(n891) );
  NAND2_X1 U993 ( .A1(G115), .A2(n903), .ZN(n890) );
  NAND2_X1 U994 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U995 ( .A(KEYINPUT47), .B(n892), .Z(n893) );
  XNOR2_X1 U996 ( .A(KEYINPUT110), .B(n893), .ZN(n894) );
  NOR2_X1 U997 ( .A1(n895), .A2(n894), .ZN(n1031) );
  XNOR2_X1 U998 ( .A(n1031), .B(n896), .ZN(n899) );
  XOR2_X1 U999 ( .A(G164), .B(n897), .Z(n898) );
  XNOR2_X1 U1000 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U1001 ( .A(n901), .B(n900), .ZN(n915) );
  NAND2_X1 U1002 ( .A1(G130), .A2(n902), .ZN(n905) );
  NAND2_X1 U1003 ( .A1(G118), .A2(n903), .ZN(n904) );
  NAND2_X1 U1004 ( .A1(n905), .A2(n904), .ZN(n912) );
  NAND2_X1 U1005 ( .A1(G106), .A2(n906), .ZN(n909) );
  NAND2_X1 U1006 ( .A1(G142), .A2(n907), .ZN(n908) );
  NAND2_X1 U1007 ( .A1(n909), .A2(n908), .ZN(n910) );
  XOR2_X1 U1008 ( .A(KEYINPUT45), .B(n910), .Z(n911) );
  NOR2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(G160), .B(n913), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(n915), .B(n914), .ZN(n916) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n916), .ZN(G395) );
  XNOR2_X1 U1013 ( .A(G171), .B(n942), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(KEYINPUT111), .B(n917), .ZN(n920) );
  XNOR2_X1 U1015 ( .A(n940), .B(n918), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(n920), .B(n919), .ZN(n921) );
  XOR2_X1 U1017 ( .A(n921), .B(G286), .Z(n922) );
  NOR2_X1 U1018 ( .A1(G37), .A2(n922), .ZN(n923) );
  XNOR2_X1 U1019 ( .A(KEYINPUT112), .B(n923), .ZN(G397) );
  XOR2_X1 U1020 ( .A(G2454), .B(G2435), .Z(n925) );
  XNOR2_X1 U1021 ( .A(G2438), .B(G2427), .ZN(n924) );
  XNOR2_X1 U1022 ( .A(n925), .B(n924), .ZN(n932) );
  XOR2_X1 U1023 ( .A(KEYINPUT105), .B(G2446), .Z(n927) );
  XNOR2_X1 U1024 ( .A(G2443), .B(G2430), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(n927), .B(n926), .ZN(n928) );
  XOR2_X1 U1026 ( .A(n928), .B(G2451), .Z(n930) );
  XNOR2_X1 U1027 ( .A(G1348), .B(G1341), .ZN(n929) );
  XNOR2_X1 U1028 ( .A(n930), .B(n929), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(n932), .B(n931), .ZN(n933) );
  NAND2_X1 U1030 ( .A1(n933), .A2(G14), .ZN(n939) );
  NAND2_X1 U1031 ( .A1(G319), .A2(n939), .ZN(n936) );
  NOR2_X1 U1032 ( .A1(G227), .A2(G229), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(KEYINPUT49), .B(n934), .ZN(n935) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(G395), .A2(G397), .ZN(n937) );
  NAND2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(G225) );
  INV_X1 U1037 ( .A(G225), .ZN(G308) );
  INV_X1 U1038 ( .A(G69), .ZN(G235) );
  INV_X1 U1039 ( .A(G96), .ZN(G221) );
  INV_X1 U1040 ( .A(n939), .ZN(G401) );
  XNOR2_X1 U1041 ( .A(G16), .B(KEYINPUT56), .ZN(n965) );
  XNOR2_X1 U1042 ( .A(G1348), .B(KEYINPUT122), .ZN(n941) );
  XNOR2_X1 U1043 ( .A(n941), .B(n940), .ZN(n944) );
  XNOR2_X1 U1044 ( .A(G1341), .B(n942), .ZN(n943) );
  NOR2_X1 U1045 ( .A1(n944), .A2(n943), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(G1961), .B(G301), .ZN(n945) );
  NOR2_X1 U1047 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1048 ( .A1(n948), .A2(n947), .ZN(n955) );
  XNOR2_X1 U1049 ( .A(KEYINPUT57), .B(KEYINPUT121), .ZN(n953) );
  XOR2_X1 U1050 ( .A(G1966), .B(KEYINPUT120), .Z(n949) );
  XNOR2_X1 U1051 ( .A(G168), .B(n949), .ZN(n950) );
  NOR2_X1 U1052 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1053 ( .A(n953), .B(n952), .Z(n954) );
  NOR2_X1 U1054 ( .A1(n955), .A2(n954), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(G299), .B(G1956), .ZN(n957) );
  NOR2_X1 U1056 ( .A1(n978), .A2(G166), .ZN(n956) );
  NOR2_X1 U1057 ( .A1(n957), .A2(n956), .ZN(n959) );
  NAND2_X1 U1058 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1059 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n1050) );
  XNOR2_X1 U1062 ( .A(G16), .B(KEYINPUT123), .ZN(n993) );
  XOR2_X1 U1063 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n991) );
  XNOR2_X1 U1064 ( .A(n966), .B(G5), .ZN(n968) );
  XNOR2_X1 U1065 ( .A(G21), .B(G1966), .ZN(n967) );
  NOR2_X1 U1066 ( .A1(n968), .A2(n967), .ZN(n989) );
  XNOR2_X1 U1067 ( .A(G20), .B(n969), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(G1341), .B(G19), .ZN(n971) );
  XNOR2_X1 U1069 ( .A(G1981), .B(G6), .ZN(n970) );
  NOR2_X1 U1070 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1071 ( .A1(n973), .A2(n972), .ZN(n976) );
  XOR2_X1 U1072 ( .A(KEYINPUT59), .B(G1348), .Z(n974) );
  XNOR2_X1 U1073 ( .A(G4), .B(n974), .ZN(n975) );
  NOR2_X1 U1074 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1075 ( .A(KEYINPUT60), .B(n977), .Z(n987) );
  XNOR2_X1 U1076 ( .A(G22), .B(n978), .ZN(n981) );
  XOR2_X1 U1077 ( .A(G1976), .B(KEYINPUT124), .Z(n979) );
  XNOR2_X1 U1078 ( .A(G23), .B(n979), .ZN(n980) );
  NAND2_X1 U1079 ( .A1(n981), .A2(n980), .ZN(n984) );
  XOR2_X1 U1080 ( .A(KEYINPUT125), .B(G1986), .Z(n982) );
  XNOR2_X1 U1081 ( .A(G24), .B(n982), .ZN(n983) );
  NOR2_X1 U1082 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1083 ( .A(KEYINPUT58), .B(n985), .Z(n986) );
  NOR2_X1 U1084 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1085 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1086 ( .A(n991), .B(n990), .ZN(n992) );
  NAND2_X1 U1087 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1088 ( .A1(n994), .A2(G11), .ZN(n1048) );
  XOR2_X1 U1089 ( .A(G34), .B(KEYINPUT118), .Z(n996) );
  XNOR2_X1 U1090 ( .A(G2084), .B(KEYINPUT54), .ZN(n995) );
  XNOR2_X1 U1091 ( .A(n996), .B(n995), .ZN(n1013) );
  XNOR2_X1 U1092 ( .A(G2090), .B(G35), .ZN(n1011) );
  XOR2_X1 U1093 ( .A(G1991), .B(G25), .Z(n997) );
  NAND2_X1 U1094 ( .A1(n997), .A2(G28), .ZN(n998) );
  XNOR2_X1 U1095 ( .A(n998), .B(KEYINPUT116), .ZN(n1008) );
  XOR2_X1 U1096 ( .A(G32), .B(G1996), .Z(n1006) );
  XNOR2_X1 U1097 ( .A(n999), .B(G27), .ZN(n1004) );
  XNOR2_X1 U1098 ( .A(G2067), .B(G26), .ZN(n1001) );
  XNOR2_X1 U1099 ( .A(G2072), .B(G33), .ZN(n1000) );
  NOR2_X1 U1100 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1101 ( .A(KEYINPUT117), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1102 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1103 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1104 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1105 ( .A(KEYINPUT53), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1106 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1107 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1108 ( .A(KEYINPUT119), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1109 ( .A1(G29), .A2(n1015), .ZN(n1016) );
  XNOR2_X1 U1110 ( .A(n1016), .B(KEYINPUT55), .ZN(n1046) );
  NOR2_X1 U1111 ( .A1(n1018), .A2(n1017), .ZN(n1026) );
  XNOR2_X1 U1112 ( .A(G160), .B(G2084), .ZN(n1022) );
  NOR2_X1 U1113 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1114 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1115 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1116 ( .A1(n1026), .A2(n1025), .ZN(n1040) );
  XOR2_X1 U1117 ( .A(G2090), .B(G162), .Z(n1027) );
  NOR2_X1 U1118 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1119 ( .A(KEYINPUT51), .B(n1029), .Z(n1030) );
  XOR2_X1 U1120 ( .A(KEYINPUT113), .B(n1030), .Z(n1038) );
  XNOR2_X1 U1121 ( .A(G2072), .B(n1031), .ZN(n1034) );
  XNOR2_X1 U1122 ( .A(G164), .B(G2078), .ZN(n1032) );
  XNOR2_X1 U1123 ( .A(n1032), .B(KEYINPUT114), .ZN(n1033) );
  NAND2_X1 U1124 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1125 ( .A(n1035), .B(KEYINPUT50), .ZN(n1036) );
  XNOR2_X1 U1126 ( .A(KEYINPUT115), .B(n1036), .ZN(n1037) );
  NAND2_X1 U1127 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NOR2_X1 U1128 ( .A1(n1040), .A2(n1039), .ZN(n1042) );
  NAND2_X1 U1129 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  XNOR2_X1 U1130 ( .A(KEYINPUT52), .B(n1043), .ZN(n1044) );
  NAND2_X1 U1131 ( .A1(G29), .A2(n1044), .ZN(n1045) );
  NAND2_X1 U1132 ( .A1(n1046), .A2(n1045), .ZN(n1047) );
  NOR2_X1 U1133 ( .A1(n1048), .A2(n1047), .ZN(n1049) );
  NAND2_X1 U1134 ( .A1(n1050), .A2(n1049), .ZN(n1051) );
  XNOR2_X1 U1135 ( .A(n1051), .B(KEYINPUT62), .ZN(n1052) );
  XNOR2_X1 U1136 ( .A(KEYINPUT127), .B(n1052), .ZN(G311) );
  INV_X1 U1137 ( .A(G311), .ZN(G150) );
endmodule

