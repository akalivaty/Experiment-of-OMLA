//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1250, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309;
  OR3_X1    g0000(.A1(KEYINPUT64), .A2(G58), .A3(G68), .ZN(new_n201));
  OAI21_X1  g0001(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n202));
  AOI21_X1  g0002(.A(G50), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g0003(.A(G77), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT65), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n208), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n217), .A2(KEYINPUT0), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n201), .A2(new_n202), .ZN(new_n219));
  INV_X1    g0019(.A(G50), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n222), .A2(new_n210), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n217), .A2(KEYINPUT0), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n218), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT66), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n228));
  INV_X1    g0028(.A(G68), .ZN(new_n229));
  INV_X1    g0029(.A(G238), .ZN(new_n230));
  INV_X1    g0030(.A(G87), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n228), .B1(new_n229), .B2(new_n230), .C1(new_n231), .C2(new_n208), .ZN(new_n232));
  AOI22_X1  g0032(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n233));
  INV_X1    g0033(.A(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G107), .ZN(new_n235));
  OAI221_X1 g0035(.A(new_n233), .B1(new_n204), .B2(new_n234), .C1(new_n235), .C2(new_n216), .ZN(new_n236));
  OAI21_X1  g0036(.A(new_n212), .B1(new_n232), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT1), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n227), .A2(new_n238), .ZN(G361));
  XOR2_X1   g0039(.A(G238), .B(G244), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT2), .B(G226), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G250), .B(G257), .Z(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(KEYINPUT67), .B(KEYINPUT68), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n243), .B(new_n248), .ZN(G358));
  XNOR2_X1  g0049(.A(G68), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT69), .ZN(new_n251));
  XOR2_X1   g0051(.A(G50), .B(G58), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(G97), .B(G107), .Z(new_n254));
  XNOR2_X1  g0054(.A(G87), .B(G116), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XOR2_X1   g0056(.A(new_n253), .B(new_n256), .Z(G351));
  XNOR2_X1  g0057(.A(KEYINPUT8), .B(G58), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G20), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n259), .A2(new_n261), .B1(G150), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n263), .B1(new_n203), .B2(new_n210), .ZN(new_n264));
  NAND3_X1  g0064(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n222), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n266), .B(KEYINPUT73), .ZN(new_n267));
  INV_X1    g0067(.A(G13), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n268), .A2(new_n210), .A3(G1), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n264), .A2(new_n267), .B1(new_n220), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n267), .A2(new_n269), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n210), .A2(G1), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(G50), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT71), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT71), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G1698), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT70), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n286), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT70), .B1(new_n288), .B2(new_n283), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n282), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G222), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n287), .A2(new_n289), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n278), .B1(new_n287), .B2(new_n289), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G223), .ZN(new_n295));
  OAI221_X1 g0095(.A(new_n291), .B1(new_n204), .B2(new_n292), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n277), .B1(new_n296), .B2(KEYINPUT72), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(KEYINPUT72), .B2(new_n296), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n277), .A2(G274), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n277), .A2(new_n300), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n301), .B1(G226), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n298), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n275), .B1(new_n306), .B2(G169), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n305), .A2(G179), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n275), .B(KEYINPUT9), .ZN(new_n310));
  INV_X1    g0110(.A(G200), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n310), .B1(new_n306), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G190), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n305), .A2(new_n313), .ZN(new_n314));
  OR3_X1    g0114(.A1(new_n312), .A2(KEYINPUT10), .A3(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT10), .B1(new_n312), .B2(new_n314), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n309), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n301), .B1(G232), .B2(new_n303), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT80), .ZN(new_n319));
  OR2_X1    g0119(.A1(KEYINPUT79), .A2(G33), .ZN(new_n320));
  NAND2_X1  g0120(.A1(KEYINPUT79), .A2(G33), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(KEYINPUT3), .A3(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n319), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  AND2_X1   g0125(.A1(KEYINPUT79), .A2(G33), .ZN(new_n326));
  NOR2_X1   g0126(.A1(KEYINPUT79), .A2(G33), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT80), .B1(new_n328), .B2(KEYINPUT3), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G226), .A2(G1698), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n282), .B2(new_n295), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n330), .A2(new_n332), .B1(G33), .B2(G87), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n318), .B1(new_n333), .B2(new_n277), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G169), .ZN(new_n335));
  INV_X1    g0135(.A(G179), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n335), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G58), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n338), .A2(new_n229), .ZN(new_n339));
  OAI21_X1  g0139(.A(G20), .B1(new_n219), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n262), .A2(G159), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT7), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n343), .A2(G20), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n286), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT3), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n345), .B1(new_n328), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n287), .A2(new_n289), .A3(new_n210), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n347), .B1(new_n348), .B2(new_n343), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n342), .B1(new_n349), .B2(new_n229), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT16), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n266), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n210), .B1(new_n325), .B2(new_n329), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n354), .A2(KEYINPUT81), .A3(new_n343), .ZN(new_n355));
  INV_X1    g0155(.A(new_n344), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT82), .B1(new_n330), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT82), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n358), .B(new_n344), .C1(new_n325), .C2(new_n329), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n355), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT81), .B1(new_n354), .B2(new_n343), .ZN(new_n361));
  OAI21_X1  g0161(.A(G68), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n342), .A2(KEYINPUT16), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n353), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n258), .A2(new_n272), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n366), .B(KEYINPUT83), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n367), .A2(new_n271), .B1(new_n269), .B2(new_n258), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n337), .B1(new_n365), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT18), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n334), .A2(new_n311), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(G190), .B2(new_n334), .ZN(new_n373));
  INV_X1    g0173(.A(new_n361), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n374), .A2(new_n355), .A3(new_n357), .A4(new_n359), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n363), .B1(new_n375), .B2(G68), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n373), .B(new_n368), .C1(new_n376), .C2(new_n353), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT17), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n362), .A2(new_n364), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n380), .A2(new_n266), .A3(new_n352), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n381), .A2(KEYINPUT17), .A3(new_n368), .A4(new_n373), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT18), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n337), .B(new_n383), .C1(new_n365), .C2(new_n369), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n371), .A2(new_n379), .A3(new_n382), .A4(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n261), .A2(G77), .B1(G20), .B2(new_n229), .ZN(new_n387));
  INV_X1    g0187(.A(new_n262), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n387), .B1(new_n220), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n267), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT11), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n268), .A2(G1), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(G20), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT75), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n269), .A2(KEYINPUT75), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n266), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n272), .A2(new_n229), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n390), .A2(new_n391), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n267), .A2(new_n389), .A3(KEYINPUT11), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n395), .A2(new_n396), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT12), .B1(new_n401), .B2(G68), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT12), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n392), .A2(new_n403), .A3(G20), .A4(new_n229), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n399), .A2(new_n400), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT77), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n399), .A2(new_n405), .A3(KEYINPUT77), .A4(new_n400), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n290), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n292), .A2(G232), .A3(G1698), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n277), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n301), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(new_n302), .B2(new_n230), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT13), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n290), .A2(G226), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G33), .A2(G97), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(new_n412), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n276), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT13), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n301), .B1(G238), .B2(new_n303), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n416), .A2(new_n423), .A3(G190), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n410), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n311), .B1(new_n416), .B2(new_n423), .ZN(new_n426));
  OAI21_X1  g0226(.A(KEYINPUT78), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n426), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT78), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n428), .A2(new_n429), .A3(new_n410), .A4(new_n424), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT14), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n416), .A2(new_n423), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n432), .B1(new_n433), .B2(G169), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n416), .A2(new_n423), .A3(G179), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n433), .A2(new_n432), .A3(G169), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n410), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  XOR2_X1   g0240(.A(KEYINPUT15), .B(G87), .Z(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n261), .ZN(new_n442));
  OAI221_X1 g0242(.A(new_n442), .B1(new_n210), .B2(new_n204), .C1(new_n388), .C2(new_n258), .ZN(new_n443));
  INV_X1    g0243(.A(new_n401), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n443), .A2(new_n266), .B1(new_n204), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n397), .A2(G77), .A3(new_n273), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n414), .B1(new_n302), .B2(new_n234), .ZN(new_n448));
  INV_X1    g0248(.A(new_n282), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n292), .A2(G232), .A3(new_n449), .ZN(new_n450));
  XOR2_X1   g0250(.A(KEYINPUT74), .B(G107), .Z(new_n451));
  OAI221_X1 g0251(.A(new_n450), .B1(new_n292), .B2(new_n451), .C1(new_n294), .C2(new_n230), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n448), .B1(new_n452), .B2(new_n276), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n447), .B1(new_n453), .B2(new_n311), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT76), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT76), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n447), .B(new_n456), .C1(new_n453), .C2(new_n311), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n453), .A2(G190), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n455), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n453), .A2(new_n336), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n445), .A2(new_n446), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(new_n453), .B2(G169), .ZN(new_n462));
  OR2_X1    g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n440), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n317), .A2(new_n386), .A3(new_n431), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n269), .A2(new_n235), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n467), .B(KEYINPUT25), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT73), .ZN(new_n469));
  XNOR2_X1  g0269(.A(new_n266), .B(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n209), .A2(G33), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n470), .A2(new_n393), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n468), .B1(new_n473), .B2(G107), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT5), .ZN(new_n475));
  OR3_X1    g0275(.A1(new_n475), .A2(KEYINPUT85), .A3(G41), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n475), .B1(KEYINPUT85), .B2(G41), .ZN(new_n477));
  INV_X1    g0277(.A(G45), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(G1), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n476), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  OR2_X1    g0280(.A1(new_n299), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n277), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n481), .B1(new_n216), .B2(new_n482), .ZN(new_n483));
  OAI22_X1  g0283(.A1(new_n282), .A2(new_n208), .B1(new_n215), .B2(new_n278), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n330), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n328), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G294), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n483), .B1(new_n488), .B2(new_n276), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n313), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n490), .B1(G200), .B2(new_n489), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT94), .ZN(new_n492));
  XOR2_X1   g0292(.A(KEYINPUT92), .B(KEYINPUT24), .Z(new_n493));
  INV_X1    g0293(.A(new_n292), .ZN(new_n494));
  NOR4_X1   g0294(.A1(new_n494), .A2(KEYINPUT22), .A3(G20), .A4(new_n231), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT22), .ZN(new_n496));
  NOR4_X1   g0296(.A1(new_n325), .A2(new_n329), .A3(G20), .A4(new_n231), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT91), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n326), .A2(new_n327), .A3(new_n346), .ZN(new_n500));
  OAI21_X1  g0300(.A(KEYINPUT80), .B1(new_n500), .B2(new_n323), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n322), .A2(new_n319), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n501), .A2(new_n210), .A3(G87), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT91), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n495), .B1(new_n499), .B2(new_n504), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n210), .A2(KEYINPUT23), .A3(G107), .ZN(new_n506));
  XOR2_X1   g0306(.A(new_n506), .B(KEYINPUT93), .Z(new_n507));
  INV_X1    g0307(.A(new_n451), .ZN(new_n508));
  OAI21_X1  g0308(.A(KEYINPUT23), .B1(new_n508), .B2(new_n210), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n486), .A2(new_n210), .A3(G116), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n507), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n493), .B1(new_n505), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n495), .ZN(new_n513));
  OAI21_X1  g0313(.A(KEYINPUT22), .B1(new_n503), .B2(KEYINPUT91), .ZN(new_n514));
  NOR3_X1   g0314(.A1(new_n325), .A2(new_n329), .A3(G20), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n498), .B1(new_n515), .B2(G87), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n513), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n511), .ZN(new_n518));
  INV_X1    g0318(.A(new_n493), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n512), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n492), .B1(new_n521), .B2(new_n266), .ZN(new_n522));
  INV_X1    g0322(.A(new_n266), .ZN(new_n523));
  AOI211_X1 g0323(.A(KEYINPUT94), .B(new_n523), .C1(new_n512), .C2(new_n520), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n474), .B(new_n491), .C1(new_n522), .C2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n474), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n515), .A2(new_n498), .A3(G87), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n527), .A2(new_n504), .A3(KEYINPUT22), .ZN(new_n528));
  AOI211_X1 g0328(.A(new_n511), .B(new_n493), .C1(new_n528), .C2(new_n513), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n519), .B1(new_n517), .B2(new_n518), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n266), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT94), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n492), .B(new_n266), .C1(new_n529), .C2(new_n530), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n526), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n489), .A2(new_n336), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(G169), .B2(new_n489), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n525), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(G169), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n482), .A2(new_n215), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n282), .A2(new_n234), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n501), .A2(new_n502), .A3(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT4), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n292), .A2(KEYINPUT4), .A3(G244), .A4(new_n449), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n293), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n539), .B1(new_n546), .B2(new_n276), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n538), .B1(new_n547), .B2(new_n481), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n292), .A2(G250), .A3(G1698), .ZN(new_n549));
  NAND2_X1  g0349(.A1(G33), .A2(G283), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n544), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n277), .B1(new_n551), .B2(new_n543), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n299), .A2(new_n480), .ZN(new_n553));
  NOR4_X1   g0353(.A1(new_n552), .A2(new_n336), .A3(new_n553), .A4(new_n539), .ZN(new_n554));
  INV_X1    g0354(.A(G97), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n269), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n472), .B2(new_n555), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT84), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT6), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n559), .A2(new_n555), .A3(G107), .ZN(new_n560));
  XNOR2_X1  g0360(.A(G97), .B(G107), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n560), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  OAI221_X1 g0362(.A(new_n558), .B1(new_n204), .B2(new_n388), .C1(new_n562), .C2(new_n210), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n559), .ZN(new_n564));
  INV_X1    g0364(.A(new_n560), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n210), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n388), .A2(new_n204), .ZN(new_n567));
  OAI21_X1  g0367(.A(KEYINPUT84), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n563), .B(new_n568), .C1(new_n451), .C2(new_n349), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n557), .B1(new_n569), .B2(new_n266), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT86), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI211_X1 g0372(.A(KEYINPUT86), .B(new_n557), .C1(new_n569), .C2(new_n266), .ZN(new_n573));
  OAI22_X1  g0373(.A1(new_n548), .A2(new_n554), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT88), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n401), .A2(new_n441), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n501), .A2(new_n210), .A3(G68), .A4(new_n502), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT19), .B1(new_n261), .B2(G97), .ZN(new_n579));
  XNOR2_X1  g0379(.A(KEYINPUT87), .B(G87), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n451), .A2(new_n555), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT19), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(new_n418), .B2(new_n210), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n579), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n575), .B(new_n577), .C1(new_n585), .C2(new_n523), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n523), .B1(new_n578), .B2(new_n584), .ZN(new_n587));
  OAI21_X1  g0387(.A(KEYINPUT88), .B1(new_n587), .B2(new_n576), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n473), .A2(new_n441), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI22_X1  g0391(.A1(new_n282), .A2(new_n230), .B1(new_n234), .B2(new_n278), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n501), .A2(new_n502), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n486), .A2(G116), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n277), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n479), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n277), .A2(G250), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n299), .B2(new_n596), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n538), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n336), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n591), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n547), .A2(G190), .A3(new_n481), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n552), .A2(new_n553), .A3(new_n539), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n604), .B(new_n570), .C1(new_n605), .C2(new_n311), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n600), .A2(G200), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n473), .A2(G87), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n599), .A2(G190), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n589), .A2(new_n607), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n574), .A2(new_n603), .A3(new_n606), .A4(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT90), .ZN(new_n612));
  INV_X1    g0412(.A(new_n482), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n553), .B1(G270), .B2(new_n613), .ZN(new_n614));
  OAI22_X1  g0414(.A1(new_n282), .A2(new_n215), .B1(new_n216), .B2(new_n278), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n330), .A2(new_n615), .B1(G303), .B2(new_n494), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n614), .B1(new_n616), .B2(new_n277), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G169), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n397), .A2(G116), .A3(new_n471), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(G116), .B2(new_n401), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n266), .B1(new_n210), .B2(G116), .ZN(new_n621));
  XNOR2_X1  g0421(.A(new_n621), .B(KEYINPUT89), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n550), .B(new_n210), .C1(G33), .C2(new_n555), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT20), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n622), .A2(KEYINPUT20), .A3(new_n623), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n620), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n612), .B1(new_n618), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT21), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT21), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n612), .B(new_n631), .C1(new_n618), .C2(new_n628), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n614), .B(G179), .C1(new_n616), .C2(new_n277), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n617), .A2(G200), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n635), .B(new_n628), .C1(new_n313), .C2(new_n617), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n630), .A2(new_n632), .A3(new_n634), .A4(new_n636), .ZN(new_n637));
  NOR4_X1   g0437(.A1(new_n466), .A2(new_n537), .A3(new_n611), .A4(new_n637), .ZN(G372));
  NAND2_X1  g0438(.A1(new_n603), .A2(new_n610), .ZN(new_n639));
  OAI21_X1  g0439(.A(KEYINPUT26), .B1(new_n639), .B2(new_n574), .ZN(new_n640));
  INV_X1    g0440(.A(new_n548), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n605), .A2(G179), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n570), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT26), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n643), .A2(new_n644), .A3(new_n603), .A4(new_n610), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n640), .A2(new_n603), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n630), .A2(new_n632), .A3(new_n634), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n648), .B1(new_n534), .B2(new_n536), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n611), .B1(new_n534), .B2(new_n491), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n646), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n466), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n652), .B(KEYINPUT95), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n371), .A2(new_n384), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n379), .A2(new_n382), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n463), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n428), .A2(new_n410), .A3(new_n424), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n438), .A2(new_n439), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n654), .B1(new_n656), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n315), .A2(new_n316), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n309), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n653), .A2(new_n662), .ZN(G369));
  OAI21_X1  g0463(.A(new_n474), .B1(new_n522), .B2(new_n524), .ZN(new_n664));
  INV_X1    g0464(.A(new_n536), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n392), .A2(new_n210), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G213), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g0470(.A(KEYINPUT96), .B(G343), .Z(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n664), .A2(new_n665), .A3(new_n672), .ZN(new_n674));
  INV_X1    g0474(.A(new_n672), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n534), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n674), .B1(new_n537), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(KEYINPUT97), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT97), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n679), .B(new_n674), .C1(new_n537), .C2(new_n676), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n647), .A2(new_n675), .ZN(new_n682));
  XOR2_X1   g0482(.A(new_n682), .B(KEYINPUT98), .Z(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n673), .B1(new_n681), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n628), .A2(new_n675), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n647), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n637), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G330), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n681), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n685), .A2(new_n691), .ZN(G399));
  NOR2_X1   g0492(.A1(new_n214), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G1), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n581), .A2(G116), .ZN(new_n696));
  INV_X1    g0496(.A(new_n221), .ZN(new_n697));
  OAI22_X1  g0497(.A1(new_n695), .A2(new_n696), .B1(new_n697), .B2(new_n694), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n603), .B(KEYINPUT100), .Z(new_n700));
  AND2_X1   g0500(.A1(new_n603), .A2(new_n610), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n644), .B1(new_n701), .B2(new_n643), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n639), .A2(KEYINPUT26), .A3(new_n574), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n700), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n649), .A2(new_n650), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n672), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT29), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n611), .A2(new_n637), .A3(new_n672), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n666), .A2(new_n709), .A3(new_n525), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT99), .ZN(new_n711));
  AOI21_X1  g0511(.A(KEYINPUT4), .B1(new_n330), .B2(new_n540), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n544), .A2(new_n550), .A3(new_n549), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n276), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n539), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n489), .A2(new_n714), .A3(new_n715), .A4(new_n599), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n711), .B1(new_n716), .B2(new_n633), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(KEYINPUT30), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n711), .B(new_n719), .C1(new_n716), .C2(new_n633), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n547), .A2(new_n481), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n489), .A2(G179), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n721), .A2(new_n722), .A3(new_n600), .A4(new_n617), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n718), .A2(new_n720), .A3(new_n723), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n672), .ZN(new_n725));
  AOI21_X1  g0525(.A(KEYINPUT31), .B1(new_n724), .B2(new_n672), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n710), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G330), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n651), .A2(KEYINPUT29), .A3(new_n672), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n708), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n699), .B1(new_n732), .B2(G1), .ZN(G364));
  NOR2_X1   g0533(.A1(new_n268), .A2(G20), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n209), .B1(new_n734), .B2(G45), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n693), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n690), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(G330), .B2(new_n688), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n210), .A2(new_n336), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n311), .A2(G190), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G190), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  OAI22_X1  g0544(.A1(new_n229), .A2(new_n742), .B1(new_n744), .B2(new_n204), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n313), .A2(G179), .A3(G200), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n210), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n740), .A2(G190), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n311), .ZN(new_n750));
  AOI22_X1  g0550(.A1(G97), .A2(new_n748), .B1(new_n750), .B2(G50), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT32), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n210), .A2(G179), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n743), .ZN(new_n754));
  INV_X1    g0554(.A(G159), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n749), .A2(G200), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n751), .B1(new_n752), .B2(new_n756), .C1(new_n338), .C2(new_n758), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n745), .B(new_n759), .C1(new_n752), .C2(new_n756), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n753), .A2(new_n741), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n753), .A2(G190), .A3(G200), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n292), .B1(new_n235), .B2(new_n761), .C1(new_n580), .C2(new_n762), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT104), .ZN(new_n764));
  INV_X1    g0564(.A(new_n750), .ZN(new_n765));
  INV_X1    g0565(.A(G326), .ZN(new_n766));
  INV_X1    g0566(.A(G294), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n765), .A2(new_n766), .B1(new_n767), .B2(new_n747), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n292), .B(new_n768), .C1(G322), .C2(new_n757), .ZN(new_n769));
  INV_X1    g0569(.A(new_n762), .ZN(new_n770));
  INV_X1    g0570(.A(new_n754), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n770), .A2(G303), .B1(new_n771), .B2(G329), .ZN(new_n772));
  INV_X1    g0572(.A(G283), .ZN(new_n773));
  INV_X1    g0573(.A(G311), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n772), .B1(new_n773), .B2(new_n761), .C1(new_n774), .C2(new_n744), .ZN(new_n775));
  XNOR2_X1  g0575(.A(KEYINPUT33), .B(G317), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(KEYINPUT105), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n776), .A2(KEYINPUT105), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n742), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n775), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n760), .A2(new_n764), .B1(new_n769), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n222), .B1(G20), .B2(new_n538), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n737), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n268), .A2(new_n260), .A3(KEYINPUT103), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT103), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(G13), .B2(G33), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n494), .A2(new_n214), .ZN(new_n791));
  INV_X1    g0591(.A(G116), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n791), .A2(G355), .B1(new_n792), .B2(new_n214), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n253), .A2(G45), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT101), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n330), .A2(new_n214), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(G45), .B2(new_n697), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n793), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n790), .B(new_n782), .C1(new_n798), .C2(KEYINPUT102), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n798), .A2(KEYINPUT102), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n784), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n790), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n688), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n739), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(G396));
  NOR2_X1   g0605(.A1(new_n463), .A2(new_n672), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n459), .B1(new_n447), .B2(new_n675), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n806), .B1(new_n807), .B2(new_n463), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n651), .B2(new_n672), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n464), .A2(new_n675), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n810), .B1(new_n651), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n737), .B1(new_n812), .B2(new_n729), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n729), .B2(new_n812), .ZN(new_n814));
  INV_X1    g0614(.A(new_n737), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n788), .A2(new_n782), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n815), .B1(new_n204), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n742), .ZN(new_n818));
  INV_X1    g0618(.A(new_n744), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G150), .A2(new_n818), .B1(new_n819), .B2(G159), .ZN(new_n820));
  INV_X1    g0620(.A(G143), .ZN(new_n821));
  INV_X1    g0621(.A(G137), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n820), .B1(new_n758), .B2(new_n821), .C1(new_n822), .C2(new_n765), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT34), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n330), .ZN(new_n826));
  INV_X1    g0626(.A(new_n761), .ZN(new_n827));
  AOI22_X1  g0627(.A1(G68), .A2(new_n827), .B1(new_n771), .B2(G132), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n828), .B1(new_n220), .B2(new_n762), .C1(new_n338), .C2(new_n747), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n825), .A2(new_n826), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n823), .A2(new_n824), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(G303), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n767), .A2(new_n758), .B1(new_n765), .B2(new_n833), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n292), .B(new_n834), .C1(G97), .C2(new_n748), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G107), .A2(new_n770), .B1(new_n818), .B2(G283), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n792), .B2(new_n744), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT106), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n761), .A2(new_n231), .B1(new_n754), .B2(new_n774), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n835), .B(new_n840), .C1(new_n838), .C2(new_n839), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n832), .A2(new_n841), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n817), .B1(new_n783), .B2(new_n842), .C1(new_n808), .C2(new_n789), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n814), .A2(new_n843), .ZN(G384));
  NOR2_X1   g0644(.A1(new_n734), .A2(new_n209), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT110), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT109), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n439), .A2(new_n672), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n437), .A2(new_n436), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n849), .A2(new_n434), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n848), .B1(new_n431), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n848), .B1(new_n425), .B2(new_n426), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(new_n438), .B2(new_n439), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n808), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n847), .B(new_n854), .C1(new_n710), .C2(new_n727), .ZN(new_n855));
  INV_X1    g0655(.A(new_n854), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT109), .B1(new_n728), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT40), .ZN(new_n859));
  INV_X1    g0659(.A(new_n670), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n365), .B2(new_n369), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n370), .A2(new_n861), .A3(new_n377), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT37), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT37), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n370), .A2(new_n861), .A3(new_n377), .A4(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n863), .A2(KEYINPUT108), .A3(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n861), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n385), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT108), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n862), .A2(new_n869), .A3(KEYINPUT37), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n866), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n362), .A2(new_n342), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n351), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n470), .B1(new_n362), .B2(new_n364), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n369), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n337), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n377), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n877), .A2(new_n670), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT37), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n865), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n385), .A2(new_n880), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n882), .A2(KEYINPUT38), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n859), .B1(new_n873), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n846), .B1(new_n858), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n728), .A2(new_n856), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n847), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n854), .B1(new_n710), .B2(new_n727), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT109), .ZN(new_n890));
  AND4_X1   g0690(.A1(new_n846), .A2(new_n888), .A3(new_n885), .A4(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n886), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n865), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n380), .A2(new_n267), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT16), .B1(new_n362), .B2(new_n342), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n368), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n860), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n337), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n897), .A2(new_n898), .A3(new_n377), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n893), .B1(new_n899), .B2(KEYINPUT37), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n897), .B1(new_n654), .B2(new_n655), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n872), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n902), .A2(new_n884), .A3(KEYINPUT107), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT107), .B1(new_n902), .B2(new_n884), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n889), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n892), .B1(new_n859), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n466), .B1(new_n710), .B2(new_n727), .ZN(new_n907));
  OAI21_X1  g0707(.A(G330), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n908), .A2(KEYINPUT111), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(KEYINPUT111), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n906), .A2(new_n907), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n902), .A2(new_n884), .A3(KEYINPUT39), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT39), .B1(new_n873), .B2(new_n884), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n438), .A2(new_n439), .A3(new_n675), .ZN(new_n915));
  OR3_X1    g0715(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n806), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n651), .B2(new_n811), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n851), .A2(new_n853), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n918), .B(new_n920), .C1(new_n903), .C2(new_n904), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n654), .A2(new_n860), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n916), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n466), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n708), .B2(new_n731), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n662), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n923), .B(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n845), .B1(new_n912), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n927), .B2(new_n912), .ZN(new_n929));
  INV_X1    g0729(.A(new_n562), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n930), .A2(KEYINPUT35), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(KEYINPUT35), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n931), .A2(G116), .A3(new_n223), .A4(new_n932), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n933), .B(KEYINPUT36), .Z(new_n934));
  OAI211_X1 g0734(.A(new_n221), .B(G77), .C1(new_n338), .C2(new_n229), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n220), .A2(G68), .ZN(new_n936));
  AOI211_X1 g0736(.A(new_n209), .B(G13), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n929), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n939), .B(KEYINPUT112), .Z(G367));
  NOR2_X1   g0740(.A1(new_n790), .A2(new_n782), .ZN(new_n941));
  INV_X1    g0741(.A(new_n441), .ZN(new_n942));
  INV_X1    g0742(.A(new_n796), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n941), .B1(new_n213), .B2(new_n942), .C1(new_n248), .C2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n747), .A2(new_n229), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n765), .A2(new_n821), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n945), .B(new_n946), .C1(G150), .C2(new_n757), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n338), .A2(new_n762), .B1(new_n742), .B2(new_n755), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(G137), .B2(new_n771), .ZN(new_n949));
  AOI22_X1  g0749(.A1(G50), .A2(new_n819), .B1(new_n827), .B2(G77), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n947), .A2(new_n292), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  XOR2_X1   g0751(.A(KEYINPUT114), .B(G311), .Z(new_n952));
  NAND2_X1  g0752(.A1(new_n750), .A2(new_n952), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n953), .B1(new_n451), .B2(new_n747), .C1(new_n758), .C2(new_n833), .ZN(new_n954));
  AOI22_X1  g0754(.A1(G283), .A2(new_n819), .B1(new_n771), .B2(G317), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n555), .B2(new_n761), .ZN(new_n956));
  OR3_X1    g0756(.A1(new_n954), .A2(new_n330), .A3(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n770), .A2(KEYINPUT46), .A3(G116), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT46), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n762), .B2(new_n792), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n958), .B(new_n960), .C1(new_n767), .C2(new_n742), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT115), .Z(new_n962));
  OAI21_X1  g0762(.A(new_n951), .B1(new_n957), .B2(new_n962), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT47), .Z(new_n964));
  OAI211_X1 g0764(.A(new_n737), .B(new_n944), .C1(new_n964), .C2(new_n783), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT116), .Z(new_n966));
  AOI21_X1  g0766(.A(new_n675), .B1(new_n589), .B2(new_n608), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n967), .A2(new_n591), .A3(new_n601), .A4(new_n602), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n639), .B2(new_n967), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n790), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n966), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n735), .B(KEYINPUT113), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n680), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n664), .A2(new_n672), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n666), .A2(new_n976), .A3(new_n525), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n679), .B1(new_n977), .B2(new_n674), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n684), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n673), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n574), .B(new_n606), .C1(new_n570), .C2(new_n675), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n643), .A2(new_n672), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(KEYINPUT44), .B1(new_n981), .B2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT44), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n987), .B(new_n984), .C1(new_n979), .C2(new_n980), .ZN(new_n988));
  AOI21_X1  g0788(.A(KEYINPUT45), .B1(new_n685), .B2(new_n984), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n683), .B1(new_n678), .B2(new_n680), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT45), .ZN(new_n991));
  NOR4_X1   g0791(.A1(new_n990), .A2(new_n991), .A3(new_n673), .A4(new_n985), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n986), .A2(new_n988), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n691), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n987), .B1(new_n685), .B2(new_n984), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n981), .A2(KEYINPUT44), .A3(new_n985), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n979), .A2(new_n980), .A3(new_n984), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n991), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n979), .A2(KEYINPUT45), .A3(new_n980), .A4(new_n984), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n998), .A2(new_n1002), .A3(new_n691), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n678), .A2(new_n680), .A3(new_n683), .ZN(new_n1004));
  AND3_X1   g0804(.A1(new_n979), .A2(new_n690), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n690), .B1(new_n979), .B2(new_n1004), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n732), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n995), .A2(new_n1003), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n732), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n693), .B(KEYINPUT41), .Z(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n974), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT43), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n970), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n970), .A2(new_n1015), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n990), .A2(new_n984), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1019), .A2(KEYINPUT42), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n574), .B1(new_n985), .B2(new_n666), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1019), .A2(KEYINPUT42), .B1(new_n675), .B2(new_n1021), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1017), .B(new_n1018), .C1(new_n1020), .C2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1020), .A2(new_n1022), .A3(new_n1015), .A4(new_n970), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n1023), .A2(new_n1025), .B1(new_n691), .B2(new_n985), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1018), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n1016), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1028), .A2(new_n994), .A3(new_n984), .A4(new_n1024), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n972), .B1(new_n1014), .B2(new_n1030), .ZN(G387));
  INV_X1    g0831(.A(new_n732), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1008), .A2(new_n693), .A3(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n678), .A2(new_n680), .A3(new_n790), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n826), .B1(new_n792), .B2(new_n761), .C1(new_n766), .C2(new_n754), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT117), .Z(new_n1037));
  AOI22_X1  g0837(.A1(G303), .A2(new_n819), .B1(new_n818), .B2(new_n952), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n757), .A2(G317), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n750), .A2(G322), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT48), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n748), .A2(G283), .B1(new_n770), .B2(G294), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT49), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1037), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n942), .A2(new_n747), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(G50), .B2(new_n757), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n744), .A2(new_n229), .B1(new_n761), .B2(new_n555), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(G159), .B2(new_n750), .ZN(new_n1054));
  INV_X1    g0854(.A(G150), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n762), .A2(new_n204), .B1(new_n754), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n259), .B2(new_n818), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1052), .A2(new_n1054), .A3(new_n330), .A4(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n783), .B1(new_n1050), .B2(new_n1058), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n243), .A2(new_n478), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1060), .A2(new_n796), .B1(new_n696), .B2(new_n791), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n258), .A2(G50), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT50), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n478), .B1(new_n229), .B2(new_n204), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n696), .B(new_n1064), .C1(new_n1063), .C2(new_n1062), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n1061), .A2(new_n1065), .B1(G107), .B2(new_n213), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n815), .B(new_n1059), .C1(new_n941), .C2(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1007), .A2(new_n974), .B1(new_n1035), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1034), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(KEYINPUT118), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT118), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1034), .A2(new_n1071), .A3(new_n1068), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1072), .ZN(G393));
  AND3_X1   g0873(.A1(new_n998), .A2(new_n691), .A3(new_n1002), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n691), .B1(new_n998), .B2(new_n1002), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1008), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1076), .A2(new_n1010), .A3(new_n693), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(G150), .A2(new_n750), .B1(new_n757), .B2(G159), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT51), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G50), .A2(new_n818), .B1(new_n771), .B2(G143), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n258), .B2(new_n744), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n748), .A2(G77), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n229), .B2(new_n762), .C1(new_n231), .C2(new_n761), .ZN(new_n1083));
  NOR4_X1   g0883(.A1(new_n1079), .A2(new_n826), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n762), .A2(new_n773), .B1(new_n761), .B2(new_n235), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n292), .B(new_n1085), .C1(G116), .C2(new_n748), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G294), .A2(new_n819), .B1(new_n771), .B2(G322), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1086), .B(new_n1087), .C1(new_n833), .C2(new_n742), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G311), .A2(new_n757), .B1(new_n750), .B2(G317), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT52), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n782), .B1(new_n1084), .B2(new_n1091), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n941), .B1(new_n555), .B2(new_n213), .C1(new_n943), .C2(new_n256), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT119), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n815), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1092), .B(new_n1095), .C1(new_n1094), .C2(new_n1093), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n985), .B2(new_n790), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1097), .B1(new_n1098), .B2(new_n974), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1077), .A2(new_n1099), .ZN(G390));
  AOI21_X1  g0900(.A(new_n815), .B1(new_n258), .B2(new_n816), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n1082), .B1(new_n758), .B2(new_n792), .C1(new_n773), .C2(new_n765), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n508), .A2(new_n818), .B1(new_n771), .B2(G294), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n231), .B2(new_n762), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n494), .B1(new_n229), .B2(new_n761), .C1(new_n555), .C2(new_n744), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n1102), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n771), .A2(G125), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1107), .B(new_n292), .C1(new_n220), .C2(new_n761), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(G159), .A2(new_n748), .B1(new_n750), .B2(G128), .ZN(new_n1109));
  INV_X1    g0909(.A(G132), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1109), .B1(new_n1110), .B2(new_n758), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT53), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n762), .B2(new_n1055), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n770), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1108), .B(new_n1111), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(KEYINPUT54), .B(G143), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n822), .A2(new_n742), .B1(new_n744), .B2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT121), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1106), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n913), .A2(new_n914), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1101), .B1(new_n783), .B2(new_n1119), .C1(new_n1120), .C2(new_n789), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n915), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n873), .B2(new_n884), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n807), .A2(new_n463), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n806), .B1(new_n706), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1123), .B1(new_n1125), .B2(new_n919), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1122), .B1(new_n918), .B2(new_n920), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n1127), .A2(KEYINPUT120), .B1(new_n913), .B2(new_n914), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT120), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1129), .B(new_n1122), .C1(new_n918), .C2(new_n920), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1126), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  NOR3_X1   g0931(.A1(new_n729), .A2(new_n809), .A3(new_n919), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1132), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1134), .B(new_n1126), .C1(new_n1128), .C2(new_n1130), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1121), .B1(new_n1136), .B2(new_n973), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n730), .A2(new_n924), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n925), .A2(new_n662), .A3(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n919), .B1(new_n729), .B2(new_n809), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n918), .B1(new_n1141), .B2(new_n1132), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1134), .A2(new_n1125), .A3(new_n1140), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1139), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1133), .A2(new_n1135), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1144), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n694), .B1(new_n1136), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1137), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(G378));
  INV_X1    g0949(.A(new_n1139), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1145), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n888), .A2(new_n885), .A3(new_n890), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(KEYINPUT110), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n858), .A2(new_n846), .A3(new_n885), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(G330), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n905), .B2(new_n859), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n275), .A2(new_n860), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n317), .B(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1160), .B(new_n1161), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n1155), .A2(new_n1157), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1162), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n1163), .A2(new_n1164), .A3(new_n923), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n923), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1162), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n902), .A2(new_n884), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT107), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n902), .A2(new_n884), .A3(KEYINPUT107), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n887), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(G330), .B1(new_n1172), .B2(KEYINPUT40), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1167), .B1(new_n892), .B2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1155), .A2(new_n1157), .A3(new_n1162), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1166), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1151), .B(KEYINPUT57), .C1(new_n1165), .C2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n923), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1174), .A2(new_n1166), .A3(new_n1175), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1178), .A2(new_n1179), .B1(new_n1145), .B2(new_n1150), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1177), .B(new_n693), .C1(KEYINPUT57), .C2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1167), .A2(new_n788), .ZN(new_n1183));
  INV_X1    g0983(.A(G41), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n826), .A2(new_n1184), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(G97), .A2(new_n818), .B1(new_n819), .B2(new_n441), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n773), .B2(new_n754), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n235), .A2(new_n758), .B1(new_n765), .B2(new_n792), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n827), .A2(G58), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(new_n204), .B2(new_n762), .C1(new_n229), .C2(new_n747), .ZN(new_n1190));
  NOR4_X1   g0990(.A1(new_n1185), .A2(new_n1187), .A3(new_n1188), .A4(new_n1190), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT58), .Z(new_n1192));
  OAI211_X1 g0992(.A(new_n1185), .B(new_n220), .C1(G33), .C2(G41), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1193), .B(KEYINPUT122), .Z(new_n1194));
  OAI22_X1  g0994(.A1(new_n762), .A2(new_n1116), .B1(new_n742), .B2(new_n1110), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G150), .A2(new_n748), .B1(new_n750), .B2(G125), .ZN(new_n1196));
  INV_X1    g0996(.A(G128), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1196), .B1(new_n1197), .B2(new_n758), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1195), .B(new_n1198), .C1(G137), .C2(new_n819), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n260), .B(new_n1184), .C1(new_n761), .C2(new_n755), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G124), .B2(new_n771), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT59), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1203), .B1(new_n1199), .B2(new_n1204), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1192), .B(new_n1194), .C1(new_n1201), .C2(new_n1205), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n1206), .A2(new_n782), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n815), .B(new_n1207), .C1(new_n220), .C2(new_n816), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1182), .A2(new_n974), .B1(new_n1183), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1181), .A2(new_n1209), .ZN(G375));
  NAND3_X1  g1010(.A1(new_n1139), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1146), .A2(new_n1013), .A3(new_n1211), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT123), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n815), .B1(new_n229), .B2(new_n816), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n773), .A2(new_n758), .B1(new_n765), .B2(new_n767), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n1215), .A2(new_n1051), .A3(new_n292), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n508), .A2(new_n819), .B1(new_n818), .B2(G116), .ZN(new_n1217));
  AND2_X1   g1017(.A1(new_n1217), .A2(KEYINPUT124), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(KEYINPUT124), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(G77), .A2(new_n827), .B1(new_n771), .B2(G303), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n555), .B2(new_n762), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n1218), .A2(new_n1219), .A3(new_n1221), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1189), .B1(new_n1197), .B2(new_n754), .C1(new_n765), .C2(new_n1110), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n819), .A2(G150), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n755), .B2(new_n762), .C1(new_n742), .C2(new_n1116), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n758), .A2(new_n822), .B1(new_n220), .B2(new_n747), .ZN(new_n1226));
  NOR3_X1   g1026(.A1(new_n1223), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1216), .A2(new_n1222), .B1(new_n1227), .B2(new_n330), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1214), .B1(new_n783), .B2(new_n1228), .C1(new_n920), .C2(new_n789), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1230), .B1(new_n1231), .B2(new_n974), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1213), .A2(new_n1232), .ZN(G381));
  NAND2_X1  g1033(.A1(new_n1182), .A2(new_n974), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1183), .A2(new_n1208), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1182), .A2(new_n1151), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT57), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1238), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n694), .B1(new_n1240), .B2(new_n1151), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1236), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n1148), .ZN(new_n1243));
  INV_X1    g1043(.A(G384), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1213), .A2(new_n1244), .A3(new_n1232), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1070), .A2(new_n804), .A3(new_n1072), .ZN(new_n1246));
  NOR4_X1   g1046(.A1(G387), .A2(new_n1245), .A3(G390), .A4(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1243), .B1(new_n1247), .B2(KEYINPUT125), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(KEYINPUT125), .B2(new_n1247), .ZN(G407));
  INV_X1    g1049(.A(new_n671), .ZN(new_n1250));
  OAI211_X1 g1050(.A(G407), .B(G213), .C1(new_n1250), .C2(new_n1243), .ZN(G409));
  OAI211_X1 g1051(.A(new_n972), .B(G390), .C1(new_n1014), .C2(new_n1030), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT127), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(G393), .B(new_n804), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(G390), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n1074), .A2(new_n1075), .A3(new_n1008), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1013), .B1(new_n1258), .B2(new_n1032), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1030), .B1(new_n1259), .B2(new_n973), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n972), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1257), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1252), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1256), .A2(new_n1263), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1262), .A2(new_n1255), .A3(KEYINPUT127), .A4(new_n1252), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT126), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1148), .B1(new_n1181), .B2(new_n1209), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1180), .A2(new_n1013), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1209), .A2(new_n1269), .A3(new_n1148), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1267), .B1(new_n1268), .B2(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(KEYINPUT126), .B(new_n1270), .C1(new_n1242), .C2(new_n1148), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT60), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(new_n1146), .B2(new_n1211), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1211), .A2(new_n1274), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n693), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1232), .B1(new_n1275), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1244), .ZN(new_n1279));
  OAI211_X1 g1079(.A(G384), .B(new_n1232), .C1(new_n1275), .C2(new_n1277), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n671), .A2(G213), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1272), .A2(new_n1273), .A3(new_n1282), .A4(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1284), .A2(KEYINPUT62), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1270), .B(new_n1283), .C1(new_n1242), .C2(new_n1148), .ZN(new_n1286));
  OAI21_X1  g1086(.A(KEYINPUT62), .B1(new_n1286), .B2(new_n1281), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n671), .A2(G213), .A3(G2897), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1281), .B(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT61), .B1(new_n1286), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1287), .A2(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1266), .B1(new_n1285), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1265), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n1254), .A2(new_n1255), .B1(new_n1262), .B2(new_n1252), .ZN(new_n1294));
  NOR3_X1   g1094(.A1(new_n1293), .A2(new_n1294), .A3(KEYINPUT61), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT63), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1284), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1272), .A2(new_n1273), .A3(new_n1283), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1289), .ZN(new_n1299));
  OR3_X1    g1099(.A1(new_n1286), .A2(new_n1296), .A3(new_n1281), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1295), .A2(new_n1297), .A3(new_n1299), .A4(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1292), .A2(new_n1301), .ZN(G405));
  INV_X1    g1102(.A(new_n1268), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1303), .A2(new_n1243), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1304), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1303), .A2(new_n1243), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1264), .A2(new_n1265), .A3(new_n1306), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1305), .A2(new_n1307), .A3(new_n1282), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1282), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1308), .A2(new_n1309), .ZN(G402));
endmodule


