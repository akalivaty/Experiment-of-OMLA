//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1247, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G226), .ZN(new_n210));
  INV_X1    g0010(.A(G116), .ZN(new_n211));
  INV_X1    g0011(.A(G270), .ZN(new_n212));
  OAI22_X1  g0012(.A1(new_n202), .A2(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G58), .B2(G232), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G107), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  OAI22_X1  g0018(.A1(new_n215), .A2(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n219), .B1(G87), .B2(G250), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT64), .B(G244), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G77), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n214), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G68), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT1), .Z(new_n228));
  NOR2_X1   g0028(.A1(new_n209), .A2(G13), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT0), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n232), .A2(new_n207), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(G50), .B1(G58), .B2(G68), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n228), .B(new_n231), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  INV_X1    g0038(.A(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT2), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n210), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G264), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n212), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(G107), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(new_n211), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  AND2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  OAI211_X1 g0055(.A(G232), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT73), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT3), .B(G33), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n259), .A2(KEYINPUT73), .A3(G232), .A4(G1698), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n259), .A2(G226), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G97), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n258), .A2(new_n260), .A3(new_n262), .A4(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  AND4_X1   g0065(.A1(KEYINPUT66), .A2(new_n265), .A3(G1), .A4(G13), .ZN(new_n266));
  AND2_X1   g0066(.A1(G1), .A2(G13), .ZN(new_n267));
  AOI21_X1  g0067(.A(KEYINPUT66), .B1(new_n267), .B2(new_n265), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n267), .A2(new_n265), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G238), .ZN(new_n275));
  INV_X1    g0075(.A(G274), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n271), .A2(new_n275), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT13), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT74), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT13), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n271), .A2(new_n282), .A3(new_n275), .A4(new_n278), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n280), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  OR3_X1    g0084(.A1(new_n279), .A2(new_n281), .A3(KEYINPUT13), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(new_n285), .A3(G169), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT14), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n280), .A2(G179), .A3(new_n283), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT14), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n284), .A2(new_n285), .A3(new_n289), .A4(G169), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n287), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n207), .A2(G33), .A3(G77), .ZN(new_n292));
  OAI21_X1  g0092(.A(KEYINPUT67), .B1(G20), .B2(G33), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NOR3_X1   g0094(.A1(KEYINPUT67), .A2(G20), .A3(G33), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI221_X1 g0096(.A(new_n292), .B1(new_n207), .B2(G68), .C1(new_n296), .C2(new_n202), .ZN(new_n297));
  NAND3_X1  g0097(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n232), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT75), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT75), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n297), .A2(new_n302), .A3(new_n299), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT11), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n206), .A2(G20), .ZN(new_n307));
  INV_X1    g0107(.A(G13), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n309), .A2(KEYINPUT12), .A3(new_n224), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n301), .A2(KEYINPUT11), .A3(new_n303), .ZN(new_n311));
  AOI21_X1  g0111(.A(KEYINPUT12), .B1(new_n309), .B2(new_n224), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n309), .A2(new_n299), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT68), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n307), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n206), .A2(KEYINPUT68), .A3(G20), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n313), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n312), .B1(new_n318), .B2(G68), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n306), .A2(new_n310), .A3(new_n311), .A4(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n291), .A2(new_n320), .ZN(new_n321));
  XOR2_X1   g0121(.A(KEYINPUT15), .B(G87), .Z(new_n322));
  NAND3_X1  g0122(.A1(new_n322), .A2(new_n207), .A3(G33), .ZN(new_n323));
  INV_X1    g0123(.A(G77), .ZN(new_n324));
  OR2_X1    g0124(.A1(KEYINPUT8), .A2(G58), .ZN(new_n325));
  NAND2_X1  g0125(.A1(KEYINPUT8), .A2(G58), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n323), .B1(new_n207), .B2(new_n324), .C1(new_n296), .C2(new_n327), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n328), .A2(new_n299), .B1(new_n324), .B2(new_n309), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(new_n324), .B2(new_n317), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G238), .A2(G1698), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n259), .B(new_n331), .C1(new_n239), .C2(G1698), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n270), .B(new_n332), .C1(G107), .C2(new_n259), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n274), .A2(new_n221), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(new_n278), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G169), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n330), .B(new_n337), .C1(G179), .C2(new_n335), .ZN(new_n338));
  AND2_X1   g0138(.A1(new_n321), .A2(new_n338), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n330), .A2(KEYINPUT69), .ZN(new_n340));
  INV_X1    g0140(.A(G190), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n330), .A2(KEYINPUT69), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n335), .A2(G200), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n340), .A2(new_n342), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(G150), .B1(new_n294), .B2(new_n295), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n203), .A2(G20), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n325), .A2(new_n207), .A3(G33), .A4(new_n326), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n299), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n309), .A2(new_n202), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n313), .A2(G50), .A3(new_n315), .A4(new_n316), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT70), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT9), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n350), .A2(new_n299), .B1(new_n202), .B2(new_n309), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT70), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n357), .A2(new_n358), .A3(new_n353), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n355), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT71), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT71), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n355), .A2(new_n362), .A3(new_n356), .A4(new_n359), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n254), .A2(new_n255), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(new_n261), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n259), .A2(G222), .A3(new_n261), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT65), .ZN(new_n367));
  AOI22_X1  g0167(.A1(G223), .A2(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n367), .B2(new_n366), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n259), .A2(new_n324), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n270), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n274), .A2(G226), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(new_n278), .A3(new_n372), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n361), .A2(new_n363), .B1(new_n373), .B2(G200), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n354), .A2(KEYINPUT70), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n358), .B1(new_n357), .B2(new_n353), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT9), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT72), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n355), .A2(new_n359), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT72), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n379), .A2(new_n380), .A3(KEYINPUT9), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n373), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G190), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n374), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT10), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n374), .A2(new_n382), .A3(KEYINPUT10), .A4(new_n384), .ZN(new_n388));
  INV_X1    g0188(.A(G179), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n383), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n390), .B(new_n354), .C1(G169), .C2(new_n383), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n387), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT18), .ZN(new_n394));
  INV_X1    g0194(.A(new_n327), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n395), .A2(new_n309), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n317), .B2(new_n395), .ZN(new_n397));
  INV_X1    g0197(.A(new_n299), .ZN(new_n398));
  XNOR2_X1  g0198(.A(G58), .B(G68), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G20), .ZN(new_n400));
  INV_X1    g0200(.A(G159), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n400), .B1(new_n296), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(G33), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT3), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT77), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT77), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT3), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n403), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT76), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n403), .ZN(new_n410));
  NAND2_X1  g0210(.A1(KEYINPUT76), .A2(G33), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n404), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n207), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n224), .B1(new_n413), .B2(KEYINPUT7), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n406), .A2(KEYINPUT3), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n404), .A2(KEYINPUT77), .ZN(new_n416));
  OAI21_X1  g0216(.A(G33), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AND2_X1   g0217(.A1(KEYINPUT76), .A2(G33), .ZN(new_n418));
  NOR2_X1   g0218(.A1(KEYINPUT76), .A2(G33), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT3), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(G20), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT7), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n402), .B1(new_n414), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n398), .B1(new_n424), .B2(KEYINPUT16), .ZN(new_n425));
  XOR2_X1   g0225(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n405), .A2(new_n407), .A3(new_n403), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n418), .A2(new_n419), .A3(KEYINPUT3), .ZN(new_n429));
  OAI211_X1 g0229(.A(KEYINPUT7), .B(new_n207), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n422), .B1(new_n259), .B2(G20), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n224), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n427), .B1(new_n432), .B2(new_n402), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n397), .B1(new_n425), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n210), .A2(G1698), .ZN(new_n435));
  OR2_X1    g0235(.A1(G223), .A2(G1698), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n417), .A2(new_n420), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G33), .A2(G87), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n269), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n274), .A2(G232), .ZN(new_n440));
  NOR4_X1   g0240(.A1(new_n439), .A2(new_n389), .A3(new_n440), .A4(new_n277), .ZN(new_n441));
  INV_X1    g0241(.A(new_n440), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n437), .A2(new_n438), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n278), .B(new_n442), .C1(new_n443), .C2(new_n269), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n441), .B1(G169), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n394), .B1(new_n434), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n402), .ZN(new_n447));
  OAI21_X1  g0247(.A(G68), .B1(new_n421), .B2(new_n422), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n413), .A2(KEYINPUT7), .ZN(new_n449));
  OAI211_X1 g0249(.A(KEYINPUT16), .B(new_n447), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(new_n433), .A3(new_n299), .ZN(new_n451));
  INV_X1    g0251(.A(new_n397), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NOR3_X1   g0253(.A1(new_n439), .A2(new_n277), .A3(new_n440), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G179), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(new_n454), .B2(new_n336), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n453), .A2(new_n456), .A3(KEYINPUT18), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n446), .A2(new_n457), .ZN(new_n458));
  OR2_X1    g0258(.A1(KEYINPUT79), .A2(G190), .ZN(new_n459));
  NAND2_X1  g0259(.A1(KEYINPUT79), .A2(G190), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NOR4_X1   g0262(.A1(new_n439), .A2(new_n277), .A3(new_n440), .A4(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n444), .A2(G200), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n451), .A2(new_n464), .A3(new_n465), .A4(new_n452), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT17), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT17), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n463), .B1(G200), .B2(new_n444), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n434), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n458), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n320), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n280), .A2(G190), .A3(new_n283), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n284), .A2(new_n285), .A3(G200), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n346), .A2(new_n393), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n309), .A2(new_n215), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n313), .B1(G1), .B2(new_n403), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n480), .B1(new_n481), .B2(new_n215), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT81), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n215), .A2(new_n217), .A3(KEYINPUT6), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT80), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT6), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G97), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n484), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n485), .B1(new_n484), .B2(new_n487), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n217), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n486), .A2(G97), .A3(G107), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n215), .A2(KEYINPUT6), .ZN(new_n492));
  OAI21_X1  g0292(.A(KEYINPUT80), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n484), .A2(new_n485), .A3(new_n487), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n493), .A2(new_n494), .A3(G107), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n207), .B1(new_n490), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n296), .A2(new_n324), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n483), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n488), .A2(new_n489), .A3(new_n217), .ZN(new_n499));
  AOI21_X1  g0299(.A(G107), .B1(new_n493), .B2(new_n494), .ZN(new_n500));
  OAI21_X1  g0300(.A(G20), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n497), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(KEYINPUT81), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n430), .A2(new_n431), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G107), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n498), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n482), .B1(new_n506), .B2(new_n299), .ZN(new_n507));
  INV_X1    g0307(.A(G45), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n508), .A2(G1), .ZN(new_n509));
  AND2_X1   g0309(.A1(KEYINPUT5), .A2(G41), .ZN(new_n510));
  NOR2_X1   g0310(.A1(KEYINPUT5), .A2(G41), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(G257), .A3(new_n272), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n509), .B(G274), .C1(new_n511), .C2(new_n510), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n259), .A2(KEYINPUT4), .A3(G244), .A4(new_n261), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G283), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n259), .A2(G250), .A3(G1698), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT4), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n417), .A2(G244), .A3(new_n261), .A4(new_n420), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n516), .B1(new_n523), .B2(new_n269), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n513), .A2(KEYINPUT82), .A3(new_n514), .ZN(new_n526));
  AOI21_X1  g0326(.A(KEYINPUT82), .B1(new_n513), .B2(new_n514), .ZN(new_n527));
  OAI22_X1  g0327(.A1(new_n523), .A2(new_n269), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n525), .A2(G190), .B1(new_n528), .B2(G200), .ZN(new_n529));
  AND2_X1   g0329(.A1(new_n507), .A2(new_n529), .ZN(new_n530));
  OAI22_X1  g0330(.A1(new_n525), .A2(G169), .B1(new_n528), .B2(G179), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n507), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n408), .A2(new_n412), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n534), .A2(new_n207), .A3(G68), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT19), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n536), .A2(new_n207), .A3(G33), .A4(G97), .ZN(new_n537));
  NOR3_X1   g0337(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(new_n207), .B2(new_n263), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n537), .B1(new_n539), .B2(new_n536), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n322), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n541), .A2(new_n299), .B1(new_n309), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n481), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n322), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n272), .B(G250), .C1(G1), .C2(new_n508), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n509), .A2(G274), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n410), .A2(G116), .A3(new_n411), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(G244), .A2(G1698), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n225), .B2(G1698), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n552), .B1(new_n534), .B2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n389), .B(new_n550), .C1(new_n555), .C2(new_n269), .ZN(new_n556));
  XNOR2_X1  g0356(.A(KEYINPUT77), .B(KEYINPUT3), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n420), .B(new_n554), .C1(new_n403), .C2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n269), .B1(new_n558), .B2(new_n551), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n336), .B1(new_n559), .B2(new_n549), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n546), .A2(new_n556), .A3(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n550), .B1(new_n555), .B2(new_n269), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(G200), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n559), .A2(new_n549), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G190), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n544), .A2(G87), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n563), .A2(new_n543), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n514), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n512), .A2(new_n272), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n570), .A2(new_n218), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n216), .A2(G1698), .ZN(new_n572));
  OR2_X1    g0372(.A1(G250), .A2(G1698), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n417), .A2(new_n420), .A3(new_n572), .A4(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n410), .A2(G294), .A3(new_n411), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI211_X1 g0376(.A(new_n569), .B(new_n571), .C1(new_n576), .C2(new_n270), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(G169), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n578), .B1(new_n389), .B2(new_n577), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT85), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT24), .ZN(new_n581));
  OAI21_X1  g0381(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n582));
  OR3_X1    g0382(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n582), .B(new_n583), .C1(new_n551), .C2(G20), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT84), .ZN(new_n585));
  XNOR2_X1  g0385(.A(new_n584), .B(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(KEYINPUT22), .A2(G20), .ZN(new_n587));
  OAI211_X1 g0387(.A(G87), .B(new_n587), .C1(new_n254), .C2(new_n255), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT83), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT83), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n259), .A2(new_n590), .A3(G87), .A4(new_n587), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n417), .A2(new_n207), .A3(G87), .A4(new_n420), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n592), .B1(KEYINPUT22), .B2(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n580), .B(new_n581), .C1(new_n586), .C2(new_n594), .ZN(new_n595));
  XNOR2_X1  g0395(.A(new_n584), .B(KEYINPUT84), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n593), .A2(KEYINPUT22), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n597), .A2(new_n589), .A3(new_n591), .ZN(new_n598));
  NAND2_X1  g0398(.A1(KEYINPUT85), .A2(KEYINPUT24), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n580), .A2(new_n581), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n596), .A2(new_n598), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n595), .A2(new_n601), .A3(new_n299), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n544), .A2(G107), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n309), .B(new_n217), .C1(KEYINPUT86), .C2(KEYINPUT25), .ZN(new_n604));
  NAND2_X1  g0404(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n605));
  XNOR2_X1  g0405(.A(new_n604), .B(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n602), .A2(new_n603), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n568), .B1(new_n579), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n577), .A2(new_n341), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n577), .B2(G200), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n610), .A2(new_n602), .A3(new_n603), .A4(new_n606), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n218), .A2(G1698), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n216), .A2(new_n261), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n417), .A2(new_n420), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n364), .A2(G303), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n269), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n570), .A2(new_n212), .ZN(new_n617));
  OR3_X1    g0417(.A1(new_n616), .A2(new_n569), .A3(new_n617), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n313), .B(G116), .C1(G1), .C2(new_n403), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n309), .A2(new_n211), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n518), .B(new_n207), .C1(G33), .C2(new_n215), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n211), .A2(G20), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n621), .A2(new_n299), .A3(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT20), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n619), .B(new_n620), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n618), .A2(KEYINPUT21), .A3(G169), .A4(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT21), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n627), .A2(G169), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n616), .A2(new_n569), .A3(new_n617), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NOR4_X1   g0432(.A1(new_n616), .A2(new_n389), .A3(new_n569), .A4(new_n617), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n627), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n628), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(G200), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  NOR4_X1   g0437(.A1(new_n616), .A2(new_n617), .A3(new_n462), .A4(new_n569), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n637), .A2(new_n627), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n533), .A2(new_n608), .A3(new_n611), .A4(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n479), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g0442(.A(new_n642), .B(KEYINPUT87), .ZN(G372));
  INV_X1    g0443(.A(new_n458), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n339), .A2(new_n477), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n644), .B1(new_n645), .B2(new_n471), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n387), .A2(new_n388), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n391), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n479), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT88), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n651), .B1(new_n556), .B2(new_n560), .ZN(new_n652));
  AOI21_X1  g0452(.A(KEYINPUT88), .B1(new_n562), .B2(new_n336), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT89), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n558), .A2(new_n551), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n270), .ZN(new_n657));
  AOI21_X1  g0457(.A(G169), .B1(new_n657), .B2(new_n550), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n559), .A2(new_n549), .A3(G179), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT88), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n560), .A2(new_n651), .ZN(new_n661));
  AOI21_X1  g0461(.A(KEYINPUT89), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n546), .B1(new_n655), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT90), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(new_n664), .A3(new_n567), .ZN(new_n665));
  INV_X1    g0465(.A(new_n546), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n660), .A2(KEYINPUT89), .A3(new_n661), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n654), .B1(new_n652), .B2(new_n653), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n567), .ZN(new_n670));
  OAI21_X1  g0470(.A(KEYINPUT90), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT26), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(new_n673), .A3(new_n532), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n507), .A2(new_n529), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n611), .B(new_n675), .C1(new_n531), .C2(new_n507), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n635), .B1(new_n607), .B2(new_n579), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n672), .A2(new_n678), .ZN(new_n679));
  NOR3_X1   g0479(.A1(new_n568), .A2(new_n507), .A3(new_n531), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n663), .B1(new_n680), .B2(new_n673), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n674), .A2(new_n679), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n650), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n649), .A2(new_n684), .ZN(G369));
  NOR2_X1   g0485(.A1(new_n308), .A2(G20), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n206), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(G213), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(G343), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n627), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g0493(.A(new_n693), .B(KEYINPUT91), .Z(new_n694));
  MUX2_X1   g0494(.A(new_n635), .B(new_n640), .S(new_n694), .Z(new_n695));
  AND2_X1   g0495(.A1(new_n695), .A2(G330), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n607), .A2(new_n579), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(new_n692), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n607), .A2(new_n692), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n611), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n698), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT92), .ZN(new_n703));
  INV_X1    g0503(.A(new_n692), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n635), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n698), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n703), .A2(new_n708), .ZN(G399));
  INV_X1    g0509(.A(new_n229), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G41), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n538), .A2(new_n211), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n712), .A2(G1), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(new_n235), .B2(new_n712), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT94), .ZN(new_n717));
  XOR2_X1   g0517(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n718));
  XNOR2_X1  g0518(.A(new_n717), .B(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT29), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n683), .A2(new_n720), .A3(new_n704), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n664), .B1(new_n663), .B2(new_n567), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n669), .A2(KEYINPUT90), .A3(new_n670), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n532), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n669), .B1(new_n725), .B2(KEYINPUT26), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n680), .A2(new_n673), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT95), .B1(new_n672), .B2(new_n678), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n672), .A2(new_n678), .A3(KEYINPUT95), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n726), .B(new_n727), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n704), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n722), .B1(new_n731), .B2(KEYINPUT29), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n522), .A2(new_n521), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n733), .A2(new_n518), .A3(new_n519), .A4(new_n517), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n270), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n526), .A2(new_n527), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n577), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n737), .A2(new_n389), .A3(new_n562), .A4(new_n618), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n571), .B1(new_n576), .B2(new_n270), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n524), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n741), .A2(KEYINPUT30), .A3(new_n564), .A4(new_n633), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT30), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n735), .A2(new_n739), .A3(new_n516), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n633), .A2(new_n564), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n738), .A2(new_n742), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n692), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n507), .A2(new_n531), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n749), .A2(new_n640), .A3(new_n675), .A4(new_n611), .ZN(new_n750));
  INV_X1    g0550(.A(new_n568), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n697), .A2(new_n751), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n750), .A2(new_n752), .A3(new_n692), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT31), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n748), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n747), .A2(KEYINPUT31), .A3(new_n692), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G330), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n732), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n719), .B1(new_n759), .B2(G1), .ZN(G364));
  AOI21_X1  g0560(.A(new_n206), .B1(new_n686), .B2(G45), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n711), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n696), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n764), .B1(G330), .B2(new_n695), .ZN(new_n765));
  INV_X1    g0565(.A(new_n763), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n232), .B1(G20), .B2(new_n336), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n207), .A2(new_n389), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G200), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(new_n461), .ZN(new_n771));
  INV_X1    g0571(.A(G322), .ZN(new_n772));
  INV_X1    g0572(.A(G283), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n207), .A2(G179), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(new_n341), .A3(G200), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n771), .A2(new_n772), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G190), .A2(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G329), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n341), .A2(G179), .A3(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n207), .ZN(new_n781));
  INV_X1    g0581(.A(G294), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n364), .B1(new_n778), .B2(new_n779), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n768), .A2(new_n777), .ZN(new_n784));
  INV_X1    g0584(.A(G311), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n774), .A2(G190), .A3(G200), .ZN(new_n787));
  INV_X1    g0587(.A(G303), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR4_X1   g0589(.A1(new_n776), .A2(new_n783), .A3(new_n786), .A4(new_n789), .ZN(new_n790));
  OR3_X1    g0590(.A1(new_n769), .A2(new_n636), .A3(KEYINPUT96), .ZN(new_n791));
  OAI21_X1  g0591(.A(KEYINPUT96), .B1(new_n769), .B2(new_n636), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n462), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G326), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n791), .A2(new_n341), .A3(new_n792), .ZN(new_n797));
  XOR2_X1   g0597(.A(KEYINPUT33), .B(G317), .Z(new_n798));
  OAI221_X1 g0598(.A(new_n790), .B1(new_n795), .B2(new_n796), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n784), .A2(new_n324), .ZN(new_n800));
  INV_X1    g0600(.A(new_n797), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n794), .A2(G50), .B1(new_n801), .B2(G68), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT32), .ZN(new_n803));
  INV_X1    g0603(.A(new_n778), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n803), .B1(new_n804), .B2(G159), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n778), .A2(KEYINPUT32), .A3(new_n401), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n775), .A2(new_n217), .ZN(new_n807));
  INV_X1    g0607(.A(G87), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n787), .A2(new_n808), .ZN(new_n809));
  NOR4_X1   g0609(.A1(new_n805), .A2(new_n806), .A3(new_n807), .A4(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n259), .B1(new_n781), .B2(new_n215), .ZN(new_n811));
  INV_X1    g0611(.A(new_n771), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n811), .B1(new_n812), .B2(G58), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n802), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n799), .B1(new_n800), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n249), .A2(G45), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n710), .A2(new_n534), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n816), .B(new_n817), .C1(G45), .C2(new_n235), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n229), .A2(G355), .A3(new_n259), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n818), .B(new_n819), .C1(G116), .C2(new_n229), .ZN(new_n820));
  NOR2_X1   g0620(.A1(G13), .A2(G33), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(G20), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(new_n767), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n767), .A2(new_n815), .B1(new_n820), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n823), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n825), .B1(new_n695), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n765), .B1(new_n766), .B2(new_n827), .ZN(G396));
  NAND2_X1  g0628(.A1(new_n330), .A2(new_n692), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n345), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n338), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n338), .A2(new_n692), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n683), .B2(new_n704), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n681), .B1(new_n672), .B2(new_n678), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n692), .B(new_n833), .C1(new_n836), .C2(new_n674), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(new_n758), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n766), .ZN(new_n840));
  INV_X1    g0640(.A(new_n784), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n794), .A2(G137), .B1(G159), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(G143), .ZN(new_n843));
  INV_X1    g0643(.A(G150), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n842), .B1(new_n843), .B2(new_n771), .C1(new_n844), .C2(new_n797), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT34), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n775), .A2(new_n224), .ZN(new_n847));
  INV_X1    g0647(.A(G132), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n534), .B1(new_n848), .B2(new_n778), .ZN(new_n849));
  INV_X1    g0649(.A(new_n781), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n847), .B(new_n849), .C1(G58), .C2(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n846), .B(new_n851), .C1(new_n202), .C2(new_n787), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n795), .A2(new_n788), .B1(new_n797), .B2(new_n773), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n364), .B1(new_n778), .B2(new_n785), .C1(new_n781), .C2(new_n215), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n775), .A2(new_n808), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n856), .B1(new_n217), .B2(new_n787), .C1(new_n771), .C2(new_n782), .ZN(new_n857));
  NOR3_X1   g0657(.A1(new_n853), .A2(new_n854), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n211), .B2(new_n784), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n852), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n767), .A2(new_n821), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n860), .A2(new_n767), .B1(new_n324), .B2(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n862), .B(new_n763), .C1(new_n822), .C2(new_n834), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n863), .B(KEYINPUT97), .Z(new_n864));
  NAND2_X1  g0664(.A1(new_n840), .A2(new_n864), .ZN(G384));
  INV_X1    g0665(.A(KEYINPUT40), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT103), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n756), .B(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n755), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n320), .A2(new_n692), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n321), .A2(new_n476), .A3(new_n871), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n320), .B(new_n692), .C1(new_n477), .C2(new_n291), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n833), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT38), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n427), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n397), .B1(new_n425), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT98), .B1(new_n878), .B2(new_n690), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n450), .A2(new_n299), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n424), .A2(new_n426), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n452), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT98), .ZN(new_n883));
  INV_X1    g0683(.A(new_n690), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n882), .A2(new_n456), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n879), .A2(new_n885), .A3(new_n466), .A4(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT99), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT37), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n466), .A2(new_n889), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n445), .A2(new_n690), .B1(new_n451), .B2(new_n452), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n453), .B1(new_n456), .B2(new_n884), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n893), .A2(KEYINPUT99), .A3(new_n889), .A4(new_n466), .ZN(new_n894));
  AOI22_X1  g0694(.A1(KEYINPUT37), .A2(new_n887), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n458), .A2(new_n471), .B1(new_n885), .B2(new_n879), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n875), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n892), .A2(new_n894), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n879), .A2(new_n885), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n472), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n900), .A2(KEYINPUT38), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n897), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n870), .A2(new_n874), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT31), .B1(new_n641), .B2(new_n692), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n868), .B1(new_n906), .B2(new_n748), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n872), .A2(new_n873), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n834), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT100), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n466), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n434), .A2(KEYINPUT100), .A3(new_n469), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n912), .A2(new_n913), .A3(new_n893), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n892), .A2(new_n894), .B1(new_n914), .B2(KEYINPUT37), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n453), .A2(new_n884), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n458), .B2(new_n471), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n875), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n866), .B1(new_n903), .B2(new_n918), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n866), .A2(new_n905), .B1(new_n910), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT104), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n650), .A2(new_n870), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n921), .B(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(G330), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT102), .B1(new_n732), .B2(new_n479), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT102), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n720), .B1(new_n730), .B2(new_n704), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n926), .B(new_n650), .C1(new_n927), .C2(new_n722), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n648), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n321), .A2(new_n692), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT101), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n895), .A2(new_n875), .A3(new_n896), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT38), .B1(new_n900), .B2(new_n902), .ZN(new_n933));
  OAI21_X1  g0733(.A(KEYINPUT39), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT39), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n903), .A2(new_n918), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n931), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n931), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n930), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n908), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n683), .A2(new_n704), .A3(new_n834), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n941), .B1(new_n942), .B2(new_n832), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n943), .A2(new_n904), .B1(new_n644), .B2(new_n690), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n929), .B(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n924), .B(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n206), .B2(new_n686), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n490), .A2(new_n495), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n211), .B1(new_n949), .B2(KEYINPUT35), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n950), .B(new_n233), .C1(KEYINPUT35), .C2(new_n949), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT36), .ZN(new_n952));
  INV_X1    g0752(.A(G58), .ZN(new_n953));
  OAI21_X1  g0753(.A(G77), .B1(new_n953), .B2(new_n224), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n954), .A2(new_n235), .B1(G50), .B2(new_n224), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n955), .A2(G1), .A3(new_n308), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n948), .A2(new_n952), .A3(new_n956), .ZN(G367));
  NOR2_X1   g0757(.A1(new_n507), .A2(new_n704), .ZN(new_n958));
  NOR3_X1   g0758(.A1(new_n530), .A2(new_n532), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(new_n532), .B2(new_n692), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n706), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT42), .ZN(new_n962));
  NOR4_X1   g0762(.A1(new_n697), .A2(new_n530), .A3(new_n532), .A4(new_n958), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n704), .B1(new_n963), .B2(new_n532), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n704), .B1(new_n543), .B2(new_n566), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n672), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n663), .B2(new_n967), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n965), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n703), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n972), .A2(new_n960), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n971), .B(new_n973), .Z(new_n974));
  NOR2_X1   g0774(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n974), .B(new_n975), .Z(new_n976));
  XNOR2_X1  g0776(.A(new_n711), .B(KEYINPUT41), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n708), .A2(new_n960), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT45), .Z(new_n980));
  NAND2_X1  g0780(.A1(new_n708), .A2(new_n960), .ZN(new_n981));
  XNOR2_X1  g0781(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n981), .B(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT106), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n972), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n701), .B(new_n705), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(new_n696), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n759), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n703), .B1(new_n980), .B2(new_n983), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n986), .B(new_n989), .C1(new_n990), .C2(new_n985), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n978), .B1(new_n991), .B2(new_n759), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n976), .B1(new_n992), .B2(new_n762), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n795), .A2(new_n843), .B1(new_n797), .B2(new_n401), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n784), .A2(new_n202), .ZN(new_n995));
  INV_X1    g0795(.A(new_n775), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(G77), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n953), .B2(new_n787), .C1(new_n771), .C2(new_n844), .ZN(new_n998));
  INV_X1    g0798(.A(G137), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n259), .B1(new_n778), .B2(new_n999), .C1(new_n781), .C2(new_n224), .ZN(new_n1000));
  NOR4_X1   g0800(.A1(new_n994), .A2(new_n995), .A3(new_n998), .A4(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n775), .A2(new_n215), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n812), .B2(G303), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n217), .B2(new_n781), .C1(new_n782), .C2(new_n797), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n787), .A2(new_n211), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n534), .B1(KEYINPUT46), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(G317), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1006), .B1(KEYINPUT46), .B2(new_n1005), .C1(new_n1007), .C2(new_n778), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1004), .B(new_n1008), .C1(G311), .C2(new_n794), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n841), .A2(G283), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1001), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n766), .B1(new_n1013), .B2(new_n767), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n817), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n824), .B1(new_n229), .B2(new_n542), .C1(new_n245), .C2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1014), .B(new_n1016), .C1(new_n826), .C2(new_n969), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT108), .Z(new_n1018));
  NAND2_X1  g0818(.A1(new_n993), .A2(new_n1018), .ZN(G387));
  AOI22_X1  g0819(.A1(new_n794), .A2(G322), .B1(G303), .B2(new_n841), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n785), .B2(new_n797), .C1(new_n1007), .C2(new_n771), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT48), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n773), .B2(new_n781), .C1(new_n782), .C2(new_n787), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT109), .Z(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT49), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n534), .B1(G116), .B2(new_n996), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(new_n796), .C2(new_n778), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n534), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1002), .B(new_n1028), .C1(G150), .C2(new_n804), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n787), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(G77), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n542), .A2(new_n781), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n812), .A2(G50), .B1(G68), .B2(new_n841), .ZN(new_n1034));
  AND4_X1   g0834(.A1(new_n1029), .A2(new_n1031), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n401), .B2(new_n795), .C1(new_n327), .C2(new_n797), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1027), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n767), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n701), .A2(new_n826), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n327), .A2(G50), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT50), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n714), .B1(new_n224), .B2(new_n324), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1042));
  AOI211_X1 g0842(.A(G45), .B(new_n1042), .C1(new_n1041), .C2(new_n1040), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n817), .B1(new_n242), .B2(new_n508), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n229), .A2(new_n259), .A3(new_n713), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n229), .A2(G107), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n824), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1038), .A2(new_n763), .A3(new_n1039), .A4(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n988), .A2(new_n762), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n711), .B1(new_n759), .B2(new_n988), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1049), .B(new_n1050), .C1(new_n989), .C2(new_n1051), .ZN(G393));
  AND2_X1   g0852(.A1(new_n990), .A2(KEYINPUT110), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n990), .A2(KEYINPUT110), .ZN(new_n1054));
  NOR3_X1   g0854(.A1(new_n980), .A2(new_n703), .A3(new_n983), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n711), .B(new_n991), .C1(new_n1056), .C2(new_n989), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n960), .A2(new_n823), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n824), .B1(new_n215), .B2(new_n229), .C1(new_n252), .C2(new_n1015), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n794), .A2(G150), .B1(new_n812), .B2(G159), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT51), .Z(new_n1061));
  OAI21_X1  g0861(.A(new_n534), .B1(new_n843), .B2(new_n778), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n856), .B1(new_n224), .B2(new_n787), .C1(new_n324), .C2(new_n781), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(G50), .C2(new_n801), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1061), .B(new_n1064), .C1(new_n327), .C2(new_n784), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n781), .A2(new_n211), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n794), .A2(G317), .B1(new_n812), .B2(G311), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT52), .Z(new_n1068));
  OAI21_X1  g0868(.A(new_n364), .B1(new_n778), .B2(new_n772), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n807), .B(new_n1069), .C1(G283), .C2(new_n1030), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT111), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n801), .A2(G303), .B1(G294), .B2(new_n841), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1068), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1065), .B1(new_n1066), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n766), .B1(new_n1074), .B2(new_n767), .ZN(new_n1075));
  AND3_X1   g0875(.A1(new_n1058), .A2(new_n1059), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n1056), .B2(new_n762), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1057), .A2(new_n1077), .ZN(G390));
  NAND3_X1  g0878(.A1(new_n730), .A2(new_n704), .A3(new_n831), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n941), .B1(new_n1079), .B2(new_n832), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n903), .A2(new_n918), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n930), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AND3_X1   g0883(.A1(new_n903), .A2(new_n918), .A3(new_n935), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n935), .B1(new_n897), .B2(new_n903), .ZN(new_n1085));
  OAI21_X1  g0885(.A(KEYINPUT101), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n938), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n942), .A2(new_n832), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n930), .B1(new_n1088), .B2(new_n908), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n1080), .A2(new_n1083), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(G330), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n833), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n870), .A2(new_n908), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n757), .A2(new_n1092), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n908), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n1097), .B1(new_n1087), .B2(new_n1089), .C1(new_n1080), .C2(new_n1083), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n762), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n794), .A2(G283), .B1(new_n801), .B2(G107), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n812), .A2(G116), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n259), .B(new_n809), .C1(G294), .C2(new_n804), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n784), .A2(new_n215), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n1104), .B(new_n847), .C1(G77), .C2(new_n850), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .A4(new_n1105), .ZN(new_n1106));
  XOR2_X1   g0906(.A(KEYINPUT54), .B(G143), .Z(new_n1107));
  AOI22_X1  g0907(.A1(new_n801), .A2(G137), .B1(new_n841), .B2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT112), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1030), .A2(G150), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT53), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n771), .A2(new_n848), .B1(new_n202), .B2(new_n775), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n259), .B1(new_n781), .B2(new_n401), .ZN(new_n1113));
  NOR3_X1   g0913(.A1(new_n1111), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(G128), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1109), .B(new_n1114), .C1(new_n1115), .C2(new_n795), .ZN(new_n1116));
  INV_X1    g0916(.A(G125), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n778), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1106), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1119), .A2(new_n767), .B1(new_n327), .B2(new_n861), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n763), .B(new_n1120), .C1(new_n1087), .C2(new_n822), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n922), .A2(new_n1091), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1093), .B1(new_n1095), .B2(new_n908), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n1088), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n870), .A2(new_n1092), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n941), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1096), .A2(new_n832), .A3(new_n1128), .A4(new_n1079), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n929), .A2(new_n1124), .A3(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n711), .B1(new_n1122), .B2(new_n1131), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n648), .B(new_n1123), .C1(new_n925), .C2(new_n928), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1099), .B1(new_n1133), .B2(new_n1130), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1100), .B(new_n1121), .C1(new_n1132), .C2(new_n1134), .ZN(G378));
  OAI22_X1  g0935(.A1(new_n795), .A2(new_n1117), .B1(new_n797), .B2(new_n848), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1030), .A2(new_n1107), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT115), .Z(new_n1138));
  OAI221_X1 g0938(.A(new_n1138), .B1(new_n1115), .B2(new_n771), .C1(new_n844), .C2(new_n781), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1136), .B(new_n1139), .C1(G137), .C2(new_n841), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT59), .ZN(new_n1141));
  AOI21_X1  g0941(.A(G33), .B1(new_n804), .B2(G124), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(G41), .B1(new_n996), .B2(G159), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT114), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n794), .A2(G116), .B1(G68), .B2(new_n850), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT113), .ZN(new_n1147));
  INV_X1    g0947(.A(G41), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1028), .B(new_n1148), .C1(new_n773), .C2(new_n778), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1031), .B1(new_n542), .B2(new_n784), .C1(new_n771), .C2(new_n217), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1149), .B(new_n1150), .C1(G97), .C2(new_n801), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1147), .B(new_n1151), .C1(new_n953), .C2(new_n775), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT58), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(G41), .B1(new_n534), .B2(G33), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1154), .B1(G50), .B2(new_n1155), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n1143), .A2(new_n1144), .B1(new_n1145), .B2(new_n1156), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(new_n1145), .B2(new_n1156), .C1(new_n1153), .C2(new_n1152), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1158), .A2(new_n767), .B1(new_n202), .B2(new_n861), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT56), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n379), .A2(new_n690), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n392), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT55), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1161), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n387), .A2(new_n388), .A3(new_n391), .A4(new_n1164), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1162), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1163), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1160), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(KEYINPUT55), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1162), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1170), .A2(KEYINPUT56), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1168), .A2(new_n1172), .A3(new_n821), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1159), .A2(new_n763), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT117), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n1168), .A2(new_n1172), .A3(KEYINPUT116), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1082), .B1(new_n1086), .B2(new_n938), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n832), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n904), .B(new_n908), .C1(new_n837), .C2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n644), .A2(new_n690), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1177), .B1(new_n1178), .B2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1168), .A2(new_n1172), .A3(KEYINPUT116), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n940), .A2(new_n944), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT116), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1168), .A2(new_n1172), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n920), .A2(G330), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n1183), .A2(new_n1185), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1188), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1176), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1188), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n1178), .A2(new_n1177), .A3(new_n1182), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1184), .B1(new_n940), .B2(new_n944), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1192), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1183), .A2(new_n1185), .A3(new_n1188), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1195), .A2(KEYINPUT117), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1191), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1175), .B1(new_n1198), .B2(new_n762), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1133), .B1(new_n1122), .B2(new_n1131), .ZN(new_n1200));
  AOI21_X1  g1000(.A(KEYINPUT57), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n749), .B1(new_n665), .B2(new_n671), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n663), .B1(new_n1202), .B2(new_n673), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT95), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n679), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n672), .A2(new_n678), .A3(KEYINPUT95), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1203), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n692), .B1(new_n1207), .B2(new_n727), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n721), .B1(new_n1208), .B2(new_n720), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n926), .B1(new_n1209), .B2(new_n650), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n928), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n649), .B(new_n1124), .C1(new_n1210), .C2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n1099), .B2(new_n1130), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1195), .A2(KEYINPUT57), .A3(new_n1196), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n711), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1199), .B1(new_n1201), .B2(new_n1215), .ZN(G375));
  INV_X1    g1016(.A(new_n1130), .ZN(new_n1217));
  OAI21_X1  g1017(.A(KEYINPUT119), .B1(new_n1217), .B2(new_n761), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n771), .A2(new_n999), .B1(new_n202), .B2(new_n781), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1028), .B(new_n1219), .C1(G58), .C2(new_n996), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n787), .A2(new_n401), .B1(new_n778), .B2(new_n1115), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT122), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n841), .A2(G150), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n801), .A2(new_n1107), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1220), .A2(new_n1222), .A3(new_n1223), .A4(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n794), .A2(G132), .ZN(new_n1226));
  XOR2_X1   g1026(.A(new_n1226), .B(KEYINPUT121), .Z(new_n1227));
  OAI21_X1  g1027(.A(new_n364), .B1(new_n778), .B2(new_n788), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n997), .B1(new_n215), .B2(new_n787), .C1(new_n217), .C2(new_n784), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1228), .B(new_n1229), .C1(G116), .C2(new_n801), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n782), .B2(new_n795), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1033), .B1(new_n773), .B2(new_n771), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT120), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n1225), .A2(new_n1227), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1234), .A2(new_n767), .B1(new_n224), .B2(new_n861), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n763), .B(new_n1235), .C1(new_n908), .C2(new_n822), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT119), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1130), .A2(new_n1237), .A3(new_n762), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1218), .A2(new_n1236), .A3(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1130), .B1(new_n929), .B2(new_n1124), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n977), .B(KEYINPUT118), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1131), .A2(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1239), .B1(new_n1240), .B2(new_n1242), .ZN(G381));
  NOR4_X1   g1043(.A1(G387), .A2(G390), .A3(G396), .A4(G393), .ZN(new_n1244));
  INV_X1    g1044(.A(G378), .ZN(new_n1245));
  INV_X1    g1045(.A(G375), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  OR3_X1    g1047(.A1(new_n1247), .A2(G384), .A3(G381), .ZN(G407));
  NAND3_X1  g1048(.A1(new_n1246), .A2(new_n691), .A3(new_n1245), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(G407), .A2(G213), .A3(new_n1249), .ZN(G409));
  INV_X1    g1050(.A(KEYINPUT61), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n691), .A2(G213), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1198), .A2(new_n1200), .A3(new_n1241), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1195), .A2(new_n762), .A3(new_n1196), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1253), .A2(new_n1174), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1245), .ZN(new_n1256));
  OAI211_X1 g1056(.A(G378), .B(new_n1199), .C1(new_n1201), .C2(new_n1215), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1252), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1252), .A2(G2897), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT60), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1261), .B1(new_n1133), .B2(new_n1130), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1212), .A2(KEYINPUT60), .A3(new_n1217), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1262), .A2(new_n711), .A3(new_n1131), .A4(new_n1263), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1264), .A2(G384), .A3(new_n1239), .ZN(new_n1265));
  AOI21_X1  g1065(.A(G384), .B1(new_n1264), .B2(new_n1239), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1260), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n711), .B(new_n1131), .C1(new_n1240), .C2(KEYINPUT60), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1263), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1239), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(G384), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1264), .A2(G384), .A3(new_n1239), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1272), .A2(new_n1273), .A3(new_n1259), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1267), .A2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1251), .B1(new_n1258), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT125), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(KEYINPUT125), .B(new_n1251), .C1(new_n1258), .C2(new_n1275), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1258), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1258), .A2(new_n1280), .ZN(new_n1283));
  XOR2_X1   g1083(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1278), .A2(new_n1279), .A3(new_n1282), .A4(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(G390), .B1(new_n993), .B2(new_n1018), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(G393), .B(G396), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n993), .A2(new_n1018), .A3(G390), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1288), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1290), .B1(new_n1288), .B2(new_n1291), .ZN(new_n1293));
  OR2_X1    g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1286), .A2(new_n1294), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(KEYINPUT123), .B(KEYINPUT63), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1276), .B1(new_n1283), .B2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1258), .A2(KEYINPUT63), .A3(new_n1280), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT124), .ZN(new_n1299));
  OR2_X1    g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1297), .A2(new_n1300), .A3(new_n1301), .A4(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1295), .A2(new_n1303), .ZN(G405));
  NAND2_X1  g1104(.A1(G375), .A2(new_n1245), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1280), .A2(new_n1245), .A3(G375), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1309), .A2(KEYINPUT127), .A3(new_n1257), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1257), .A2(KEYINPUT127), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1307), .A2(new_n1308), .A3(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(new_n1313), .B(new_n1294), .ZN(G402));
endmodule


