//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0 1 0 0 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n991, new_n992, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1009,
    new_n1010, new_n1011, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1026, new_n1027, new_n1028, new_n1029, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1036, new_n1037, new_n1038,
    new_n1039;
  XNOR2_X1  g000(.A(KEYINPUT87), .B(G36gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G29gat), .ZN(new_n203));
  INV_X1    g002(.A(G50gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G43gat), .ZN(new_n205));
  INV_X1    g004(.A(G43gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G50gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  AND3_X1   g008(.A1(new_n203), .A2(KEYINPUT15), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT15), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  OR3_X1    g011(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n212), .A2(new_n203), .A3(new_n215), .A4(KEYINPUT88), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n213), .A2(KEYINPUT86), .A3(new_n214), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n214), .A2(KEYINPUT86), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n210), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n212), .A2(new_n203), .A3(new_n215), .ZN(new_n220));
  OAI22_X1  g019(.A1(new_n220), .A2(KEYINPUT88), .B1(new_n211), .B2(new_n208), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT89), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n219), .A2(new_n221), .A3(KEYINPUT89), .ZN(new_n225));
  XNOR2_X1  g024(.A(G15gat), .B(G22gat), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n226), .A2(G1gat), .ZN(new_n227));
  INV_X1    g026(.A(G8gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT16), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n226), .B1(new_n229), .B2(G1gat), .ZN(new_n230));
  AND3_X1   g029(.A1(new_n227), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n228), .B1(new_n227), .B2(new_n230), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n224), .A2(new_n225), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT90), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n224), .A2(new_n225), .ZN(new_n236));
  INV_X1    g035(.A(new_n233), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  AOI211_X1 g037(.A(KEYINPUT90), .B(new_n233), .C1(new_n224), .C2(new_n225), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n234), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G229gat), .A2(G233gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(KEYINPUT13), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n225), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT89), .B1(new_n219), .B2(new_n221), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n237), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT90), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n236), .A2(new_n235), .A3(new_n237), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT17), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n251), .B1(new_n245), .B2(new_n246), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n222), .A2(KEYINPUT17), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(new_n233), .A3(new_n253), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n250), .A2(KEYINPUT18), .A3(new_n241), .A4(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G113gat), .B(G141gat), .ZN(new_n256));
  INV_X1    g055(.A(G197gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(KEYINPUT11), .B(G169gat), .Z(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n260), .B(KEYINPUT12), .Z(new_n261));
  AND3_X1   g060(.A1(new_n244), .A2(new_n255), .A3(new_n261), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n254), .B(new_n241), .C1(new_n238), .C2(new_n239), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT91), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT18), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT91), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n250), .A2(new_n266), .A3(new_n241), .A4(new_n254), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n264), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n262), .A2(KEYINPUT93), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT93), .B1(new_n262), .B2(new_n268), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n244), .A2(new_n255), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT92), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n272), .B1(new_n268), .B2(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n264), .A2(KEYINPUT92), .A3(new_n265), .A4(new_n267), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n261), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n271), .A2(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(G190gat), .B(G218gat), .Z(new_n278));
  INV_X1    g077(.A(G85gat), .ZN(new_n279));
  INV_X1    g078(.A(G92gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OR2_X1    g080(.A1(KEYINPUT99), .A2(KEYINPUT7), .ZN(new_n282));
  NAND2_X1  g081(.A1(KEYINPUT99), .A2(KEYINPUT7), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT100), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT100), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n281), .A2(new_n282), .A3(new_n286), .A4(new_n283), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT7), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n285), .B(new_n287), .C1(new_n288), .C2(new_n281), .ZN(new_n289));
  XOR2_X1   g088(.A(G99gat), .B(G106gat), .Z(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT101), .B(G85gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(G99gat), .A2(G106gat), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n292), .A2(new_n280), .B1(KEYINPUT8), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n289), .A2(new_n291), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n291), .B1(new_n289), .B2(new_n294), .ZN(new_n297));
  OR3_X1    g096(.A1(new_n296), .A2(KEYINPUT102), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT102), .B1(new_n296), .B2(new_n297), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n252), .A2(new_n253), .A3(new_n298), .A4(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n296), .A2(new_n297), .ZN(new_n301));
  NAND2_X1  g100(.A1(G232gat), .A2(G233gat), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n236), .A2(new_n301), .B1(KEYINPUT41), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n278), .B1(new_n300), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n300), .A2(new_n278), .A3(new_n304), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n303), .A2(KEYINPUT41), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n309), .B(G134gat), .ZN(new_n310));
  INV_X1    g109(.A(G162gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n312), .B1(new_n305), .B2(KEYINPUT103), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n306), .A2(new_n307), .A3(KEYINPUT103), .A4(new_n312), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT96), .B(KEYINPUT20), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT95), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  XOR2_X1   g120(.A(G57gat), .B(G64gat), .Z(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n320), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT94), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G71gat), .B(G78gat), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT21), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(new_n233), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT98), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT98), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n332), .A2(new_n335), .A3(new_n233), .ZN(new_n336));
  INV_X1    g135(.A(G231gat), .ZN(new_n337));
  INV_X1    g136(.A(G233gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n334), .A2(new_n336), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n339), .B1(new_n334), .B2(new_n336), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n318), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n342), .ZN(new_n344));
  INV_X1    g143(.A(new_n318), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n344), .A2(new_n340), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G183gat), .B(G211gat), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n331), .A2(KEYINPUT21), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n350), .A2(new_n352), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n349), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n355), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(new_n348), .A3(new_n353), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(G127gat), .B(G155gat), .Z(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n360), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n356), .A2(new_n358), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n361), .A2(new_n343), .A3(new_n346), .A4(new_n363), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT104), .B1(new_n317), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n367), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT104), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(new_n370), .A3(new_n316), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n329), .B(new_n330), .C1(new_n296), .C2(new_n297), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n373));
  INV_X1    g172(.A(new_n297), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n374), .A2(new_n295), .A3(new_n331), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n372), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n301), .A2(KEYINPUT10), .A3(new_n331), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G230gat), .A2(G233gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n372), .A2(new_n375), .ZN(new_n381));
  INV_X1    g180(.A(new_n379), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G120gat), .B(G148gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(G176gat), .B(G204gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n380), .A2(new_n383), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT105), .B1(new_n378), .B2(new_n379), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT105), .ZN(new_n392));
  AOI211_X1 g191(.A(new_n392), .B(new_n382), .C1(new_n376), .C2(new_n377), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n391), .A2(new_n394), .A3(new_n383), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n389), .B1(new_n395), .B2(new_n386), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n368), .A2(new_n371), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(G127gat), .ZN(new_n398));
  INV_X1    g197(.A(G134gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(G127gat), .A2(G134gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G120gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(G113gat), .ZN(new_n404));
  INV_X1    g203(.A(G113gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(G120gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT1), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n402), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G113gat), .B(G120gat), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n400), .B1(new_n411), .B2(KEYINPUT1), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n398), .A2(KEYINPUT69), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n398), .A2(KEYINPUT69), .ZN(new_n414));
  NOR3_X1   g213(.A1(new_n413), .A2(new_n414), .A3(new_n399), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n412), .A2(new_n415), .A3(KEYINPUT70), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT70), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n407), .A2(new_n408), .B1(new_n398), .B2(new_n399), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT69), .B(G127gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(G134gat), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n417), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n410), .B1(new_n416), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT23), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n423), .B1(G169gat), .B2(G176gat), .ZN(new_n424));
  AND2_X1   g223(.A1(G169gat), .A2(G176gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(G169gat), .A2(G176gat), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n425), .B1(KEYINPUT23), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT65), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n424), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G183gat), .A2(G190gat), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT24), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(KEYINPUT66), .A3(new_n431), .ZN(new_n432));
  OR2_X1    g231(.A1(G183gat), .A2(G190gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n431), .B1(new_n430), .B2(KEYINPUT66), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT25), .B1(new_n429), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT67), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT28), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(G190gat), .ZN(new_n441));
  AND2_X1   g240(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n442));
  NOR2_X1   g241(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n440), .B(new_n441), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT68), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT68), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n447), .A2(KEYINPUT67), .A3(KEYINPUT28), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n444), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT27), .B(G183gat), .ZN(new_n451));
  AOI21_X1  g250(.A(G190gat), .B1(new_n438), .B2(new_n439), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n451), .A2(new_n446), .A3(new_n448), .A4(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n425), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n426), .A2(KEYINPUT26), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT26), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n456), .A2(G169gat), .A3(G176gat), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n454), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n450), .A2(new_n453), .A3(new_n458), .A4(new_n430), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n437), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n427), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT25), .ZN(new_n462));
  NAND3_X1  g261(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n433), .B(new_n463), .C1(new_n464), .C2(KEYINPUT64), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(KEYINPUT64), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n462), .B(new_n424), .C1(new_n465), .C2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n462), .A2(KEYINPUT65), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n461), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n422), .B1(new_n460), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n444), .A2(new_n449), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n451), .A2(new_n452), .B1(new_n446), .B2(new_n448), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n458), .A2(new_n430), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n423), .A2(G169gat), .A3(G176gat), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT65), .B1(new_n477), .B2(new_n425), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n478), .B(new_n424), .C1(new_n435), .C2(new_n434), .ZN(new_n479));
  AOI22_X1  g278(.A1(new_n475), .A2(new_n476), .B1(new_n479), .B2(KEYINPUT25), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT70), .B1(new_n412), .B2(new_n415), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n418), .A2(new_n417), .A3(new_n420), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n409), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n424), .A2(new_n462), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n463), .B1(G183gat), .B2(G190gat), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT64), .B1(new_n430), .B2(new_n431), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n484), .B1(new_n487), .B2(new_n466), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n427), .B1(new_n488), .B2(new_n469), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n480), .A2(new_n483), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(G227gat), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n491), .A2(new_n338), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n472), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n494), .B(KEYINPUT34), .ZN(new_n495));
  XNOR2_X1  g294(.A(G15gat), .B(G43gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(G71gat), .B(G99gat), .ZN(new_n497));
  XOR2_X1   g296(.A(new_n496), .B(new_n497), .Z(new_n498));
  AOI21_X1  g297(.A(new_n493), .B1(new_n472), .B2(new_n490), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n498), .B1(new_n499), .B2(KEYINPUT33), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT32), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n472), .A2(new_n490), .ZN(new_n504));
  AOI221_X4 g303(.A(new_n501), .B1(KEYINPUT33), .B2(new_n498), .C1(new_n504), .C2(new_n492), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n495), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n492), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT32), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT33), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n508), .A2(new_n510), .A3(new_n498), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT34), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n494), .B(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n500), .A2(new_n502), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n511), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n495), .A2(KEYINPUT71), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n506), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  OAI211_X1 g316(.A(KEYINPUT71), .B(new_n495), .C1(new_n503), .C2(new_n505), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT36), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n515), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n522), .A2(KEYINPUT36), .ZN(new_n523));
  OR2_X1    g322(.A1(KEYINPUT72), .A2(G197gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(KEYINPUT72), .A2(G197gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(G204gat), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(G204gat), .ZN(new_n527));
  AND2_X1   g326(.A1(KEYINPUT72), .A2(G197gat), .ZN(new_n528));
  NOR2_X1   g327(.A1(KEYINPUT72), .A2(G197gat), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT22), .ZN(new_n531));
  INV_X1    g330(.A(G211gat), .ZN(new_n532));
  INV_X1    g331(.A(G218gat), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n526), .A2(new_n530), .A3(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G211gat), .B(G218gat), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n526), .A2(new_n530), .A3(new_n536), .A4(new_n534), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(G226gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n542), .A2(new_n338), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n489), .A2(new_n437), .A3(new_n459), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT29), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n543), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n547), .B1(new_n480), .B2(new_n489), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n541), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT74), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT73), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n551), .B1(new_n546), .B2(new_n548), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n545), .B1(new_n460), .B2(new_n471), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n551), .B1(new_n553), .B2(new_n547), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n550), .B1(new_n556), .B2(new_n541), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT30), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n544), .A2(new_n543), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT29), .B1(new_n480), .B2(new_n489), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n559), .B1(new_n560), .B2(new_n543), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n554), .B1(new_n561), .B2(new_n551), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n562), .A2(KEYINPUT74), .A3(new_n540), .ZN(new_n563));
  XNOR2_X1  g362(.A(G8gat), .B(G36gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(G64gat), .B(G92gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n557), .A2(new_n558), .A3(new_n563), .A4(new_n567), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n562), .A2(new_n540), .B1(KEYINPUT74), .B2(new_n549), .ZN(new_n569));
  AND4_X1   g368(.A1(KEYINPUT74), .A2(new_n552), .A3(new_n555), .A4(new_n540), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n566), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n557), .A2(new_n563), .A3(new_n567), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(KEYINPUT30), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G1gat), .B(G29gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(new_n279), .ZN(new_n575));
  XNOR2_X1  g374(.A(KEYINPUT0), .B(G57gat), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n575), .B(new_n576), .Z(new_n577));
  NAND2_X1  g376(.A1(G225gat), .A2(G233gat), .ZN(new_n578));
  XOR2_X1   g377(.A(G155gat), .B(G162gat), .Z(new_n579));
  XNOR2_X1  g378(.A(G141gat), .B(G148gat), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n579), .B1(KEYINPUT2), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT2), .ZN(new_n582));
  AND2_X1   g381(.A1(KEYINPUT75), .A2(G155gat), .ZN(new_n583));
  NOR2_X1   g382(.A1(KEYINPUT75), .A2(G155gat), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n582), .B1(new_n585), .B2(G162gat), .ZN(new_n586));
  OR2_X1    g385(.A1(G155gat), .A2(G162gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(G155gat), .A2(G162gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(G148gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(G141gat), .ZN(new_n591));
  INV_X1    g390(.A(G141gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(G148gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n581), .B1(new_n586), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n422), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT75), .B(G155gat), .ZN(new_n598));
  OAI21_X1  g397(.A(KEYINPUT2), .B1(new_n598), .B2(new_n311), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n591), .A2(new_n593), .B1(new_n587), .B2(new_n588), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n594), .A2(new_n582), .ZN(new_n601));
  AOI22_X1  g400(.A1(new_n599), .A2(new_n600), .B1(new_n601), .B2(new_n579), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n410), .B(new_n602), .C1(new_n416), .C2(new_n421), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n578), .B1(new_n597), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT5), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT78), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n578), .ZN(new_n607));
  INV_X1    g406(.A(new_n603), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n481), .A2(new_n482), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n602), .B1(new_n609), .B2(new_n410), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n607), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT78), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(new_n612), .A3(KEYINPUT5), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT4), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n607), .B1(new_n603), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT77), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n602), .A2(new_n616), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n581), .B(new_n616), .C1(new_n586), .C2(new_n595), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n483), .B(KEYINPUT4), .C1(new_n617), .C2(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n596), .A2(KEYINPUT3), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT3), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n581), .B(new_n623), .C1(new_n586), .C2(new_n595), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(KEYINPUT76), .B1(new_n625), .B2(new_n483), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT76), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n422), .A2(new_n627), .A3(new_n624), .A4(new_n622), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  AOI22_X1  g428(.A1(new_n606), .A2(new_n613), .B1(new_n621), .B2(new_n629), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n483), .B(new_n614), .C1(new_n617), .C2(new_n619), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n603), .A2(KEYINPUT4), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT79), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n631), .A2(new_n632), .A3(KEYINPUT79), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n607), .A2(KEYINPUT5), .ZN(new_n637));
  AND4_X1   g436(.A1(new_n629), .A2(new_n635), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n577), .B1(new_n630), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT6), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n621), .A2(new_n629), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n604), .A2(KEYINPUT78), .A3(new_n605), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n612), .B1(new_n611), .B2(KEYINPUT5), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n577), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n635), .A2(new_n629), .A3(new_n636), .A4(new_n637), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n639), .A2(new_n640), .A3(new_n647), .ZN(new_n648));
  OAI211_X1 g447(.A(KEYINPUT6), .B(new_n577), .C1(new_n630), .C2(new_n638), .ZN(new_n649));
  AOI22_X1  g448(.A1(new_n568), .A2(new_n573), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT29), .B1(new_n538), .B2(new_n539), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n623), .B1(new_n651), .B2(KEYINPUT80), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT80), .ZN(new_n653));
  AOI211_X1 g452(.A(new_n653), .B(KEYINPUT29), .C1(new_n538), .C2(new_n539), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n596), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(G228gat), .A2(G233gat), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n624), .A2(new_n545), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n656), .B1(new_n541), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(G22gat), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n596), .A2(KEYINPUT77), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n661), .B(new_n618), .C1(new_n651), .C2(KEYINPUT3), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n541), .A2(new_n657), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n656), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n659), .A2(new_n660), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(KEYINPUT82), .ZN(new_n667));
  AOI22_X1  g466(.A1(new_n655), .A2(new_n658), .B1(new_n664), .B2(new_n656), .ZN(new_n668));
  OAI21_X1  g467(.A(G22gat), .B1(new_n668), .B2(KEYINPUT81), .ZN(new_n669));
  INV_X1    g468(.A(new_n656), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n663), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n540), .A2(new_n545), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n653), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n651), .A2(KEYINPUT80), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n673), .A2(new_n623), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n671), .B1(new_n675), .B2(new_n596), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT81), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n670), .B1(new_n662), .B2(new_n663), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n667), .B1(new_n669), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(G78gat), .B(G106gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT31), .B(G50gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n668), .A2(KEYINPUT81), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n677), .B1(new_n676), .B2(new_n678), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n684), .A2(new_n685), .A3(KEYINPUT82), .A4(G22gat), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n680), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n683), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n668), .A2(new_n660), .ZN(new_n689));
  INV_X1    g488(.A(new_n666), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n521), .B(new_n523), .C1(new_n650), .C2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n692), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT39), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n608), .A2(new_n610), .A3(new_n607), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n635), .A2(new_n629), .A3(new_n636), .ZN(new_n698));
  AOI211_X1 g497(.A(new_n696), .B(new_n697), .C1(new_n698), .C2(new_n607), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(new_n696), .A3(new_n607), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n577), .B(KEYINPUT83), .Z(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(KEYINPUT40), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT84), .B1(new_n630), .B2(new_n638), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT84), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n644), .A2(new_n707), .A3(new_n646), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n702), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT40), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n699), .A2(new_n703), .A3(new_n710), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n705), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n573), .A2(new_n568), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n695), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n569), .A2(new_n570), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT37), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n567), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n562), .A2(new_n541), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n718), .B1(new_n561), .B2(new_n540), .ZN(new_n721));
  AOI21_X1  g520(.A(KEYINPUT38), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n572), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n647), .A2(new_n640), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n649), .B1(new_n709), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT38), .ZN(new_n727));
  OAI21_X1  g526(.A(KEYINPUT37), .B1(new_n569), .B2(new_n570), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n727), .B1(new_n719), .B2(new_n728), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n724), .A2(new_n726), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n694), .B1(new_n716), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n695), .A2(new_n522), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT35), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n732), .A2(new_n726), .A3(new_n733), .A4(new_n713), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT85), .ZN(new_n735));
  AOI22_X1  g534(.A1(new_n518), .A2(new_n517), .B1(new_n687), .B2(new_n691), .ZN(new_n736));
  AOI211_X1 g535(.A(new_n735), .B(new_n733), .C1(new_n650), .C2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n648), .A2(new_n649), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n713), .A2(new_n738), .A3(new_n692), .A4(new_n519), .ZN(new_n739));
  AOI21_X1  g538(.A(KEYINPUT85), .B1(new_n739), .B2(KEYINPUT35), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n734), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  AOI211_X1 g540(.A(new_n277), .B(new_n397), .C1(new_n731), .C2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n738), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g544(.A1(new_n742), .A2(new_n714), .ZN(new_n746));
  OAI21_X1  g545(.A(KEYINPUT42), .B1(new_n746), .B2(new_n228), .ZN(new_n747));
  XOR2_X1   g546(.A(KEYINPUT16), .B(G8gat), .Z(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  MUX2_X1   g548(.A(KEYINPUT42), .B(new_n747), .S(new_n749), .Z(G1325gat));
  INV_X1    g549(.A(new_n522), .ZN(new_n751));
  AOI21_X1  g550(.A(G15gat), .B1(new_n742), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n521), .A2(new_n523), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n753), .A2(G15gat), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n752), .B1(new_n742), .B2(new_n754), .ZN(G1326gat));
  NAND2_X1  g554(.A1(new_n742), .A2(new_n695), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT106), .ZN(new_n757));
  XOR2_X1   g556(.A(KEYINPUT43), .B(G22gat), .Z(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(G1327gat));
  AOI21_X1  g558(.A(new_n316), .B1(new_n731), .B2(new_n741), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n760), .A2(KEYINPUT44), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n739), .A2(KEYINPUT35), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n735), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n739), .A2(KEYINPUT85), .A3(KEYINPUT35), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT108), .B1(new_n765), .B2(new_n734), .ZN(new_n766));
  OAI211_X1 g565(.A(KEYINPUT108), .B(new_n734), .C1(new_n737), .C2(new_n740), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n731), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n317), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n761), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n396), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n277), .A2(new_n369), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(G29gat), .B1(new_n775), .B2(new_n738), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n774), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n777), .A2(G29gat), .A3(new_n738), .ZN(new_n778));
  XNOR2_X1  g577(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n776), .A2(new_n780), .ZN(G1328gat));
  OAI21_X1  g580(.A(new_n202), .B1(new_n775), .B2(new_n713), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n777), .A2(new_n713), .A3(new_n202), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT46), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n785), .A2(KEYINPUT109), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n783), .A2(new_n784), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(KEYINPUT109), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n782), .A2(new_n786), .A3(new_n787), .A4(new_n788), .ZN(G1329gat));
  INV_X1    g588(.A(new_n730), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n693), .B1(new_n790), .B2(new_n715), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT108), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n741), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n791), .B1(new_n793), .B2(new_n767), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n771), .B1(new_n794), .B2(new_n316), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n760), .A2(KEYINPUT44), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n795), .A2(new_n753), .A3(new_n796), .A4(new_n774), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(G43gat), .ZN(new_n798));
  INV_X1    g597(.A(new_n777), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n799), .A2(new_n206), .A3(new_n751), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT47), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n801), .B(new_n802), .ZN(G1330gat));
  NAND4_X1  g602(.A1(new_n795), .A2(new_n695), .A3(new_n796), .A4(new_n774), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(G50gat), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n799), .A2(new_n204), .A3(new_n695), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT48), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n807), .B(new_n808), .ZN(G1331gat));
  AND2_X1   g608(.A1(new_n368), .A2(new_n371), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n810), .A2(new_n277), .A3(new_n773), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n794), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n743), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(G57gat), .ZN(G1332gat));
  INV_X1    g613(.A(KEYINPUT49), .ZN(new_n815));
  INV_X1    g614(.A(G64gat), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n714), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(KEYINPUT110), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n812), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n815), .A2(new_n816), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n819), .B(new_n820), .ZN(G1333gat));
  NAND2_X1  g620(.A1(new_n812), .A2(new_n753), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n522), .A2(G71gat), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n822), .A2(G71gat), .B1(new_n812), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g624(.A1(new_n812), .A2(new_n695), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(G78gat), .ZN(G1335gat));
  INV_X1    g626(.A(new_n277), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(new_n369), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(new_n396), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n772), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n832), .A2(new_n738), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n793), .A2(new_n767), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n316), .B1(new_n834), .B2(new_n731), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT51), .B1(new_n835), .B2(new_n829), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n769), .A2(KEYINPUT51), .A3(new_n317), .A4(new_n829), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT111), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT111), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n835), .A2(new_n839), .A3(KEYINPUT51), .A4(new_n829), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n836), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n743), .A2(new_n773), .A3(new_n292), .ZN(new_n842));
  OAI22_X1  g641(.A1(new_n833), .A2(new_n292), .B1(new_n841), .B2(new_n842), .ZN(G1336gat));
  NAND3_X1  g642(.A1(new_n714), .A2(new_n280), .A3(new_n773), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n838), .A2(new_n840), .ZN(new_n845));
  XOR2_X1   g644(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n846));
  OAI21_X1  g645(.A(new_n846), .B1(new_n770), .B2(new_n830), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n844), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n795), .A2(new_n714), .A3(new_n796), .A4(new_n831), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n849), .A2(G92gat), .ZN(new_n850));
  OAI21_X1  g649(.A(KEYINPUT52), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT52), .B1(new_n849), .B2(G92gat), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n852), .B1(new_n841), .B2(new_n844), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(G1337gat));
  XOR2_X1   g653(.A(KEYINPUT113), .B(G99gat), .Z(new_n855));
  INV_X1    g654(.A(new_n753), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n832), .B2(new_n856), .ZN(new_n857));
  OR3_X1    g656(.A1(new_n396), .A2(new_n522), .A3(new_n855), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n857), .B1(new_n841), .B2(new_n858), .ZN(G1338gat));
  NAND4_X1  g658(.A1(new_n795), .A2(new_n695), .A3(new_n796), .A4(new_n831), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n860), .A2(G106gat), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n847), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n396), .A2(new_n692), .A3(G106gat), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n865));
  INV_X1    g664(.A(G106gat), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n866), .B1(new_n860), .B2(new_n867), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n772), .A2(KEYINPUT114), .A3(new_n695), .A4(new_n831), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n863), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n865), .B1(new_n841), .B2(new_n871), .ZN(new_n872));
  OAI22_X1  g671(.A1(new_n864), .A2(new_n865), .B1(new_n870), .B2(new_n872), .ZN(G1339gat));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n874), .B1(new_n390), .B2(new_n393), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n874), .B1(new_n378), .B2(new_n379), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n376), .A2(new_n377), .A3(new_n382), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n387), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT55), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n875), .A2(new_n878), .A3(KEYINPUT55), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(new_n388), .A3(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n884), .B1(new_n271), .B2(new_n276), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n250), .A2(new_n254), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(G229gat), .A3(G233gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n250), .A2(new_n234), .A3(new_n242), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n260), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT93), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n264), .A2(new_n265), .A3(new_n267), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n244), .A2(new_n255), .A3(new_n261), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n262), .A2(KEYINPUT93), .A3(new_n268), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n889), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(new_n773), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n317), .B1(new_n885), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n895), .A2(new_n884), .A3(new_n317), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n367), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n828), .A2(new_n397), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n903), .A2(new_n732), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n714), .A2(new_n738), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(G113gat), .B1(new_n906), .B2(new_n277), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n268), .A2(new_n273), .ZN(new_n908));
  INV_X1    g707(.A(new_n272), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n909), .A3(new_n275), .ZN(new_n910));
  INV_X1    g709(.A(new_n261), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n893), .A2(new_n894), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n883), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI211_X1 g713(.A(new_n396), .B(new_n889), .C1(new_n893), .C2(new_n894), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n316), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n369), .B1(new_n916), .B2(new_n898), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n917), .A2(new_n901), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n905), .A2(new_n736), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(new_n405), .A3(new_n828), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n907), .A2(new_n921), .ZN(G1340gat));
  OAI21_X1  g721(.A(G120gat), .B1(new_n906), .B2(new_n396), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n920), .A2(new_n403), .A3(new_n773), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(G1341gat));
  AOI21_X1  g724(.A(new_n419), .B1(new_n920), .B2(new_n369), .ZN(new_n926));
  INV_X1    g725(.A(new_n906), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n367), .A2(new_n413), .A3(new_n414), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(G1342gat));
  INV_X1    g728(.A(KEYINPUT115), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n920), .A2(new_n399), .A3(new_n317), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT56), .ZN(new_n932));
  OAI21_X1  g731(.A(G134gat), .B1(new_n906), .B2(new_n316), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n930), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n931), .A2(KEYINPUT56), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n931), .A2(KEYINPUT56), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n936), .A2(KEYINPUT115), .A3(new_n933), .A4(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n935), .A2(new_n938), .ZN(G1343gat));
  INV_X1    g738(.A(KEYINPUT58), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n918), .A2(new_n692), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n753), .A2(new_n738), .A3(new_n714), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n943), .A2(G141gat), .A3(new_n277), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  XOR2_X1   g744(.A(new_n942), .B(KEYINPUT116), .Z(new_n946));
  AOI21_X1  g745(.A(new_n899), .B1(new_n916), .B2(KEYINPUT118), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT118), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n897), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n369), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  OAI211_X1 g749(.A(KEYINPUT57), .B(new_n695), .C1(new_n950), .C2(new_n901), .ZN(new_n951));
  XOR2_X1   g750(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n953), .B1(new_n918), .B2(new_n692), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n946), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n955), .A2(new_n828), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n940), .B(new_n945), .C1(new_n956), .C2(new_n592), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n592), .B1(new_n955), .B2(new_n828), .ZN(new_n958));
  OAI21_X1  g757(.A(KEYINPUT58), .B1(new_n958), .B2(new_n944), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n959), .ZN(G1344gat));
  INV_X1    g759(.A(new_n943), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n961), .A2(new_n590), .A3(new_n773), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT59), .ZN(new_n963));
  OAI21_X1  g762(.A(KEYINPUT120), .B1(new_n883), .B2(new_n316), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT120), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n389), .B1(new_n879), .B2(new_n880), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n317), .A2(new_n965), .A3(new_n882), .A4(new_n966), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n964), .A2(new_n895), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n367), .B1(new_n897), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n692), .B1(new_n969), .B2(new_n902), .ZN(new_n970));
  OAI21_X1  g769(.A(KEYINPUT121), .B1(new_n970), .B2(KEYINPUT57), .ZN(new_n971));
  OAI211_X1 g770(.A(new_n695), .B(new_n952), .C1(new_n917), .C2(new_n901), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT119), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT121), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT57), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n964), .A2(new_n895), .A3(new_n967), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n916), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n901), .B1(new_n978), .B2(new_n367), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n975), .B(new_n976), .C1(new_n979), .C2(new_n692), .ZN(new_n980));
  NAND4_X1  g779(.A1(new_n903), .A2(KEYINPUT119), .A3(new_n695), .A4(new_n952), .ZN(new_n981));
  NAND4_X1  g780(.A1(new_n971), .A2(new_n974), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  INV_X1    g781(.A(new_n946), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n982), .A2(new_n773), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n963), .B1(new_n984), .B2(G148gat), .ZN(new_n985));
  AOI211_X1 g784(.A(KEYINPUT59), .B(new_n590), .C1(new_n955), .C2(new_n773), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n962), .B1(new_n985), .B2(new_n986), .ZN(G1345gat));
  AOI21_X1  g786(.A(new_n585), .B1(new_n961), .B2(new_n369), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n367), .A2(new_n598), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n988), .B1(new_n955), .B2(new_n989), .ZN(G1346gat));
  AOI21_X1  g789(.A(G162gat), .B1(new_n961), .B2(new_n317), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n316), .A2(new_n311), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n991), .B1(new_n955), .B2(new_n992), .ZN(G1347gat));
  NOR2_X1   g792(.A1(new_n918), .A2(new_n743), .ZN(new_n994));
  NOR3_X1   g793(.A1(new_n520), .A2(new_n695), .A3(new_n713), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NOR3_X1   g795(.A1(new_n996), .A2(G169gat), .A3(new_n277), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n997), .B(KEYINPUT122), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n714), .A2(new_n738), .ZN(new_n999));
  XNOR2_X1  g798(.A(new_n999), .B(KEYINPUT123), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n904), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g800(.A(G169gat), .B1(new_n1001), .B2(new_n277), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n998), .A2(new_n1002), .ZN(G1348gat));
  OAI21_X1  g802(.A(G176gat), .B1(new_n1001), .B2(new_n396), .ZN(new_n1004));
  INV_X1    g803(.A(G176gat), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n773), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1004), .B1(new_n996), .B2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g806(.A(new_n1007), .B(KEYINPUT124), .ZN(G1349gat));
  OAI21_X1  g807(.A(G183gat), .B1(new_n1001), .B2(new_n367), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n369), .A2(new_n451), .ZN(new_n1010));
  OAI21_X1  g809(.A(new_n1009), .B1(new_n996), .B2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g810(.A(new_n1011), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g811(.A(G190gat), .B1(new_n1001), .B2(new_n316), .ZN(new_n1013));
  AND2_X1   g812(.A1(new_n1013), .A2(KEYINPUT61), .ZN(new_n1014));
  NOR2_X1   g813(.A1(new_n1013), .A2(KEYINPUT61), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n317), .A2(new_n441), .ZN(new_n1016));
  OAI22_X1  g815(.A1(new_n1014), .A2(new_n1015), .B1(new_n996), .B2(new_n1016), .ZN(G1351gat));
  NAND3_X1  g816(.A1(new_n856), .A2(new_n714), .A3(new_n695), .ZN(new_n1018));
  XNOR2_X1  g817(.A(new_n1018), .B(KEYINPUT125), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n994), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g819(.A(new_n1020), .ZN(new_n1021));
  NAND3_X1  g820(.A1(new_n1021), .A2(new_n257), .A3(new_n828), .ZN(new_n1022));
  AND2_X1   g821(.A1(new_n1000), .A2(new_n856), .ZN(new_n1023));
  AND3_X1   g822(.A1(new_n982), .A2(new_n828), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g823(.A(new_n1022), .B1(new_n1024), .B2(new_n257), .ZN(G1352gat));
  NAND2_X1  g824(.A1(new_n773), .A2(new_n527), .ZN(new_n1026));
  OAI21_X1  g825(.A(KEYINPUT62), .B1(new_n1020), .B2(new_n1026), .ZN(new_n1027));
  OR3_X1    g826(.A1(new_n1020), .A2(KEYINPUT62), .A3(new_n1026), .ZN(new_n1028));
  AND3_X1   g827(.A1(new_n982), .A2(new_n773), .A3(new_n1023), .ZN(new_n1029));
  OAI211_X1 g828(.A(new_n1027), .B(new_n1028), .C1(new_n1029), .C2(new_n527), .ZN(G1353gat));
  NAND3_X1  g829(.A1(new_n1021), .A2(new_n532), .A3(new_n369), .ZN(new_n1031));
  NAND3_X1  g830(.A1(new_n982), .A2(new_n369), .A3(new_n1023), .ZN(new_n1032));
  AND3_X1   g831(.A1(new_n1032), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1033));
  AOI21_X1  g832(.A(KEYINPUT63), .B1(new_n1032), .B2(G211gat), .ZN(new_n1034));
  OAI21_X1  g833(.A(new_n1031), .B1(new_n1033), .B2(new_n1034), .ZN(G1354gat));
  NAND2_X1  g834(.A1(new_n317), .A2(G218gat), .ZN(new_n1036));
  XNOR2_X1  g835(.A(new_n1036), .B(KEYINPUT126), .ZN(new_n1037));
  NAND3_X1  g836(.A1(new_n982), .A2(new_n1023), .A3(new_n1037), .ZN(new_n1038));
  OAI21_X1  g837(.A(new_n533), .B1(new_n1020), .B2(new_n316), .ZN(new_n1039));
  AND2_X1   g838(.A1(new_n1038), .A2(new_n1039), .ZN(G1355gat));
endmodule


