//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n627, new_n628, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n791, new_n792, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n848, new_n849, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT5), .ZN(new_n203));
  NAND2_X1  g002(.A1(G225gat), .A2(G233gat), .ZN(new_n204));
  XOR2_X1   g003(.A(G127gat), .B(G134gat), .Z(new_n205));
  INV_X1    g004(.A(KEYINPUT1), .ZN(new_n206));
  XNOR2_X1  g005(.A(G113gat), .B(G120gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT67), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G113gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G120gat), .ZN(new_n211));
  INV_X1    g010(.A(G120gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G113gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n213), .A3(new_n208), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n205), .B1(new_n209), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT69), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n211), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n210), .A2(KEYINPUT69), .A3(G120gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT68), .B(G120gat), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n218), .B(new_n219), .C1(new_n220), .C2(new_n210), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n205), .A2(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n216), .A2(new_n223), .ZN(new_n224));
  OR2_X1    g023(.A1(G141gat), .A2(G148gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(G141gat), .A2(G148gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(KEYINPUT77), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT77), .ZN(new_n228));
  AND2_X1   g027(.A1(G141gat), .A2(G148gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(G141gat), .A2(G148gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G155gat), .A2(G162gat), .ZN(new_n232));
  OR3_X1    g031(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n227), .A2(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G155gat), .ZN(new_n235));
  INV_X1    g034(.A(G162gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(new_n232), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n229), .A2(new_n230), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT76), .B(KEYINPUT2), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  OAI211_X1 g040(.A(KEYINPUT78), .B(KEYINPUT3), .C1(new_n234), .C2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n231), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n233), .A2(new_n232), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n239), .A2(new_n240), .ZN(new_n247));
  INV_X1    g046(.A(new_n238), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n245), .A2(new_n246), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n224), .A2(new_n242), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n245), .A2(new_n249), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT78), .B1(new_n252), .B2(KEYINPUT3), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n203), .B(new_n204), .C1(new_n251), .C2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n243), .A2(new_n244), .B1(new_n247), .B2(new_n248), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n256), .A2(new_n216), .A3(new_n223), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT80), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(new_n258), .A3(KEYINPUT4), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(KEYINPUT4), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n211), .A2(new_n213), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT67), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n262), .A2(new_n206), .A3(new_n214), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n263), .A2(new_n205), .B1(new_n221), .B2(new_n222), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(new_n265), .A3(new_n256), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n260), .A2(new_n266), .A3(KEYINPUT80), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n255), .A2(new_n259), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n224), .A2(new_n252), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(new_n257), .ZN(new_n270));
  INV_X1    g069(.A(new_n204), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n203), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n260), .A2(KEYINPUT79), .A3(new_n266), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT79), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n264), .A2(new_n274), .A3(new_n265), .A4(new_n256), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n275), .B(new_n204), .C1(new_n251), .C2(new_n253), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n272), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n268), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G1gat), .B(G29gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT0), .ZN(new_n280));
  XNOR2_X1  g079(.A(G57gat), .B(G85gat), .ZN(new_n281));
  XOR2_X1   g080(.A(new_n280), .B(new_n281), .Z(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n278), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n268), .A2(new_n277), .A3(new_n282), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT81), .ZN(new_n288));
  AND4_X1   g087(.A1(new_n288), .A2(new_n278), .A3(KEYINPUT6), .A4(new_n283), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n282), .B1(new_n268), .B2(new_n277), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n288), .B1(new_n290), .B2(KEYINPUT6), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n287), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G8gat), .B(G36gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(G64gat), .B(G92gat), .ZN(new_n294));
  XOR2_X1   g093(.A(new_n293), .B(new_n294), .Z(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G226gat), .ZN(new_n297));
  INV_X1    g096(.A(G233gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AND2_X1   g098(.A1(G183gat), .A2(G190gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT24), .ZN(new_n301));
  AOI22_X1  g100(.A1(new_n300), .A2(new_n301), .B1(G169gat), .B2(G176gat), .ZN(new_n302));
  INV_X1    g101(.A(G183gat), .ZN(new_n303));
  INV_X1    g102(.A(G190gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G183gat), .A2(G190gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(KEYINPUT24), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G169gat), .ZN(new_n308));
  INV_X1    g107(.A(G176gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT23), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT23), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n302), .A2(new_n307), .A3(new_n312), .A4(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT25), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT64), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n315), .A2(KEYINPUT64), .A3(new_n316), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT65), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n313), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n322), .A2(KEYINPUT23), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT25), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n302), .A2(new_n307), .A3(new_n312), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n319), .A2(new_n320), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT26), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n322), .A2(new_n331), .A3(new_n323), .ZN(new_n332));
  NAND2_X1  g131(.A1(G169gat), .A2(G176gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n310), .A2(KEYINPUT26), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(new_n306), .ZN(new_n336));
  NAND2_X1  g135(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n337));
  AOI21_X1  g136(.A(G190gat), .B1(new_n337), .B2(KEYINPUT27), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT27), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n339), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT28), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT27), .B(G183gat), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n304), .A2(KEYINPUT28), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n336), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT29), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n299), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT64), .B1(new_n315), .B2(new_n316), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n325), .A2(new_n327), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n345), .B1(new_n352), .B2(new_n320), .ZN(new_n353));
  INV_X1    g152(.A(new_n299), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G197gat), .B(G204gat), .ZN(new_n356));
  INV_X1    g155(.A(G211gat), .ZN(new_n357));
  INV_X1    g156(.A(G218gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n356), .B1(KEYINPUT22), .B2(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G211gat), .B(G218gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n349), .A2(new_n355), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n362), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n354), .B1(new_n353), .B2(KEYINPUT29), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n347), .A2(new_n299), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n296), .B1(new_n363), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT75), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n362), .B1(new_n349), .B2(new_n355), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n365), .A2(new_n364), .A3(new_n366), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n373), .A2(KEYINPUT75), .A3(new_n296), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n371), .A2(new_n372), .A3(new_n295), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT30), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT30), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n371), .A2(new_n372), .A3(new_n377), .A4(new_n295), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n370), .A2(new_n374), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT82), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n292), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n380), .B1(new_n292), .B2(new_n379), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n315), .A2(KEYINPUT64), .A3(new_n316), .ZN(new_n383));
  NOR3_X1   g182(.A1(new_n383), .A2(new_n350), .A3(new_n351), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n264), .B1(new_n384), .B2(new_n345), .ZN(new_n385));
  INV_X1    g184(.A(G227gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n386), .A2(new_n298), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n330), .A2(new_n346), .A3(new_n224), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n385), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT32), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT33), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  XOR2_X1   g191(.A(G15gat), .B(G43gat), .Z(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT70), .ZN(new_n394));
  XOR2_X1   g193(.A(G71gat), .B(G99gat), .Z(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n390), .A2(new_n392), .A3(new_n397), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n389), .B(KEYINPUT32), .C1(new_n391), .C2(new_n396), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n353), .A2(new_n224), .ZN(new_n403));
  INV_X1    g202(.A(new_n388), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n402), .B1(new_n405), .B2(new_n387), .ZN(new_n406));
  OAI221_X1 g205(.A(new_n401), .B1(new_n386), .B2(new_n298), .C1(new_n403), .C2(new_n404), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n400), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT72), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n398), .A2(new_n399), .A3(new_n406), .A4(new_n407), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT72), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n400), .A2(new_n412), .A3(new_n408), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n364), .A2(new_n348), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n256), .B1(new_n414), .B2(new_n246), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n364), .B1(new_n348), .B2(new_n250), .ZN(new_n416));
  XNOR2_X1  g215(.A(G78gat), .B(G106gat), .ZN(new_n417));
  OR3_X1    g216(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n417), .B1(new_n415), .B2(new_n416), .ZN(new_n419));
  NAND2_X1  g218(.A1(G228gat), .A2(G233gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(G22gat), .ZN(new_n421));
  XOR2_X1   g220(.A(KEYINPUT31), .B(G50gat), .Z(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n418), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n423), .B1(new_n418), .B2(new_n419), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n410), .A2(new_n411), .A3(new_n413), .A4(new_n426), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n381), .A2(new_n382), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT35), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n202), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n291), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n290), .A2(new_n288), .A3(KEYINPUT6), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n290), .A2(KEYINPUT6), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n431), .A2(new_n432), .B1(new_n286), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n370), .A2(new_n374), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n376), .A2(new_n378), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT82), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n292), .A2(new_n379), .A3(new_n380), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(KEYINPUT85), .B(KEYINPUT35), .C1(new_n440), .C2(new_n427), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n437), .A2(KEYINPUT83), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT83), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n379), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n409), .A2(KEYINPUT73), .A3(new_n411), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT73), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n400), .A2(new_n447), .A3(new_n408), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n426), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n450), .A2(KEYINPUT35), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n445), .A2(new_n449), .A3(new_n292), .A4(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n430), .A2(new_n441), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n434), .A2(new_n375), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n373), .A2(KEYINPUT37), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT37), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n371), .A2(new_n372), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(new_n296), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT38), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n459), .B1(new_n457), .B2(KEYINPUT84), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n458), .B(new_n460), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n267), .B(new_n259), .C1(new_n253), .C2(new_n251), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n271), .ZN(new_n463));
  OR2_X1    g262(.A1(new_n463), .A2(KEYINPUT39), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n463), .B(KEYINPUT39), .C1(new_n271), .C2(new_n270), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(new_n465), .A3(new_n282), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT40), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n290), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n468), .B1(new_n467), .B2(new_n466), .ZN(new_n469));
  OAI221_X1 g268(.A(new_n426), .B1(new_n454), .B2(new_n461), .C1(new_n445), .C2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT74), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n471), .B1(new_n449), .B2(KEYINPUT36), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT36), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n446), .A2(KEYINPUT74), .A3(new_n473), .A4(new_n448), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n410), .A2(KEYINPUT36), .A3(new_n411), .A4(new_n413), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n450), .B1(new_n381), .B2(new_n382), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n470), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n453), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(G15gat), .B(G22gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n480), .B(KEYINPUT88), .ZN(new_n481));
  INV_X1    g280(.A(G1gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n482), .A2(KEYINPUT16), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n483), .B(KEYINPUT89), .C1(new_n481), .C2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(G8gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(G71gat), .B(G78gat), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n489), .B1(KEYINPUT91), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(G64gat), .ZN(new_n492));
  OR2_X1    g291(.A1(new_n492), .A2(G57gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(G57gat), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n491), .B(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(new_n496), .B(KEYINPUT94), .Z(new_n497));
  AOI21_X1  g296(.A(new_n488), .B1(KEYINPUT21), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n496), .A2(KEYINPUT21), .ZN(new_n499));
  XNOR2_X1  g298(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n498), .B(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(G127gat), .B(G155gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n503), .B(KEYINPUT93), .ZN(new_n504));
  NAND2_X1  g303(.A1(G231gat), .A2(G233gat), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n505), .B(KEYINPUT92), .Z(new_n506));
  XNOR2_X1  g305(.A(new_n504), .B(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G183gat), .B(G211gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n502), .B(new_n509), .ZN(new_n510));
  AND2_X1   g309(.A1(G232gat), .A2(G233gat), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n511), .A2(KEYINPUT41), .ZN(new_n512));
  XNOR2_X1  g311(.A(G134gat), .B(G162gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(G29gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n516), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n517));
  XOR2_X1   g316(.A(KEYINPUT14), .B(G29gat), .Z(new_n518));
  OAI21_X1  g317(.A(new_n517), .B1(new_n518), .B2(G36gat), .ZN(new_n519));
  AND2_X1   g318(.A1(G43gat), .A2(G50gat), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n520), .A2(KEYINPUT15), .ZN(new_n521));
  XNOR2_X1  g320(.A(KEYINPUT86), .B(G43gat), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n521), .B1(new_n522), .B2(G50gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(G43gat), .A2(G50gat), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT15), .B1(new_n520), .B2(new_n524), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n519), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT87), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n519), .A2(new_n525), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n529), .A2(KEYINPUT87), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n528), .B1(new_n530), .B2(new_n526), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n532), .ZN(new_n534));
  NAND2_X1  g333(.A1(G99gat), .A2(G106gat), .ZN(new_n535));
  INV_X1    g334(.A(G85gat), .ZN(new_n536));
  INV_X1    g335(.A(G92gat), .ZN(new_n537));
  AOI22_X1  g336(.A1(KEYINPUT8), .A2(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(KEYINPUT95), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(KEYINPUT95), .A2(G85gat), .A3(G92gat), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT7), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n538), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(G99gat), .B(G106gat), .Z(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n533), .A2(new_n534), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n545), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n531), .A2(new_n547), .B1(KEYINPUT41), .B2(new_n511), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G190gat), .B(G218gat), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n550), .B(KEYINPUT96), .Z(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n549), .A2(new_n551), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n515), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n554), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n556), .A2(new_n514), .A3(new_n552), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n510), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n488), .A2(new_n531), .ZN(new_n561));
  NAND2_X1  g360(.A1(G229gat), .A2(G233gat), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n533), .A2(new_n487), .A3(new_n534), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT90), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT18), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n487), .B(new_n531), .Z(new_n568));
  XOR2_X1   g367(.A(new_n562), .B(KEYINPUT13), .Z(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n565), .A2(new_n566), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n561), .A2(new_n562), .A3(new_n563), .A4(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n567), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G113gat), .B(G141gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(G197gat), .ZN(new_n575));
  XOR2_X1   g374(.A(KEYINPUT11), .B(G169gat), .Z(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n577), .B(KEYINPUT12), .Z(new_n578));
  NAND2_X1  g377(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n578), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n567), .A2(new_n570), .A3(new_n580), .A4(new_n572), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n497), .A2(KEYINPUT10), .A3(new_n547), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n543), .A2(new_n544), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n496), .B1(KEYINPUT97), .B2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(new_n545), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n584), .B1(KEYINPUT10), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G230gat), .A2(G233gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(G120gat), .B(G148gat), .Z(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT99), .ZN(new_n592));
  XOR2_X1   g391(.A(G176gat), .B(G204gat), .Z(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n586), .B(new_n547), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n595), .A2(new_n589), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n594), .B1(new_n596), .B2(KEYINPUT98), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n587), .A2(G230gat), .A3(G233gat), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT98), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n590), .A2(new_n597), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT100), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT100), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n590), .A2(new_n597), .A3(new_n603), .A4(new_n600), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n589), .B(KEYINPUT101), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n588), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(new_n598), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(new_n594), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  NOR3_X1   g410(.A1(new_n560), .A2(new_n583), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n479), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n613), .A2(new_n292), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(new_n482), .ZN(G1324gat));
  INV_X1    g414(.A(new_n613), .ZN(new_n616));
  INV_X1    g415(.A(new_n445), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n486), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(KEYINPUT16), .B(G8gat), .ZN(new_n619));
  NOR3_X1   g418(.A1(new_n613), .A2(new_n445), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(KEYINPUT42), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n621), .B1(KEYINPUT42), .B2(new_n620), .ZN(G1325gat));
  OAI21_X1  g421(.A(G15gat), .B1(new_n613), .B2(new_n476), .ZN(new_n623));
  INV_X1    g422(.A(G15gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n449), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n623), .B1(new_n613), .B2(new_n625), .ZN(G1326gat));
  NOR2_X1   g425(.A1(new_n613), .A2(new_n426), .ZN(new_n627));
  XOR2_X1   g426(.A(KEYINPUT43), .B(G22gat), .Z(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(G1327gat));
  AOI21_X1  g428(.A(new_n559), .B1(new_n453), .B2(new_n478), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n583), .A2(new_n510), .A3(new_n611), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n630), .A2(new_n516), .A3(new_n434), .A4(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT45), .ZN(new_n633));
  INV_X1    g432(.A(new_n631), .ZN(new_n634));
  XOR2_X1   g433(.A(KEYINPUT102), .B(KEYINPUT44), .Z(new_n635));
  AOI21_X1  g434(.A(new_n635), .B1(new_n479), .B2(new_n558), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT102), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT44), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI211_X1 g439(.A(new_n559), .B(new_n640), .C1(new_n453), .C2(new_n478), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n634), .B1(new_n637), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(new_n292), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n645), .A2(KEYINPUT103), .ZN(new_n646));
  OAI21_X1  g445(.A(G29gat), .B1(new_n645), .B2(KEYINPUT103), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n633), .B1(new_n646), .B2(new_n647), .ZN(G1328gat));
  OAI21_X1  g447(.A(G36gat), .B1(new_n644), .B2(new_n445), .ZN(new_n649));
  INV_X1    g448(.A(new_n630), .ZN(new_n650));
  NOR4_X1   g449(.A1(new_n650), .A2(G36gat), .A3(new_n445), .A4(new_n634), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT46), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n649), .A2(new_n652), .ZN(G1329gat));
  AOI21_X1  g452(.A(new_n522), .B1(new_n446), .B2(new_n448), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n630), .A2(new_n631), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n476), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n656), .B(new_n631), .C1(new_n636), .C2(new_n641), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(KEYINPUT106), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n522), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n657), .A2(KEYINPUT106), .ZN(new_n660));
  OAI211_X1 g459(.A(KEYINPUT47), .B(new_n655), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n655), .B(KEYINPUT104), .Z(new_n662));
  NAND2_X1  g461(.A1(new_n657), .A2(new_n522), .ZN(new_n663));
  AOI21_X1  g462(.A(KEYINPUT47), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI211_X1 g465(.A(KEYINPUT105), .B(KEYINPUT47), .C1(new_n662), .C2(new_n663), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n661), .B1(new_n666), .B2(new_n667), .ZN(G1330gat));
  NAND3_X1  g467(.A1(new_n643), .A2(G50gat), .A3(new_n450), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n650), .A2(new_n426), .A3(new_n634), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n670), .A2(G50gat), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n672));
  NAND3_X1  g471(.A1(new_n669), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(KEYINPUT108), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT108), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n669), .A2(new_n675), .A3(new_n671), .A4(new_n672), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT48), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n669), .A2(new_n671), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n674), .B(new_n676), .C1(new_n677), .C2(new_n678), .ZN(G1331gat));
  INV_X1    g478(.A(new_n611), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n560), .A2(new_n582), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n479), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n434), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g484(.A(new_n445), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(KEYINPUT109), .Z(new_n687));
  NAND2_X1  g486(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n688), .B(new_n689), .Z(G1333gat));
  OAI21_X1  g489(.A(G71gat), .B1(new_n682), .B2(new_n476), .ZN(new_n691));
  INV_X1    g490(.A(G71gat), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n449), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n691), .B1(new_n682), .B2(new_n693), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n694), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g494(.A1(new_n683), .A2(new_n450), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g496(.A1(new_n510), .A2(new_n582), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n630), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT51), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n680), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(new_n536), .A3(new_n434), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT110), .ZN(new_n703));
  INV_X1    g502(.A(new_n698), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(new_n680), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n705), .B1(new_n636), .B2(new_n641), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n703), .B1(new_n706), .B2(new_n292), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(G85gat), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n706), .A2(new_n703), .A3(new_n292), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n702), .B1(new_n708), .B2(new_n709), .ZN(G1336gat));
  NOR2_X1   g509(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  AND4_X1   g511(.A1(new_n479), .A2(new_n558), .A3(new_n698), .A4(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n712), .B1(new_n630), .B2(new_n698), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n617), .A2(new_n537), .A3(new_n611), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n706), .A2(new_n445), .ZN(new_n718));
  OAI22_X1  g517(.A1(new_n717), .A2(KEYINPUT112), .B1(new_n718), .B2(new_n537), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n717), .A2(KEYINPUT112), .ZN(new_n720));
  OAI21_X1  g519(.A(KEYINPUT52), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT52), .ZN(new_n722));
  OAI221_X1 g521(.A(new_n722), .B1(new_n700), .B2(new_n716), .C1(new_n718), .C2(new_n537), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(G1337gat));
  INV_X1    g523(.A(G99gat), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n701), .A2(new_n725), .A3(new_n449), .ZN(new_n726));
  OAI21_X1  g525(.A(G99gat), .B1(new_n706), .B2(new_n476), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(G1338gat));
  INV_X1    g527(.A(G106gat), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n450), .B(new_n705), .C1(new_n636), .C2(new_n641), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n729), .B1(new_n730), .B2(KEYINPUT116), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(KEYINPUT116), .B2(new_n730), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT53), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n611), .A2(new_n729), .A3(new_n450), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT113), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n732), .B(new_n733), .C1(new_n700), .C2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n735), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(new_n713), .B2(new_n714), .ZN(new_n738));
  AOI22_X1  g537(.A1(new_n738), .A2(KEYINPUT114), .B1(new_n730), .B2(G106gat), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT114), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n740), .B(new_n737), .C1(new_n713), .C2(new_n714), .ZN(new_n741));
  AOI211_X1 g540(.A(KEYINPUT115), .B(new_n733), .C1(new_n739), .C2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT115), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n738), .A2(KEYINPUT114), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n730), .A2(G106gat), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n744), .A2(new_n741), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n743), .B1(new_n746), .B2(KEYINPUT53), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n736), .B1(new_n742), .B2(new_n747), .ZN(G1339gat));
  INV_X1    g547(.A(KEYINPUT117), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n568), .A2(new_n569), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n562), .B1(new_n561), .B2(new_n563), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n577), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n752), .A2(new_n581), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n558), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT55), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n584), .B(new_n606), .C1(KEYINPUT10), .C2(new_n587), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n590), .A2(new_n756), .A3(KEYINPUT54), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n594), .B1(new_n608), .B2(KEYINPUT54), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n755), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OR2_X1    g558(.A1(new_n608), .A2(KEYINPUT54), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n590), .A2(new_n756), .A3(KEYINPUT54), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n760), .A2(KEYINPUT55), .A3(new_n594), .A4(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n759), .A2(new_n605), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n749), .B1(new_n754), .B2(new_n763), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n759), .A2(new_n605), .A3(new_n762), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n765), .A2(KEYINPUT117), .A3(new_n753), .A4(new_n558), .ZN(new_n766));
  AOI22_X1  g565(.A1(new_n765), .A2(new_n582), .B1(new_n753), .B2(new_n611), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n764), .B(new_n766), .C1(new_n767), .C2(new_n558), .ZN(new_n768));
  INV_X1    g567(.A(new_n510), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n560), .A2(new_n582), .A3(new_n611), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n617), .A2(new_n292), .A3(new_n427), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n776), .A2(new_n210), .A3(new_n582), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n771), .B1(new_n768), .B2(new_n769), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(new_n450), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n617), .A2(new_n292), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n780), .A2(new_n449), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(G113gat), .B1(new_n783), .B2(new_n583), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n784), .A2(KEYINPUT118), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n784), .A2(KEYINPUT118), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n777), .B1(new_n785), .B2(new_n786), .ZN(G1340gat));
  AOI21_X1  g586(.A(new_n212), .B1(new_n782), .B2(new_n611), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n775), .A2(new_n220), .A3(new_n680), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n788), .A2(new_n789), .ZN(G1341gat));
  OAI21_X1  g589(.A(G127gat), .B1(new_n783), .B2(new_n769), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n769), .A2(G127gat), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n775), .B2(new_n792), .ZN(G1342gat));
  NAND2_X1  g592(.A1(new_n782), .A2(new_n558), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT56), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n775), .A2(G134gat), .A3(new_n559), .ZN(new_n796));
  AOI22_X1  g595(.A1(new_n794), .A2(G134gat), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT119), .ZN(new_n798));
  OR3_X1    g597(.A1(new_n775), .A2(G134gat), .A3(new_n559), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n798), .B1(new_n799), .B2(KEYINPUT56), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n796), .A2(KEYINPUT119), .A3(new_n795), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n797), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT120), .ZN(G1343gat));
  AOI21_X1  g602(.A(new_n426), .B1(new_n770), .B2(new_n772), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n780), .A2(new_n476), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n583), .A2(G141gat), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n804), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT58), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT121), .B1(new_n804), .B2(KEYINPUT57), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n753), .A2(new_n611), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n812), .B1(new_n583), .B2(new_n763), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT122), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n767), .A2(KEYINPUT122), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n815), .A2(new_n816), .A3(new_n559), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n764), .A2(new_n766), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n510), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI211_X1 g618(.A(KEYINPUT57), .B(new_n450), .C1(new_n819), .C2(new_n771), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n821), .B(new_n822), .C1(new_n778), .C2(new_n426), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n811), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n824), .A2(new_n582), .A3(new_n806), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n810), .B1(new_n825), .B2(G141gat), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT124), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI211_X1 g627(.A(KEYINPUT124), .B(new_n810), .C1(new_n825), .C2(G141gat), .ZN(new_n829));
  XOR2_X1   g628(.A(new_n808), .B(KEYINPUT123), .Z(new_n830));
  AOI21_X1  g629(.A(new_n830), .B1(G141gat), .B2(new_n825), .ZN(new_n831));
  OAI22_X1  g630(.A1(new_n828), .A2(new_n829), .B1(new_n809), .B2(new_n831), .ZN(G1344gat));
  INV_X1    g631(.A(new_n804), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n805), .ZN(new_n834));
  INV_X1    g633(.A(G148gat), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n835), .A3(new_n611), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n824), .A2(new_n806), .ZN(new_n837));
  AOI211_X1 g636(.A(KEYINPUT59), .B(new_n835), .C1(new_n837), .C2(new_n611), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n765), .A2(new_n558), .A3(new_n753), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n817), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n772), .B1(new_n841), .B2(new_n510), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT57), .B1(new_n842), .B2(new_n450), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n778), .A2(new_n822), .A3(new_n426), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n611), .B(new_n806), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n839), .B1(new_n845), .B2(G148gat), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n836), .B1(new_n838), .B2(new_n846), .ZN(G1345gat));
  NAND3_X1  g646(.A1(new_n834), .A2(new_n235), .A3(new_n510), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n837), .A2(new_n510), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n848), .B1(new_n849), .B2(new_n235), .ZN(G1346gat));
  AOI21_X1  g649(.A(G162gat), .B1(new_n834), .B2(new_n558), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n559), .A2(new_n236), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n837), .B2(new_n852), .ZN(G1347gat));
  NOR4_X1   g652(.A1(new_n778), .A2(new_n434), .A3(new_n445), .A4(new_n427), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n308), .A3(new_n582), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT125), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n445), .A2(new_n434), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n779), .A2(new_n449), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(G169gat), .B1(new_n858), .B2(new_n583), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n856), .A2(new_n859), .ZN(G1348gat));
  OAI21_X1  g659(.A(G176gat), .B1(new_n858), .B2(new_n680), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n854), .A2(new_n309), .A3(new_n611), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1349gat));
  OAI21_X1  g662(.A(G183gat), .B1(new_n858), .B2(new_n769), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n854), .A2(new_n342), .A3(new_n510), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g665(.A(KEYINPUT126), .B(KEYINPUT60), .ZN(new_n867));
  XOR2_X1   g666(.A(new_n866), .B(new_n867), .Z(G1350gat));
  NAND3_X1  g667(.A1(new_n854), .A2(new_n304), .A3(new_n558), .ZN(new_n869));
  OAI21_X1  g668(.A(G190gat), .B1(new_n858), .B2(new_n559), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n870), .A2(KEYINPUT61), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(KEYINPUT61), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(G1351gat));
  NAND2_X1  g672(.A1(new_n476), .A2(new_n857), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n833), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(G197gat), .B1(new_n875), .B2(new_n582), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n843), .A2(new_n844), .ZN(new_n877));
  INV_X1    g676(.A(new_n874), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n582), .A2(G197gat), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n876), .B1(new_n880), .B2(new_n881), .ZN(G1352gat));
  OAI21_X1  g681(.A(G204gat), .B1(new_n879), .B2(new_n680), .ZN(new_n883));
  NOR4_X1   g682(.A1(new_n833), .A2(G204gat), .A3(new_n680), .A4(new_n874), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(KEYINPUT62), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(G1353gat));
  NAND3_X1  g685(.A1(new_n875), .A2(new_n357), .A3(new_n510), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT127), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n510), .B(new_n878), .C1(new_n843), .C2(new_n844), .ZN(new_n889));
  AND4_X1   g688(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT63), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n357), .B1(KEYINPUT127), .B2(new_n891), .ZN(new_n892));
  AOI22_X1  g691(.A1(new_n889), .A2(new_n892), .B1(new_n888), .B2(KEYINPUT63), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n887), .B1(new_n890), .B2(new_n893), .ZN(G1354gat));
  OAI21_X1  g693(.A(G218gat), .B1(new_n879), .B2(new_n559), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n875), .A2(new_n358), .A3(new_n558), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(G1355gat));
endmodule


