//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  OR2_X1    g003(.A1(KEYINPUT70), .A2(KEYINPUT22), .ZN(new_n205));
  NAND2_X1  g004(.A1(KEYINPUT70), .A2(KEYINPUT22), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n205), .B(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G197gat), .B(G204gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G211gat), .B(G218gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n209), .A2(new_n212), .A3(new_n210), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT2), .ZN(new_n218));
  INV_X1    g017(.A(G155gat), .ZN(new_n219));
  INV_X1    g018(.A(G162gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OR2_X1    g022(.A1(G141gat), .A2(G148gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(G141gat), .A2(G148gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT73), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(new_n218), .ZN(new_n228));
  NAND2_X1  g027(.A1(KEYINPUT73), .A2(KEYINPUT2), .ZN(new_n229));
  AND4_X1   g028(.A1(new_n224), .A2(new_n228), .A3(new_n225), .A4(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT74), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT72), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n232), .A2(new_n219), .A3(new_n220), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT72), .B1(G155gat), .B2(G162gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n222), .A3(new_n234), .ZN(new_n235));
  NOR3_X1   g034(.A1(new_n230), .A2(new_n231), .A3(new_n235), .ZN(new_n236));
  AND3_X1   g035(.A1(new_n233), .A2(new_n222), .A3(new_n234), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n224), .A2(new_n228), .A3(new_n225), .A4(new_n229), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT74), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n226), .B1(new_n236), .B2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n240), .A2(KEYINPUT3), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT71), .B(KEYINPUT29), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n217), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n215), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n212), .B1(new_n209), .B2(new_n210), .ZN(new_n246));
  OAI211_X1 g045(.A(KEYINPUT75), .B(new_n242), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT75), .B1(new_n216), .B2(new_n242), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n240), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G228gat), .A2(G233gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n244), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n252), .ZN(new_n254));
  INV_X1    g053(.A(new_n226), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n231), .B1(new_n230), .B2(new_n235), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n237), .A2(KEYINPUT74), .A3(new_n238), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(new_n248), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n216), .B1(new_n259), .B2(new_n242), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT29), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n216), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n258), .B1(new_n262), .B2(new_n248), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n254), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT31), .B(G50gat), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n253), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n266), .B1(new_n253), .B2(new_n264), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n204), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n264), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(new_n265), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n253), .A2(new_n264), .A3(new_n266), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(new_n203), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(G226gat), .A2(G233gat), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G169gat), .ZN(new_n277));
  INV_X1    g076(.A(G176gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT26), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n281), .B1(G169gat), .B2(G176gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(G183gat), .A2(G190gat), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n283), .B1(new_n279), .B2(new_n280), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n286));
  INV_X1    g085(.A(G183gat), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT66), .B1(new_n287), .B2(KEYINPUT27), .ZN(new_n288));
  AOI21_X1  g087(.A(G190gat), .B1(new_n287), .B2(KEYINPUT27), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT66), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT27), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n291), .A3(G183gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n288), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT67), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT67), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n288), .A2(new_n289), .A3(new_n292), .A4(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n286), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n291), .A2(G183gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n289), .A2(KEYINPUT28), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT69), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n289), .A2(new_n301), .A3(KEYINPUT28), .A4(new_n298), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n285), .B1(new_n297), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n277), .A2(new_n278), .A3(KEYINPUT23), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT23), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(G169gat), .B2(G176gat), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n305), .B(new_n307), .C1(new_n277), .C2(new_n278), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT25), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n311), .B1(G183gat), .B2(G190gat), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n283), .A2(KEYINPUT65), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n283), .A2(KEYINPUT65), .ZN(new_n314));
  NOR3_X1   g113(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT24), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n310), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT24), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n312), .B1(new_n317), .B2(new_n283), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n309), .B1(new_n318), .B2(new_n308), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n276), .B1(new_n321), .B2(new_n242), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n275), .B1(new_n304), .B2(new_n320), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n217), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n321), .A2(new_n276), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT29), .B1(new_n304), .B2(new_n320), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n325), .B(new_n216), .C1(new_n276), .C2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G8gat), .B(G36gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(G64gat), .B(G92gat), .ZN(new_n329));
  XOR2_X1   g128(.A(new_n328), .B(new_n329), .Z(new_n330));
  AND3_X1   g129(.A1(new_n324), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n330), .B1(new_n324), .B2(new_n327), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT30), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n324), .A2(new_n327), .ZN(new_n335));
  INV_X1    g134(.A(new_n330), .ZN(new_n336));
  NOR3_X1   g135(.A1(new_n335), .A2(KEYINPUT30), .A3(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G1gat), .B(G29gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT0), .ZN(new_n340));
  XNOR2_X1  g139(.A(G57gat), .B(G85gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n240), .A2(KEYINPUT3), .ZN(new_n344));
  INV_X1    g143(.A(G134gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G127gat), .ZN(new_n346));
  INV_X1    g145(.A(G127gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(G134gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G113gat), .B(G120gat), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n349), .B1(new_n350), .B2(KEYINPUT1), .ZN(new_n351));
  INV_X1    g150(.A(G120gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(G113gat), .ZN(new_n353));
  INV_X1    g152(.A(G113gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(G120gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G127gat), .B(G134gat), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT1), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n351), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n344), .A2(new_n259), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(G225gat), .A2(G233gat), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n360), .B(new_n226), .C1(new_n236), .C2(new_n239), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n258), .A2(KEYINPUT4), .A3(new_n360), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n362), .A2(new_n363), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT5), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n240), .A2(new_n361), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n364), .ZN(new_n371));
  INV_X1    g170(.A(new_n363), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n366), .A2(new_n367), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n375), .A2(new_n369), .A3(new_n363), .A4(new_n362), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n343), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n370), .A2(new_n363), .A3(new_n364), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT76), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n370), .A2(KEYINPUT76), .A3(new_n363), .A4(new_n364), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n361), .B1(new_n258), .B2(new_n248), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n383), .A2(new_n241), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n366), .A2(new_n367), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n372), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n382), .A2(new_n386), .A3(KEYINPUT39), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n343), .B1(new_n386), .B2(KEYINPUT39), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT40), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n363), .B1(new_n375), .B2(new_n362), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT39), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n342), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT40), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n382), .A2(new_n386), .A3(KEYINPUT39), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n377), .B1(new_n389), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n274), .B1(new_n338), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n374), .A2(new_n376), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n343), .A2(KEYINPUT6), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT6), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n342), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n398), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n374), .A2(new_n400), .A3(new_n376), .A4(new_n342), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n324), .A2(new_n327), .A3(new_n330), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n216), .B1(new_n322), .B2(new_n323), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n325), .B(new_n217), .C1(new_n276), .C2(new_n326), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n406), .A2(KEYINPUT37), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT77), .ZN(new_n409));
  OR2_X1    g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n335), .A2(new_n336), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n336), .A2(KEYINPUT37), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT38), .B1(new_n408), .B2(new_n409), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n410), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  AND2_X1   g214(.A1(new_n335), .A2(KEYINPUT37), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n336), .B1(new_n335), .B2(KEYINPUT37), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT38), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n405), .A2(new_n415), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G227gat), .A2(G233gat), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n420), .B(KEYINPUT64), .Z(new_n421));
  AND3_X1   g220(.A1(new_n304), .A2(new_n360), .A3(new_n320), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n360), .B1(new_n304), .B2(new_n320), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT32), .ZN(new_n425));
  XOR2_X1   g224(.A(G15gat), .B(G43gat), .Z(new_n426));
  XNOR2_X1  g225(.A(G71gat), .B(G99gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n421), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n321), .A2(new_n361), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n304), .A2(new_n360), .A3(new_n320), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n428), .B1(new_n432), .B2(KEYINPUT33), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n430), .A2(new_n429), .A3(new_n431), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT34), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT34), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n430), .A2(new_n436), .A3(new_n429), .A4(new_n431), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n433), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n435), .A2(new_n437), .ZN(new_n439));
  INV_X1    g238(.A(new_n428), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT33), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n440), .B1(new_n424), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n425), .B1(new_n438), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n433), .A2(new_n435), .A3(new_n437), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n422), .A2(new_n423), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n436), .B1(new_n446), .B2(new_n429), .ZN(new_n447));
  INV_X1    g246(.A(new_n437), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n442), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n425), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n445), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n444), .A2(KEYINPUT36), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT36), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n445), .A2(new_n449), .A3(new_n450), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n450), .B1(new_n445), .B2(new_n449), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n397), .A2(new_n419), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n411), .A2(KEYINPUT30), .A3(new_n404), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n458), .A2(new_n459), .B1(new_n403), .B2(new_n402), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n269), .A2(new_n273), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n461), .A2(new_n451), .A3(new_n444), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n402), .A2(new_n403), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n465), .B1(new_n334), .B2(new_n337), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT35), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT78), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n468), .B1(new_n454), .B2(new_n455), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n444), .A2(KEYINPUT78), .A3(new_n451), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n274), .A2(KEYINPUT35), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n469), .A2(new_n470), .A3(new_n460), .A4(new_n471), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n457), .A2(new_n463), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G15gat), .B(G22gat), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT16), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n474), .B1(new_n475), .B2(G1gat), .ZN(new_n476));
  INV_X1    g275(.A(G8gat), .ZN(new_n477));
  OAI221_X1 g276(.A(new_n476), .B1(KEYINPUT80), .B2(new_n477), .C1(G1gat), .C2(new_n474), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(KEYINPUT80), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n478), .B(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(G29gat), .A2(G36gat), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT14), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(G36gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(KEYINPUT79), .B(G29gat), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT15), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n483), .B(KEYINPUT15), .C1(new_n484), .C2(new_n485), .ZN(new_n489));
  XNOR2_X1  g288(.A(G43gat), .B(G50gat), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  OR2_X1    g290(.A1(new_n489), .A2(new_n490), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n480), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n480), .A2(new_n493), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT83), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n480), .A2(new_n493), .A3(KEYINPUT83), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n494), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(G229gat), .A2(G233gat), .ZN(new_n500));
  XOR2_X1   g299(.A(new_n500), .B(KEYINPUT13), .Z(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT81), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT17), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n504), .B1(new_n493), .B2(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT81), .A4(KEYINPUT17), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT17), .B1(new_n491), .B2(new_n492), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n509), .A2(new_n480), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT82), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n508), .A2(KEYINPUT82), .A3(new_n510), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n513), .A2(new_n500), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT18), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n503), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n515), .A2(new_n514), .ZN(new_n519));
  INV_X1    g318(.A(new_n500), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT82), .B1(new_n508), .B2(new_n510), .ZN(new_n521));
  NOR3_X1   g320(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT84), .B1(new_n522), .B2(KEYINPUT18), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT84), .ZN(new_n524));
  NOR3_X1   g323(.A1(new_n516), .A2(new_n524), .A3(new_n517), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n518), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G113gat), .B(G141gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(G197gat), .ZN(new_n528));
  XOR2_X1   g327(.A(KEYINPUT11), .B(G169gat), .Z(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n530), .B(KEYINPUT12), .Z(new_n531));
  NAND2_X1  g330(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n531), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n533), .B(new_n518), .C1(new_n523), .C2(new_n525), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n473), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(G85gat), .A2(G92gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  NAND2_X1  g338(.A1(G99gat), .A2(G106gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT8), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n539), .B(new_n541), .C1(G85gat), .C2(G92gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(G99gat), .B(G106gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT90), .ZN(new_n545));
  NOR2_X1   g344(.A1(G71gat), .A2(G78gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT9), .ZN(new_n547));
  NAND2_X1  g346(.A1(G71gat), .A2(G78gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(G57gat), .B(G64gat), .Z(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(KEYINPUT87), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT85), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n548), .B1(new_n546), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n554), .B1(new_n553), .B2(new_n546), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n550), .A2(KEYINPUT86), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT9), .B1(new_n550), .B2(KEYINPUT86), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n552), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n545), .A2(KEYINPUT10), .A3(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n559), .B(new_n544), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT10), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G230gat), .A2(G233gat), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n566), .B(KEYINPUT93), .Z(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G120gat), .B(G148gat), .Z(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT94), .ZN(new_n571));
  XOR2_X1   g370(.A(G176gat), .B(G204gat), .Z(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n569), .B(new_n574), .C1(new_n568), .C2(new_n562), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n562), .A2(new_n568), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n569), .A2(KEYINPUT95), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT95), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n565), .A2(new_n578), .A3(new_n568), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n576), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n575), .B1(new_n580), .B2(new_n574), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n560), .A2(KEYINPUT21), .ZN(new_n583));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n583), .B(new_n584), .Z(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(G127gat), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n560), .A2(KEYINPUT21), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n587), .A2(new_n480), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n588), .B(KEYINPUT88), .Z(new_n589));
  OR2_X1    g388(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n586), .A2(new_n589), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G183gat), .B(G211gat), .Z(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT89), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(new_n219), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n594), .B(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n592), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n590), .A2(new_n591), .A3(new_n597), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n545), .A2(new_n509), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(new_n508), .ZN(new_n603));
  AND2_X1   g402(.A1(G232gat), .A2(G233gat), .ZN(new_n604));
  AOI22_X1  g403(.A1(new_n545), .A2(new_n493), .B1(KEYINPUT41), .B2(new_n604), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G190gat), .B(G218gat), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n607), .A2(KEYINPUT91), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(KEYINPUT91), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n606), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G134gat), .B(G162gat), .Z(new_n611));
  NOR2_X1   g410(.A1(new_n604), .A2(KEYINPUT41), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT92), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n610), .B(new_n615), .C1(new_n608), .C2(new_n606), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n614), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  AND4_X1   g418(.A1(new_n537), .A2(new_n582), .A3(new_n601), .A4(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n465), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g422(.A1(new_n620), .A2(new_n338), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(G8gat), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n625), .B(KEYINPUT96), .Z(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT16), .B(G8gat), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT42), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT97), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(G1325gat));
  INV_X1    g431(.A(G15gat), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n620), .A2(new_n633), .A3(new_n470), .A4(new_n469), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n456), .A2(new_n452), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n620), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n634), .B1(new_n637), .B2(new_n633), .ZN(G1326gat));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n274), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT98), .ZN(new_n640));
  XOR2_X1   g439(.A(KEYINPUT43), .B(G22gat), .Z(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(G1327gat));
  AND2_X1   g441(.A1(new_n599), .A2(new_n600), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n643), .A2(new_n582), .A3(new_n618), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT99), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n645), .A2(new_n537), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n646), .A2(new_n621), .A3(new_n485), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT45), .ZN(new_n648));
  OAI21_X1  g447(.A(KEYINPUT44), .B1(new_n473), .B2(new_n619), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n467), .A2(new_n472), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n405), .A2(new_n415), .A3(new_n418), .ZN(new_n652));
  INV_X1    g451(.A(new_n377), .ZN(new_n653));
  AND3_X1   g452(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n393), .B1(new_n392), .B2(new_n394), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n458), .A2(new_n459), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n461), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n635), .B1(new_n652), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(KEYINPUT101), .B1(new_n460), .B2(new_n461), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n466), .A2(new_n661), .A3(new_n274), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(KEYINPUT102), .B1(new_n659), .B2(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT101), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n661), .B1(new_n466), .B2(new_n274), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT102), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n457), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n651), .B1(new_n664), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n618), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n649), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n581), .A2(KEYINPUT100), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n581), .A2(KEYINPUT100), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n678), .A2(new_n536), .A3(new_n601), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n673), .A2(new_n674), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n674), .B1(new_n673), .B2(new_n679), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(new_n465), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n648), .B1(new_n684), .B2(new_n485), .ZN(G1328gat));
  NAND3_X1  g484(.A1(new_n646), .A2(new_n484), .A3(new_n338), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(KEYINPUT46), .Z(new_n687));
  OAI21_X1  g486(.A(G36gat), .B1(new_n683), .B2(new_n657), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(G1329gat));
  NAND2_X1  g488(.A1(new_n469), .A2(new_n470), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(G43gat), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n646), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n673), .A2(new_n679), .ZN(new_n694));
  OAI21_X1  g493(.A(G43gat), .B1(new_n694), .B2(new_n635), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n693), .A2(KEYINPUT47), .A3(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT104), .B(KEYINPUT47), .Z(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n650), .B1(new_n659), .B2(new_n462), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n671), .B1(new_n700), .B2(new_n618), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n659), .A2(KEYINPUT102), .A3(new_n663), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n668), .B1(new_n457), .B2(new_n667), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n650), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n672), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n701), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n679), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT103), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n673), .A2(new_n674), .A3(new_n679), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n708), .A2(new_n636), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(G43gat), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n692), .B1(new_n711), .B2(KEYINPUT105), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT105), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n710), .A2(new_n713), .A3(G43gat), .ZN(new_n714));
  AOI211_X1 g513(.A(new_n697), .B(new_n699), .C1(new_n712), .C2(new_n714), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n680), .A2(new_n681), .A3(new_n635), .ZN(new_n716));
  INV_X1    g515(.A(G43gat), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT105), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n718), .A2(new_n714), .A3(new_n693), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT106), .B1(new_n719), .B2(new_n698), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n696), .B1(new_n715), .B2(new_n720), .ZN(G1330gat));
  NOR2_X1   g520(.A1(new_n461), .A2(G50gat), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n646), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G50gat), .B1(new_n694), .B2(new_n461), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n723), .A2(KEYINPUT48), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n682), .A2(new_n274), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n726), .A2(G50gat), .B1(new_n646), .B2(new_n722), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n727), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g527(.A1(new_n643), .A2(new_n535), .A3(new_n618), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n678), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT107), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(new_n670), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n465), .B(KEYINPUT108), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  AND2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n732), .B(new_n338), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n731), .A2(new_n657), .A3(new_n670), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n740), .B2(new_n737), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1333gat));
  INV_X1    g542(.A(G71gat), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n732), .A2(new_n744), .A3(new_n470), .A4(new_n469), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n731), .A2(new_n635), .A3(new_n670), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n746), .B2(new_n744), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n274), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G78gat), .ZN(G1335gat));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n601), .A2(new_n535), .A3(new_n582), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n673), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n751), .B1(new_n753), .B2(new_n465), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G85gat), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n753), .A2(new_n751), .A3(new_n465), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n619), .A2(new_n601), .A3(new_n535), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n704), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n704), .A2(KEYINPUT51), .A3(new_n757), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  OR3_X1    g562(.A1(new_n582), .A2(G85gat), .A3(new_n465), .ZN(new_n764));
  OAI22_X1  g563(.A1(new_n755), .A2(new_n756), .B1(new_n763), .B2(new_n764), .ZN(G1336gat));
  OAI21_X1  g564(.A(KEYINPUT112), .B1(new_n753), .B2(new_n657), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n766), .A2(G92gat), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT112), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n673), .A2(new_n768), .A3(new_n338), .A4(new_n752), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n677), .B1(new_n760), .B2(new_n761), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n657), .A2(G92gat), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(G92gat), .B1(new_n753), .B2(new_n657), .ZN(new_n776));
  AOI22_X1  g575(.A1(KEYINPUT111), .A2(new_n776), .B1(new_n771), .B2(new_n772), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n776), .A2(KEYINPUT111), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI221_X1 g578(.A(KEYINPUT113), .B1(new_n770), .B2(new_n775), .C1(new_n779), .C2(new_n774), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n770), .A2(new_n775), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n774), .B1(new_n777), .B2(new_n778), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n780), .A2(new_n784), .ZN(G1337gat));
  OAI21_X1  g584(.A(G99gat), .B1(new_n753), .B2(new_n635), .ZN(new_n786));
  OR3_X1    g585(.A1(new_n582), .A2(new_n690), .A3(G99gat), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n763), .B2(new_n787), .ZN(G1338gat));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(KEYINPUT53), .ZN(new_n790));
  INV_X1    g589(.A(G106gat), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n771), .A2(new_n791), .A3(new_n274), .ZN(new_n792));
  OAI21_X1  g591(.A(G106gat), .B1(new_n753), .B2(new_n461), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n789), .A2(KEYINPUT53), .ZN(new_n795));
  XOR2_X1   g594(.A(new_n794), .B(new_n795), .Z(G1339gat));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n520), .B1(new_n519), .B2(new_n521), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n499), .A2(new_n502), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n530), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n534), .A2(new_n581), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n577), .A2(new_n804), .A3(new_n579), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n804), .B1(new_n565), .B2(new_n568), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n561), .A2(new_n564), .A3(new_n567), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n574), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n805), .A2(KEYINPUT55), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n575), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n805), .A2(new_n808), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n534), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n522), .A2(KEYINPUT84), .A3(KEYINPUT18), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n524), .B1(new_n516), .B2(new_n517), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n533), .B1(new_n818), .B2(new_n518), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n811), .B(new_n814), .C1(new_n815), .C2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n618), .B1(new_n803), .B2(new_n820), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n534), .A2(new_n801), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n822), .A2(new_n618), .A3(new_n814), .A4(new_n811), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n797), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n810), .B1(new_n532), .B2(new_n534), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n802), .B1(new_n826), .B2(new_n814), .ZN(new_n827));
  OAI211_X1 g626(.A(KEYINPUT115), .B(new_n823), .C1(new_n827), .C2(new_n618), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n825), .A2(new_n828), .A3(new_n643), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n729), .A2(new_n582), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n733), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n464), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n338), .ZN(new_n834));
  AOI21_X1  g633(.A(G113gat), .B1(new_n834), .B2(new_n535), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n274), .B1(new_n829), .B2(new_n830), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n690), .A2(new_n465), .A3(new_n338), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT116), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n836), .A2(new_n841), .A3(new_n837), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n536), .A2(new_n354), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n835), .B1(new_n844), .B2(new_n845), .ZN(G1340gat));
  NAND3_X1  g645(.A1(new_n834), .A2(new_n352), .A3(new_n581), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n839), .A2(new_n678), .A3(new_n842), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n848), .A2(KEYINPUT117), .A3(G120gat), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT117), .B1(new_n848), .B2(G120gat), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n847), .B1(new_n849), .B2(new_n850), .ZN(G1341gat));
  NAND3_X1  g650(.A1(new_n834), .A2(new_n347), .A3(new_n601), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n840), .A2(new_n843), .A3(new_n643), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(new_n347), .ZN(G1342gat));
  NAND2_X1  g653(.A1(new_n618), .A2(new_n657), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n833), .A2(G134gat), .A3(new_n855), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT56), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n840), .A2(new_n843), .A3(new_n619), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n857), .B1(new_n345), .B2(new_n858), .ZN(G1343gat));
  NAND3_X1  g658(.A1(new_n635), .A2(new_n621), .A3(new_n657), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT118), .ZN(new_n861));
  XNOR2_X1  g660(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n829), .A2(new_n830), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n863), .B1(new_n864), .B2(new_n274), .ZN(new_n865));
  XNOR2_X1  g664(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n812), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n535), .A2(new_n811), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n803), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n619), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n601), .B1(new_n870), .B2(new_n823), .ZN(new_n871));
  INV_X1    g670(.A(new_n830), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n274), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n535), .B(new_n861), .C1(new_n865), .C2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(G141gat), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n831), .A2(KEYINPUT121), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n635), .A2(new_n274), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n879), .B1(new_n831), .B2(KEYINPUT121), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n536), .A2(G141gat), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n878), .A2(new_n880), .A3(new_n657), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT58), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT58), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n877), .A2(new_n885), .A3(new_n882), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(G1344gat));
  NAND2_X1  g686(.A1(new_n878), .A2(new_n880), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(new_n338), .ZN(new_n889));
  INV_X1    g688(.A(G148gat), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n889), .A2(new_n890), .A3(new_n581), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n864), .A2(new_n274), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n893), .A2(new_n862), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n873), .A2(new_n874), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n581), .B(new_n861), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n892), .B1(new_n896), .B2(G148gat), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n861), .B1(new_n865), .B2(new_n875), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n898), .A2(new_n582), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n892), .A2(G148gat), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n891), .B1(new_n897), .B2(new_n901), .ZN(G1345gat));
  NAND3_X1  g701(.A1(new_n889), .A2(new_n219), .A3(new_n601), .ZN(new_n903));
  OAI21_X1  g702(.A(G155gat), .B1(new_n898), .B2(new_n643), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1346gat));
  OR3_X1    g704(.A1(new_n888), .A2(G162gat), .A3(new_n855), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT122), .B1(new_n898), .B2(new_n619), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(G162gat), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n898), .A2(KEYINPUT122), .A3(new_n619), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(G1347gat));
  NOR2_X1   g709(.A1(new_n734), .A2(new_n657), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n836), .A2(new_n470), .A3(new_n469), .A4(new_n911), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n912), .A2(new_n277), .A3(new_n536), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n621), .B1(new_n829), .B2(new_n830), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n464), .A2(new_n657), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT123), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(G169gat), .B1(new_n917), .B2(new_n535), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n913), .A2(new_n918), .ZN(G1348gat));
  OAI21_X1  g718(.A(G176gat), .B1(new_n912), .B2(new_n677), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n917), .A2(new_n278), .A3(new_n581), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1349gat));
  NAND2_X1  g721(.A1(new_n287), .A2(KEYINPUT27), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n917), .A2(new_n298), .A3(new_n923), .A4(new_n601), .ZN(new_n924));
  OAI21_X1  g723(.A(G183gat), .B1(new_n912), .B2(new_n643), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g726(.A(G190gat), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n917), .A2(new_n928), .A3(new_n618), .ZN(new_n929));
  OAI21_X1  g728(.A(G190gat), .B1(new_n912), .B2(new_n619), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n930), .A2(KEYINPUT61), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n930), .A2(KEYINPUT61), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(G1351gat));
  NOR2_X1   g732(.A1(new_n879), .A2(new_n657), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n914), .A2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(G197gat), .B1(new_n936), .B2(new_n535), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n894), .A2(new_n895), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n911), .A2(new_n635), .ZN(new_n939));
  XOR2_X1   g738(.A(new_n939), .B(KEYINPUT124), .Z(new_n940));
  AND2_X1   g739(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n535), .A2(G197gat), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n937), .B1(new_n941), .B2(new_n942), .ZN(G1352gat));
  NOR2_X1   g742(.A1(new_n582), .A2(G204gat), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n936), .A2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n946), .A2(KEYINPUT125), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  XOR2_X1   g747(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n949));
  AOI21_X1  g748(.A(new_n948), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n938), .A2(new_n678), .A3(new_n940), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(G204gat), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(G1353gat));
  NAND3_X1  g752(.A1(new_n936), .A2(new_n207), .A3(new_n601), .ZN(new_n954));
  OAI211_X1 g753(.A(new_n601), .B(new_n940), .C1(new_n894), .C2(new_n895), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n955), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n956));
  AOI21_X1  g755(.A(KEYINPUT63), .B1(new_n955), .B2(G211gat), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(G1354gat));
  NAND4_X1  g757(.A1(new_n938), .A2(G218gat), .A3(new_n618), .A4(new_n940), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n208), .B1(new_n935), .B2(new_n619), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(KEYINPUT126), .ZN(new_n961));
  OR2_X1    g760(.A1(new_n960), .A2(KEYINPUT126), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(G1355gat));
endmodule


