//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 0 1 0 0 1 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n584, new_n585, new_n586, new_n588, new_n589,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n819, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888;
  XNOR2_X1  g000(.A(KEYINPUT70), .B(G197gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G204gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT71), .B(G218gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(KEYINPUT22), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G211gat), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n203), .A2(KEYINPUT22), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G218gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT72), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT24), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n214), .B(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OR3_X1    g017(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT65), .B(G190gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n225), .A2(G183gat), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT25), .B1(new_n226), .B2(new_n216), .ZN(new_n227));
  OAI22_X1  g026(.A1(new_n224), .A2(KEYINPUT25), .B1(new_n223), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n228), .B(KEYINPUT66), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT27), .B(G183gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT28), .B1(new_n233), .B2(new_n225), .ZN(new_n234));
  INV_X1    g033(.A(new_n225), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT28), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(new_n236), .A3(new_n230), .ZN(new_n237));
  OR3_X1    g036(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(new_n222), .A3(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n234), .A2(new_n214), .A3(new_n237), .A4(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n229), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G226gat), .A2(G233gat), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n244), .A2(KEYINPUT29), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n241), .A2(new_n228), .ZN(new_n247));
  OAI22_X1  g046(.A1(new_n242), .A2(new_n243), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  OR2_X1    g047(.A1(new_n213), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n242), .A2(new_n245), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n247), .A2(new_n244), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n213), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G8gat), .B(G36gat), .ZN(new_n255));
  INV_X1    g054(.A(G64gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G92gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  OR2_X1    g060(.A1(new_n261), .A2(KEYINPUT30), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(KEYINPUT30), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n249), .A2(new_n253), .A3(new_n259), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT73), .ZN(new_n266));
  OR2_X1    g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n266), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n264), .A2(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(G141gat), .B(G148gat), .Z(new_n271));
  INV_X1    g070(.A(KEYINPUT74), .ZN(new_n272));
  INV_X1    g071(.A(G155gat), .ZN(new_n273));
  INV_X1    g072(.A(G162gat), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT2), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n271), .A2(new_n272), .A3(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G155gat), .B(G162gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT1), .ZN(new_n279));
  XNOR2_X1  g078(.A(G127gat), .B(G134gat), .ZN(new_n280));
  INV_X1    g079(.A(G120gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n281), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(G113gat), .B2(new_n281), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT68), .B1(new_n281), .B2(G113gat), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n279), .B(new_n280), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n280), .ZN(new_n286));
  XNOR2_X1  g085(.A(G113gat), .B(G120gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n286), .B1(KEYINPUT1), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n278), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT4), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT3), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n278), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n293), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(new_n289), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(G225gat), .A2(G233gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(new_n300), .B(KEYINPUT79), .Z(new_n301));
  OR2_X1    g100(.A1(new_n301), .A2(KEYINPUT39), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n278), .B(new_n290), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n301), .B(KEYINPUT39), .C1(new_n299), .C2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT0), .B(G57gat), .ZN(new_n305));
  INV_X1    g104(.A(G85gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G1gat), .B(G29gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n302), .A2(new_n304), .A3(new_n309), .ZN(new_n310));
  OR2_X1    g109(.A1(KEYINPUT80), .A2(KEYINPUT40), .ZN(new_n311));
  OR2_X1    g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT5), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n313), .B1(new_n303), .B2(new_n299), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n298), .B1(new_n278), .B2(new_n290), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n314), .B1(new_n297), .B2(new_n315), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n292), .A2(new_n313), .A3(new_n298), .A4(new_n296), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n309), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n318), .B1(new_n310), .B2(new_n311), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n270), .A2(new_n312), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT29), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n211), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n278), .B1(new_n322), .B2(new_n293), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n295), .A2(new_n321), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n323), .B1(new_n213), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G228gat), .A2(G233gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(G22gat), .ZN(new_n327));
  OR2_X1    g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT77), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n325), .A2(new_n327), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(KEYINPUT76), .B(KEYINPUT31), .ZN(new_n332));
  INV_X1    g131(.A(G50gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n332), .B(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n334), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n328), .A2(new_n329), .A3(new_n336), .A4(new_n330), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G78gat), .B(G106gat), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n339), .B(KEYINPUT78), .Z(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n335), .A2(new_n337), .A3(new_n340), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT37), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n254), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT38), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n213), .A2(new_n248), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n348), .B(KEYINPUT37), .C1(new_n213), .C2(new_n252), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n346), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n254), .B(KEYINPUT37), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n259), .B(new_n350), .C1(new_n351), .C2(new_n347), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n249), .A2(new_n347), .A3(new_n253), .A4(new_n260), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XOR2_X1   g153(.A(KEYINPUT75), .B(KEYINPUT6), .Z(new_n355));
  NOR2_X1   g154(.A1(new_n318), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n316), .A2(new_n317), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n357), .B(new_n309), .Z(new_n358));
  AOI21_X1  g157(.A(new_n356), .B1(new_n358), .B2(new_n355), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n320), .B(new_n344), .C1(new_n354), .C2(new_n359), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n335), .A2(new_n337), .A3(new_n340), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n340), .B1(new_n335), .B2(new_n337), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n262), .A2(new_n263), .B1(new_n267), .B2(new_n268), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n359), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT36), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n242), .B(new_n289), .ZN(new_n368));
  NAND2_X1  g167(.A1(G227gat), .A2(G233gat), .ZN(new_n369));
  XOR2_X1   g168(.A(new_n369), .B(KEYINPUT64), .Z(new_n370));
  OR3_X1    g169(.A1(new_n368), .A2(KEYINPUT34), .A3(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT34), .B1(new_n368), .B2(new_n370), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n368), .A2(new_n370), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT32), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n371), .A2(new_n375), .A3(new_n372), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT33), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT69), .B(G71gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(G99gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(G15gat), .B(G43gat), .ZN(new_n383));
  XOR2_X1   g182(.A(new_n382), .B(new_n383), .Z(new_n384));
  NAND2_X1  g183(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n377), .A2(new_n378), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n386), .B1(new_n377), .B2(new_n378), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n367), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n377), .A2(new_n378), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n385), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n392), .A2(KEYINPUT36), .A3(new_n387), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n360), .A2(new_n366), .A3(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n388), .A2(new_n389), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(new_n361), .B2(new_n362), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT35), .B1(new_n397), .B2(new_n365), .ZN(new_n398));
  INV_X1    g197(.A(new_n365), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT35), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n399), .A2(new_n344), .A3(new_n400), .A4(new_n396), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n395), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G183gat), .B(G211gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(G231gat), .A2(G233gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n404), .B(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(G1gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT16), .ZN(new_n408));
  XNOR2_X1  g207(.A(G15gat), .B(G22gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(KEYINPUT85), .ZN(new_n410));
  MUX2_X1   g209(.A(new_n408), .B(new_n407), .S(new_n410), .Z(new_n411));
  INV_X1    g210(.A(G8gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT21), .ZN(new_n414));
  AND2_X1   g213(.A1(G71gat), .A2(G78gat), .ZN(new_n415));
  NOR2_X1   g214(.A1(G71gat), .A2(G78gat), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G57gat), .B(G64gat), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(G57gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(G64gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n256), .A2(G57gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G71gat), .B(G78gat), .ZN(new_n425));
  INV_X1    g224(.A(new_n419), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n420), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n413), .B1(new_n414), .B2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(KEYINPUT86), .ZN(new_n430));
  XOR2_X1   g229(.A(G127gat), .B(G155gat), .Z(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n430), .A2(new_n431), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n406), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n434), .ZN(new_n436));
  INV_X1    g235(.A(new_n406), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(new_n437), .A3(new_n432), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n428), .A2(new_n414), .ZN(new_n439));
  XOR2_X1   g238(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(new_n440), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n435), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n441), .B1(new_n435), .B2(new_n438), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT14), .ZN(new_n446));
  NOR2_X1   g245(.A1(G29gat), .A2(G36gat), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT83), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT83), .B1(G29gat), .B2(G36gat), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n449), .B(new_n451), .ZN(new_n452));
  XOR2_X1   g251(.A(G43gat), .B(G50gat), .Z(new_n453));
  INV_X1    g252(.A(KEYINPUT15), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(G29gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(KEYINPUT84), .B(G36gat), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n452), .B(new_n455), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  OR2_X1    g257(.A1(new_n453), .A2(new_n454), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n458), .B(new_n459), .ZN(new_n460));
  OR2_X1    g259(.A1(new_n460), .A2(KEYINPUT17), .ZN(new_n461));
  XOR2_X1   g260(.A(G99gat), .B(G106gat), .Z(new_n462));
  NAND2_X1  g261(.A1(G85gat), .A2(G92gat), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT7), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT87), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT87), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT7), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n464), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n469), .B1(new_n464), .B2(new_n466), .ZN(new_n470));
  NAND2_X1  g269(.A1(G99gat), .A2(G106gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT8), .ZN(new_n472));
  XNOR2_X1  g271(.A(KEYINPUT88), .B(G92gat), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n472), .B1(new_n473), .B2(G85gat), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n462), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n463), .A2(KEYINPUT87), .A3(new_n465), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT87), .B(KEYINPUT7), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n476), .B1(new_n464), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n258), .A2(KEYINPUT88), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT88), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(G92gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n482), .A2(new_n306), .B1(KEYINPUT8), .B2(new_n471), .ZN(new_n483));
  INV_X1    g282(.A(new_n462), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n478), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n475), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n460), .A2(KEYINPUT17), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n461), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AND2_X1   g287(.A1(G232gat), .A2(G233gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT41), .ZN(new_n490));
  XOR2_X1   g289(.A(G190gat), .B(G218gat), .Z(new_n491));
  NOR2_X1   g290(.A1(new_n491), .A2(KEYINPUT89), .ZN(new_n492));
  INV_X1    g291(.A(new_n460), .ZN(new_n493));
  INV_X1    g292(.A(new_n486), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n488), .A2(new_n490), .A3(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(G134gat), .B(G162gat), .Z(new_n497));
  OR2_X1    g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n491), .A2(KEYINPUT89), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n489), .A2(KEYINPUT41), .ZN(new_n500));
  XOR2_X1   g299(.A(new_n499), .B(new_n500), .Z(new_n501));
  NAND2_X1  g300(.A1(new_n496), .A2(new_n497), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n498), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n501), .B1(new_n498), .B2(new_n502), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n411), .B(G8gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n493), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n413), .A2(new_n460), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(G229gat), .A2(G233gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(KEYINPUT13), .ZN(new_n512));
  OR2_X1    g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n461), .A2(new_n413), .A3(new_n487), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n514), .A2(new_n508), .A3(new_n511), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT18), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n514), .A2(KEYINPUT18), .A3(new_n508), .A4(new_n511), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n513), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(G113gat), .B(G141gat), .Z(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(KEYINPUT82), .ZN(new_n521));
  XOR2_X1   g320(.A(G169gat), .B(G197gat), .Z(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  XOR2_X1   g322(.A(KEYINPUT81), .B(KEYINPUT11), .Z(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT12), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n519), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n513), .A2(new_n517), .A3(new_n518), .A4(new_n526), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NOR3_X1   g330(.A1(new_n470), .A2(new_n474), .A3(new_n462), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n484), .B1(new_n478), .B2(new_n483), .ZN(new_n533));
  OAI22_X1  g332(.A1(new_n532), .A2(new_n533), .B1(KEYINPUT90), .B2(new_n428), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT90), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n420), .A2(new_n427), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n535), .B1(new_n420), .B2(new_n427), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n485), .B(new_n475), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT10), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n534), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT91), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n534), .A2(new_n538), .A3(KEYINPUT91), .A4(new_n539), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n486), .A2(new_n539), .A3(new_n428), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(G230gat), .A2(G233gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n538), .ZN(new_n550));
  INV_X1    g349(.A(new_n548), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n549), .A2(KEYINPUT92), .A3(new_n552), .ZN(new_n553));
  OR2_X1    g352(.A1(new_n552), .A2(KEYINPUT92), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(G120gat), .B(G148gat), .Z(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(G176gat), .ZN(new_n557));
  INV_X1    g356(.A(G204gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n559), .B(KEYINPUT93), .Z(new_n560));
  NAND2_X1  g359(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT94), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n553), .A2(new_n554), .ZN(new_n563));
  INV_X1    g362(.A(new_n559), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT94), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n555), .A2(new_n566), .A3(new_n560), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n562), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  NOR4_X1   g367(.A1(new_n445), .A2(new_n506), .A3(new_n531), .A4(new_n568), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n403), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n359), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g372(.A1(new_n570), .A2(new_n270), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n574), .B(KEYINPUT96), .Z(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(G8gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(KEYINPUT16), .B(G8gat), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT42), .ZN(new_n579));
  NAND2_X1  g378(.A1(KEYINPUT95), .A2(KEYINPUT42), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n580), .B1(new_n575), .B2(new_n577), .ZN(new_n581));
  NOR2_X1   g380(.A1(KEYINPUT95), .A2(KEYINPUT42), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n576), .B(new_n579), .C1(new_n581), .C2(new_n582), .ZN(G1325gat));
  AOI21_X1  g382(.A(G15gat), .B1(new_n570), .B2(new_n396), .ZN(new_n584));
  INV_X1    g383(.A(new_n394), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n570), .A2(G15gat), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(G1326gat));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n363), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT43), .B(G22gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(G1327gat));
  NOR2_X1   g389(.A1(new_n505), .A2(KEYINPUT44), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n395), .A2(new_n402), .A3(KEYINPUT97), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT97), .B1(new_n395), .B2(new_n402), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n591), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n505), .B1(new_n395), .B2(new_n402), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT44), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NOR3_X1   g399(.A1(new_n444), .A2(new_n531), .A3(new_n568), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(G29gat), .B1(new_n602), .B2(new_n359), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n596), .A2(new_n601), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n604), .A2(new_n456), .A3(new_n571), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT45), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(G1328gat));
  NAND3_X1  g406(.A1(new_n604), .A2(new_n270), .A3(new_n457), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n608), .B(KEYINPUT46), .Z(new_n609));
  NOR2_X1   g408(.A1(new_n602), .A2(new_n364), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n609), .B1(new_n457), .B2(new_n610), .ZN(G1329gat));
  NAND3_X1  g410(.A1(new_n600), .A2(G43gat), .A3(new_n601), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n604), .A2(new_n396), .ZN(new_n613));
  OAI22_X1  g412(.A1(new_n612), .A2(new_n394), .B1(G43gat), .B2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g414(.A1(new_n363), .A2(G50gat), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n604), .A2(new_n363), .ZN(new_n617));
  OAI22_X1  g416(.A1(new_n602), .A2(new_n616), .B1(G50gat), .B2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g418(.A(KEYINPUT97), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n403), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(new_n592), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n444), .A2(new_n505), .A3(new_n531), .ZN(new_n623));
  INV_X1    g422(.A(new_n568), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n625), .B(KEYINPUT98), .Z(new_n626));
  AND2_X1   g425(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n571), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT99), .B(G57gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(G1332gat));
  NAND2_X1  g429(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n627), .A2(new_n270), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(KEYINPUT100), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT100), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n627), .A2(new_n634), .A3(new_n270), .A4(new_n631), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n636), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n637));
  NOR2_X1   g436(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n633), .A2(new_n638), .A3(new_n635), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(G1333gat));
  NAND3_X1  g439(.A1(new_n627), .A2(G71gat), .A3(new_n585), .ZN(new_n641));
  INV_X1    g440(.A(G71gat), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n622), .A2(new_n626), .ZN(new_n643));
  INV_X1    g442(.A(new_n396), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g446(.A1(new_n627), .A2(new_n363), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g448(.A1(new_n445), .A2(new_n531), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n591), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n652), .B1(new_n621), .B2(new_n592), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n568), .B(new_n651), .C1(new_n653), .C2(new_n598), .ZN(new_n654));
  OAI21_X1  g453(.A(G85gat), .B1(new_n654), .B2(new_n359), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n596), .A2(new_n651), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT101), .B(KEYINPUT51), .Z(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT51), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n656), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n571), .A2(new_n306), .A3(new_n568), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT102), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n655), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT103), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n655), .B(KEYINPUT103), .C1(new_n663), .C2(new_n665), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(G1336gat));
  OAI21_X1  g469(.A(new_n661), .B1(new_n657), .B2(KEYINPUT104), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n656), .A2(new_n672), .A3(KEYINPUT51), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n364), .A2(new_n624), .A3(G92gat), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n600), .A2(new_n270), .A3(new_n568), .A4(new_n651), .ZN(new_n676));
  AOI22_X1  g475(.A1(new_n674), .A2(new_n675), .B1(new_n676), .B2(new_n473), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT52), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n676), .A2(new_n473), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n675), .B1(new_n659), .B2(new_n662), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n678), .ZN(new_n681));
  OAI22_X1  g480(.A1(new_n677), .A2(new_n678), .B1(new_n679), .B2(new_n681), .ZN(G1337gat));
  OR4_X1    g481(.A1(G99gat), .A2(new_n663), .A3(new_n644), .A4(new_n624), .ZN(new_n683));
  OAI21_X1  g482(.A(G99gat), .B1(new_n654), .B2(new_n394), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(G1338gat));
  INV_X1    g484(.A(G106gat), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n686), .A2(KEYINPUT105), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(KEYINPUT105), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n687), .B(new_n688), .C1(new_n654), .C2(new_n344), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT53), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n344), .A2(G106gat), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n568), .B(new_n691), .C1(new_n659), .C2(new_n662), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n671), .A2(new_n568), .A3(new_n673), .A4(new_n691), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n693), .B1(new_n695), .B2(new_n690), .ZN(G1339gat));
  AOI21_X1  g495(.A(new_n511), .B1(new_n514), .B2(new_n508), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n508), .A2(new_n509), .A3(new_n512), .ZN(new_n698));
  OAI211_X1 g497(.A(KEYINPUT109), .B(new_n525), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n525), .B1(new_n697), .B2(new_n698), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT109), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n529), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n568), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n544), .A2(new_n551), .A3(new_n546), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n549), .A2(KEYINPUT106), .A3(KEYINPUT54), .A4(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n551), .B1(new_n544), .B2(new_n546), .ZN(new_n707));
  AOI211_X1 g506(.A(new_n548), .B(new_n545), .C1(new_n542), .C2(new_n543), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT54), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n711), .B1(new_n707), .B2(new_n709), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n706), .B(new_n559), .C1(new_n710), .C2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT55), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n565), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n713), .A2(new_n714), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT108), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n713), .A2(new_n720), .A3(new_n714), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n565), .B(KEYINPUT107), .C1(new_n713), .C2(new_n714), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n717), .A2(new_n719), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n704), .B1(new_n723), .B2(new_n531), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI211_X1 g525(.A(KEYINPUT110), .B(new_n704), .C1(new_n723), .C2(new_n531), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n726), .A2(new_n505), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n506), .A2(new_n703), .ZN(new_n729));
  OR2_X1    g528(.A1(new_n729), .A2(new_n723), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n444), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n623), .A2(new_n568), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n733), .A2(new_n571), .A3(new_n364), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n397), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n530), .ZN(new_n736));
  XNOR2_X1  g535(.A(KEYINPUT111), .B(G113gat), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1340gat));
  NAND2_X1  g537(.A1(new_n735), .A2(new_n568), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g539(.A1(new_n735), .A2(new_n444), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(G127gat), .ZN(G1342gat));
  NOR3_X1   g541(.A1(new_n734), .A2(new_n397), .A3(new_n505), .ZN(new_n743));
  INV_X1    g542(.A(G134gat), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n745), .A2(KEYINPUT56), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(KEYINPUT56), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n746), .B(new_n747), .C1(new_n744), .C2(new_n743), .ZN(G1343gat));
  OAI21_X1  g547(.A(new_n571), .B1(new_n731), .B2(new_n732), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT114), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI211_X1 g550(.A(KEYINPUT114), .B(new_n571), .C1(new_n731), .C2(new_n732), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n270), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(G141gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n394), .A2(new_n363), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT115), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n753), .A2(new_n754), .A3(new_n530), .A4(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT58), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT57), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n759), .B(new_n363), .C1(new_n731), .C2(new_n732), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n388), .A2(new_n389), .A3(new_n367), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT36), .B1(new_n392), .B2(new_n387), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n571), .B(new_n364), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT112), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n394), .A2(new_n765), .A3(new_n571), .A4(new_n364), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n530), .A2(new_n718), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n704), .B1(new_n715), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n505), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n444), .B1(new_n770), .B2(new_n730), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n363), .B1(new_n771), .B2(new_n732), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n767), .B1(new_n772), .B2(KEYINPUT57), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n760), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(G141gat), .B1(new_n774), .B2(new_n531), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n757), .A2(new_n758), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT116), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT113), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n760), .A2(new_n773), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n778), .B1(new_n760), .B2(new_n773), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n530), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G141gat), .ZN(new_n782));
  AOI211_X1 g581(.A(new_n777), .B(new_n758), .C1(new_n782), .C2(new_n757), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n774), .A2(KEYINPUT113), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n760), .A2(new_n773), .A3(new_n778), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n531), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n757), .B1(new_n786), .B2(new_n754), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT116), .B1(new_n787), .B2(KEYINPUT58), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n776), .B1(new_n783), .B2(new_n788), .ZN(G1344gat));
  OAI21_X1  g588(.A(new_n568), .B1(new_n779), .B2(new_n780), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT59), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n790), .A2(new_n791), .A3(G148gat), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT117), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n790), .A2(KEYINPUT117), .A3(new_n791), .A4(G148gat), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n733), .A2(new_n363), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT57), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n732), .B(KEYINPUT118), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n759), .B(new_n363), .C1(new_n799), .C2(new_n771), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n767), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n568), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n791), .B1(new_n803), .B2(G148gat), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n753), .A2(new_n756), .ZN(new_n805));
  OR2_X1    g604(.A1(new_n624), .A2(G148gat), .ZN(new_n806));
  OAI22_X1  g605(.A1(new_n796), .A2(new_n804), .B1(new_n805), .B2(new_n806), .ZN(G1345gat));
  OAI21_X1  g606(.A(new_n444), .B1(new_n779), .B2(new_n780), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n805), .A2(new_n445), .ZN(new_n809));
  MUX2_X1   g608(.A(new_n808), .B(new_n809), .S(new_n273), .Z(G1346gat));
  NAND4_X1  g609(.A1(new_n753), .A2(new_n274), .A3(new_n506), .A4(new_n756), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n505), .B1(new_n784), .B2(new_n785), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n811), .B1(new_n812), .B2(new_n274), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT119), .ZN(G1347gat));
  INV_X1    g613(.A(new_n397), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n364), .A2(new_n571), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n815), .B(new_n816), .C1(new_n731), .C2(new_n732), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n530), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n568), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g621(.A1(new_n818), .A2(new_n232), .A3(new_n444), .ZN(new_n823));
  OAI21_X1  g622(.A(G183gat), .B1(new_n817), .B2(new_n445), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n825), .A2(KEYINPUT120), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(KEYINPUT120), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT60), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n826), .A2(KEYINPUT60), .A3(new_n827), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(G1350gat));
  OAI21_X1  g631(.A(G190gat), .B1(new_n817), .B2(new_n505), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT121), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT121), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n835), .B(G190gat), .C1(new_n817), .C2(new_n505), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT122), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT61), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n818), .A2(new_n235), .A3(new_n506), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n838), .A2(new_n839), .ZN(new_n842));
  NAND2_X1  g641(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n834), .A2(new_n842), .A3(new_n843), .A4(new_n836), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n840), .A2(new_n841), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT123), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT123), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n840), .A2(new_n847), .A3(new_n841), .A4(new_n844), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(G1351gat));
  INV_X1    g648(.A(G197gat), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n798), .A2(new_n800), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n394), .A2(new_n816), .ZN(new_n852));
  XOR2_X1   g651(.A(new_n852), .B(KEYINPUT124), .Z(new_n853));
  NOR2_X1   g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n850), .B1(new_n854), .B2(new_n530), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n733), .A2(new_n363), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n852), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n857), .A2(G197gat), .A3(new_n531), .ZN(new_n858));
  OAI21_X1  g657(.A(KEYINPUT125), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n858), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT125), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n851), .A2(new_n531), .A3(new_n853), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n860), .B(new_n861), .C1(new_n862), .C2(new_n850), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n859), .A2(new_n863), .ZN(G1352gat));
  INV_X1    g663(.A(KEYINPUT126), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n851), .A2(new_n624), .ZN(new_n866));
  INV_X1    g665(.A(new_n853), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n558), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n624), .A2(G204gat), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT62), .B1(new_n857), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT62), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n856), .A2(new_n872), .A3(new_n852), .A4(new_n869), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n865), .B1(new_n868), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n801), .A2(new_n568), .A3(new_n867), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(G204gat), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n871), .A2(new_n873), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n877), .A2(new_n878), .A3(KEYINPUT126), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n875), .A2(new_n879), .ZN(G1353gat));
  INV_X1    g679(.A(new_n857), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n207), .A3(new_n444), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n801), .A2(new_n444), .A3(new_n867), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n883), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT63), .B1(new_n883), .B2(G211gat), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(G1354gat));
  AOI21_X1  g685(.A(G218gat), .B1(new_n881), .B2(new_n506), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n506), .A2(new_n204), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n854), .B2(new_n888), .ZN(G1355gat));
endmodule


