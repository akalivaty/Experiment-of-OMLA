//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT87), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(G110), .B(G140), .ZN(new_n191));
  INV_X1    g005(.A(G227), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G953), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n191), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n196));
  INV_X1    g010(.A(G104), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(G107), .ZN(new_n198));
  INV_X1    g012(.A(G107), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(KEYINPUT3), .A3(G104), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT88), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n202), .B1(new_n199), .B2(G104), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n197), .A2(KEYINPUT88), .A3(G107), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n201), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G101), .ZN(new_n206));
  INV_X1    g020(.A(G101), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n201), .A2(new_n207), .A3(new_n203), .A4(new_n204), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(KEYINPUT4), .A3(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT0), .B(G128), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n211), .A2(G143), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G143), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT64), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n210), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n216), .A2(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n212), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT0), .ZN(new_n222));
  INV_X1    g036(.A(G128), .ZN(new_n223));
  NOR3_X1   g037(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT4), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n205), .A2(new_n226), .A3(G101), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n209), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT1), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n229), .B1(G143), .B2(new_n211), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT89), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n223), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT1), .B1(new_n216), .B2(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT89), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n232), .A2(new_n234), .B1(new_n212), .B2(new_n220), .ZN(new_n235));
  NOR3_X1   g049(.A1(new_n221), .A2(KEYINPUT1), .A3(new_n223), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n199), .A2(G104), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n197), .A2(G107), .ZN(new_n239));
  OAI21_X1  g053(.A(G101), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n208), .A2(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n228), .B1(new_n242), .B2(KEYINPUT10), .ZN(new_n243));
  INV_X1    g057(.A(new_n236), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n245));
  AOI221_X4 g059(.A(new_n245), .B1(G128), .B2(new_n233), .C1(new_n215), .C2(new_n218), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n214), .B1(new_n216), .B2(G146), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n218), .B1(new_n217), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n233), .A2(G128), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT69), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n244), .B1(new_n246), .B2(new_n250), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n208), .A2(new_n240), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n251), .A2(KEYINPUT10), .A3(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n243), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT66), .B(G134), .ZN(new_n255));
  AOI21_X1  g069(.A(KEYINPUT67), .B1(new_n255), .B2(G137), .ZN(new_n256));
  INV_X1    g070(.A(G134), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT66), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT66), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G134), .ZN(new_n260));
  AND4_X1   g074(.A1(KEYINPUT67), .A2(new_n258), .A3(new_n260), .A4(G137), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G137), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(KEYINPUT11), .A3(G134), .ZN(new_n264));
  AOI21_X1  g078(.A(G137), .B1(new_n258), .B2(new_n260), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT65), .B(KEYINPUT11), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(G131), .B1(new_n262), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT68), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT67), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n258), .A2(new_n260), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n270), .B1(new_n271), .B2(new_n263), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n255), .A2(KEYINPUT67), .A3(G137), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n264), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n271), .A2(new_n263), .ZN(new_n276));
  INV_X1    g090(.A(new_n266), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G131), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n274), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n268), .A2(new_n269), .A3(new_n280), .ZN(new_n281));
  OAI211_X1 g095(.A(KEYINPUT68), .B(G131), .C1(new_n262), .C2(new_n267), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n254), .A2(new_n283), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n281), .A2(new_n282), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n285), .B1(new_n243), .B2(new_n253), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n195), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n244), .B(new_n241), .C1(new_n246), .C2(new_n250), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n252), .B1(new_n236), .B2(new_n235), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n285), .A2(KEYINPUT90), .A3(KEYINPUT12), .A4(new_n290), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n290), .A2(KEYINPUT12), .A3(new_n282), .A4(new_n281), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT90), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT12), .ZN(new_n295));
  INV_X1    g109(.A(new_n290), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n295), .B1(new_n296), .B2(new_n283), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n291), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n194), .B1(new_n254), .B2(new_n283), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT91), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n287), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n298), .A2(KEYINPUT91), .A3(new_n299), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G469), .ZN(new_n305));
  INV_X1    g119(.A(G902), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n195), .B1(new_n298), .B2(new_n284), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n299), .A2(new_n286), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G469), .B1(new_n310), .B2(G902), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n190), .B1(new_n307), .B2(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(G128), .B(G143), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n271), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n255), .A2(new_n313), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G116), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT100), .B1(new_n318), .B2(G122), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT100), .ZN(new_n320));
  INV_X1    g134(.A(G122), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G116), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n318), .A2(G122), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n317), .B1(G107), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n324), .B(KEYINPUT14), .ZN(new_n327));
  INV_X1    g141(.A(new_n323), .ZN(new_n328));
  OAI21_X1  g142(.A(G107), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT102), .ZN(new_n330));
  OR2_X1    g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n330), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n326), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  XOR2_X1   g148(.A(KEYINPUT101), .B(KEYINPUT13), .Z(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(G128), .A3(new_n216), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n336), .B(G134), .C1(new_n335), .C2(new_n314), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n316), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n325), .B(new_n199), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G953), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G217), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n188), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n334), .A2(new_n341), .A3(new_n344), .ZN(new_n345));
  OAI22_X1  g159(.A1(new_n333), .A2(new_n340), .B1(new_n188), .B2(new_n343), .ZN(new_n346));
  AOI21_X1  g160(.A(G902), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G478), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n348), .A2(KEYINPUT15), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  AOI211_X1 g165(.A(G902), .B(new_n349), .C1(new_n345), .C2(new_n346), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G237), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(new_n342), .A3(G214), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n216), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n354), .A2(new_n342), .A3(G143), .A4(G214), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n279), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT96), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n279), .A3(new_n357), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT17), .ZN(new_n362));
  OR2_X1    g176(.A1(new_n360), .A2(new_n359), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT98), .ZN(new_n365));
  INV_X1    g179(.A(G125), .ZN(new_n366));
  NOR3_X1   g180(.A1(new_n366), .A2(KEYINPUT16), .A3(G140), .ZN(new_n367));
  XNOR2_X1  g181(.A(G125), .B(G140), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n367), .B1(new_n368), .B2(KEYINPUT16), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n369), .B(new_n211), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT97), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n370), .A2(new_n371), .B1(KEYINPUT17), .B2(new_n358), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT98), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n361), .A2(new_n363), .A3(new_n373), .A4(new_n362), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n369), .B(G146), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT97), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n365), .A2(new_n372), .A3(new_n374), .A4(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(G113), .B(G122), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n378), .B(new_n197), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT95), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n358), .A2(new_n380), .A3(KEYINPUT18), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n368), .B(new_n211), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(KEYINPUT18), .A3(G131), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n356), .A2(new_n357), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n381), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n377), .A2(new_n379), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n379), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n369), .A2(G146), .ZN(new_n388));
  XOR2_X1   g202(.A(new_n368), .B(KEYINPUT19), .Z(new_n389));
  OAI21_X1  g203(.A(new_n388), .B1(new_n389), .B2(G146), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n390), .B1(new_n363), .B2(new_n361), .ZN(new_n391));
  INV_X1    g205(.A(new_n385), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n387), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n386), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT20), .ZN(new_n395));
  NOR2_X1   g209(.A1(G475), .A2(G902), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(KEYINPUT99), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n394), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  XOR2_X1   g213(.A(KEYINPUT94), .B(KEYINPUT20), .Z(new_n400));
  AOI21_X1  g214(.A(new_n397), .B1(new_n386), .B2(new_n393), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n386), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n379), .B1(new_n377), .B2(new_n385), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n306), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G475), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n353), .A2(new_n402), .A3(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(G110), .B(G122), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT71), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT2), .ZN(new_n410));
  INV_X1    g224(.A(G113), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(KEYINPUT71), .A2(KEYINPUT2), .A3(G113), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n412), .A2(new_n413), .B1(new_n410), .B2(new_n411), .ZN(new_n414));
  INV_X1    g228(.A(G119), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G116), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n318), .A2(G119), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT72), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n414), .B(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n209), .A2(new_n420), .A3(new_n227), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n414), .A2(new_n416), .A3(new_n417), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n416), .A2(new_n417), .A3(KEYINPUT5), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n423), .B(G113), .C1(KEYINPUT5), .C2(new_n416), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n252), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n408), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT6), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT6), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n421), .A2(new_n408), .A3(new_n425), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT92), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT92), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n421), .A2(new_n425), .A3(new_n431), .A4(new_n408), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n428), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n427), .B1(new_n433), .B2(new_n426), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n251), .A2(new_n366), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n219), .A2(new_n224), .A3(new_n366), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n342), .A2(G224), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n438), .B(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n434), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G210), .B1(G237), .B2(G902), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n435), .A2(new_n437), .B1(KEYINPUT7), .B2(new_n439), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n439), .A2(KEYINPUT7), .ZN(new_n444));
  AOI211_X1 g258(.A(new_n436), .B(new_n444), .C1(new_n251), .C2(new_n366), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n422), .A2(new_n424), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n252), .B(new_n446), .ZN(new_n447));
  XOR2_X1   g261(.A(new_n408), .B(KEYINPUT8), .Z(new_n448));
  OAI22_X1  g262(.A1(new_n443), .A2(new_n445), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n430), .A2(new_n432), .ZN(new_n451));
  AOI21_X1  g265(.A(G902), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n441), .A2(new_n442), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n451), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n306), .B1(new_n454), .B2(new_n449), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(new_n434), .B2(new_n440), .ZN(new_n456));
  XOR2_X1   g270(.A(new_n442), .B(KEYINPUT93), .Z(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n453), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G952), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(G953), .ZN(new_n461));
  INV_X1    g275(.A(G234), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n461), .B1(new_n462), .B2(new_n354), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT21), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n465), .A2(G898), .ZN(new_n466));
  OAI21_X1  g280(.A(G953), .B1(new_n465), .B2(G898), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n306), .B1(G234), .B2(G237), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(G214), .B1(G237), .B2(G902), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n407), .A2(new_n459), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n312), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n281), .A2(new_n282), .A3(new_n225), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT70), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n263), .A2(G134), .ZN(new_n478));
  OAI21_X1  g292(.A(G131), .B1(new_n265), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n280), .A2(new_n479), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n214), .A2(new_n216), .A3(G146), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n481), .B1(new_n212), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n249), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n245), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n248), .A2(KEYINPUT69), .A3(new_n249), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n236), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n477), .B1(new_n480), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n251), .A2(KEYINPUT70), .A3(new_n280), .A4(new_n479), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n476), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n420), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n420), .B(KEYINPUT75), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT73), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n480), .B2(new_n487), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n251), .A2(KEYINPUT73), .A3(new_n280), .A4(new_n479), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n476), .A2(new_n492), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT77), .B1(new_n497), .B2(KEYINPUT28), .ZN(new_n498));
  XOR2_X1   g312(.A(new_n420), .B(KEYINPUT75), .Z(new_n499));
  NOR2_X1   g313(.A1(new_n480), .A2(new_n487), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n476), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT28), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n476), .A2(new_n494), .A3(new_n495), .ZN(new_n505));
  AOI22_X1  g319(.A1(new_n505), .A2(new_n492), .B1(new_n490), .B2(new_n420), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n504), .B1(new_n506), .B2(new_n503), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n498), .B1(new_n507), .B2(KEYINPUT77), .ZN(new_n508));
  XOR2_X1   g322(.A(KEYINPUT26), .B(G101), .Z(new_n509));
  NAND3_X1  g323(.A1(new_n354), .A2(new_n342), .A3(G210), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n509), .B(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT76), .B(KEYINPUT27), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n511), .B(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(KEYINPUT78), .B1(new_n508), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n503), .B1(new_n491), .B2(new_n496), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT28), .B1(new_n501), .B2(new_n476), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT77), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT77), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n518), .B1(new_n506), .B2(new_n503), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT78), .ZN(new_n521));
  INV_X1    g335(.A(new_n513), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT30), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n490), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n476), .A2(new_n494), .A3(KEYINPUT30), .A4(new_n495), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n420), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT74), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n525), .A2(KEYINPUT74), .A3(new_n420), .A4(new_n526), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n529), .A2(new_n513), .A3(new_n496), .A4(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT31), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n530), .A2(new_n496), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n534), .A2(KEYINPUT31), .A3(new_n513), .A4(new_n529), .ZN(new_n535));
  AOI22_X1  g349(.A1(new_n514), .A2(new_n523), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(G472), .A2(G902), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(KEYINPUT32), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n533), .A2(new_n535), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n521), .B1(new_n520), .B2(new_n522), .ZN(new_n541));
  AOI211_X1 g355(.A(KEYINPUT78), .B(new_n513), .C1(new_n517), .C2(new_n519), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT32), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n544), .A3(new_n537), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n476), .A2(new_n494), .A3(new_n495), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n499), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n547), .A2(KEYINPUT79), .A3(new_n496), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT79), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n546), .A2(new_n549), .A3(new_n499), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n548), .A2(KEYINPUT28), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT29), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n522), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n551), .A2(new_n504), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n306), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n529), .A2(new_n496), .A3(new_n530), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT29), .B1(new_n556), .B2(new_n522), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n517), .A2(new_n513), .A3(new_n519), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n555), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(G472), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT80), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n527), .A2(new_n528), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n530), .A2(new_n496), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n522), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n564), .A2(new_n558), .A3(new_n552), .ZN(new_n565));
  INV_X1    g379(.A(new_n555), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT80), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(new_n568), .A3(G472), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n539), .A2(new_n545), .B1(new_n561), .B2(new_n569), .ZN(new_n570));
  XOR2_X1   g384(.A(KEYINPUT24), .B(G110), .Z(new_n571));
  XNOR2_X1  g385(.A(G119), .B(G128), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT82), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(KEYINPUT23), .B1(new_n223), .B2(G119), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT83), .B1(new_n223), .B2(G119), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(G110), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n575), .A2(new_n375), .A3(new_n579), .ZN(new_n580));
  OAI22_X1  g394(.A1(new_n578), .A2(G110), .B1(new_n572), .B2(new_n571), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n368), .A2(new_n211), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(new_n388), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n342), .A2(G221), .A3(G234), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(KEYINPUT84), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT22), .B(G137), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n584), .B(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT25), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(new_n590), .A3(new_n306), .ZN(new_n591));
  INV_X1    g405(.A(G217), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n592), .B1(G234), .B2(new_n306), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(KEYINPUT81), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n590), .B1(new_n589), .B2(new_n306), .ZN(new_n596));
  OR3_X1    g410(.A1(new_n595), .A2(KEYINPUT85), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT85), .B1(new_n595), .B2(new_n596), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n594), .A2(G902), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n589), .A2(new_n599), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n597), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(KEYINPUT86), .B1(new_n570), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n561), .A2(new_n569), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n543), .A2(new_n544), .A3(new_n537), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n544), .B1(new_n543), .B2(new_n537), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT86), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(new_n608), .A3(new_n601), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n475), .B1(new_n603), .B2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(new_n207), .ZN(G3));
  OAI21_X1  g425(.A(G472), .B1(new_n536), .B2(G902), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n543), .A2(new_n537), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n307), .A2(new_n311), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n189), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n614), .A2(new_n602), .A3(new_n616), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n402), .A2(new_n406), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n345), .A2(new_n346), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT33), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT33), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n345), .A2(new_n346), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n620), .A2(G478), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n348), .A2(new_n306), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n347), .B2(new_n348), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n618), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n456), .A2(new_n442), .ZN(new_n629));
  INV_X1    g443(.A(new_n453), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n471), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n628), .A2(new_n631), .A3(new_n470), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n617), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT34), .B(G104), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  NAND2_X1  g449(.A1(new_n394), .A2(new_n398), .ZN(new_n636));
  INV_X1    g450(.A(new_n400), .ZN(new_n637));
  OAI21_X1  g451(.A(KEYINPUT104), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n401), .A2(new_n639), .A3(new_n400), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n641), .B(KEYINPUT103), .C1(new_n400), .C2(new_n401), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT103), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n401), .A2(new_n400), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n638), .B(new_n640), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n353), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n642), .A2(new_n406), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n647), .A2(new_n470), .A3(new_n631), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n617), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT35), .B(G107), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G9));
  XNOR2_X1  g465(.A(new_n584), .B(KEYINPUT105), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT36), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n588), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n652), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n599), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n597), .A2(new_n598), .A3(new_n656), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n312), .A2(new_n474), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n658), .A2(new_n612), .A3(new_n613), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT37), .B(G110), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  OAI211_X1 g475(.A(new_n657), .B(new_n471), .C1(new_n630), .C2(new_n629), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n616), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n342), .A2(G900), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n469), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n666), .A2(KEYINPUT106), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(KEYINPUT106), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n667), .A2(new_n463), .A3(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n647), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n663), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g486(.A(KEYINPUT107), .B1(new_n570), .B2(new_n672), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n663), .A2(new_n671), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT107), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n674), .A2(new_n607), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  XOR2_X1   g492(.A(new_n459), .B(KEYINPUT38), .Z(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n657), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n618), .A2(new_n353), .ZN(new_n682));
  AND4_X1   g496(.A1(new_n471), .A2(new_n680), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n539), .A2(new_n545), .ZN(new_n684));
  INV_X1    g498(.A(new_n556), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n522), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n548), .A2(new_n550), .ZN(new_n687));
  AOI21_X1  g501(.A(G902), .B1(new_n687), .B2(new_n522), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(G472), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n684), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n669), .B(KEYINPUT39), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n312), .A2(new_n692), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n693), .A2(KEYINPUT40), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(KEYINPUT40), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n683), .A2(new_n691), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G143), .ZN(G45));
  NAND2_X1  g511(.A1(new_n627), .A2(new_n669), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n663), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(KEYINPUT108), .B1(new_n570), .B2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n616), .A2(new_n662), .A3(new_n698), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n607), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  AOI21_X1  g520(.A(G902), .B1(new_n302), .B2(new_n303), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n190), .B1(new_n707), .B2(new_n305), .ZN(new_n708));
  OAI21_X1  g522(.A(G469), .B1(new_n707), .B2(KEYINPUT109), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n710));
  AOI211_X1 g524(.A(new_n710), .B(G902), .C1(new_n302), .C2(new_n303), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n708), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(KEYINPUT110), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n714), .B(new_n708), .C1(new_n709), .C2(new_n711), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n713), .A2(new_n632), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n607), .A3(new_n601), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  AND3_X1   g533(.A1(new_n648), .A2(new_n713), .A3(new_n715), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n607), .A3(new_n601), .ZN(new_n721));
  XOR2_X1   g535(.A(KEYINPUT111), .B(G116), .Z(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G18));
  INV_X1    g537(.A(new_n631), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n713), .A2(new_n724), .A3(new_n715), .ZN(new_n725));
  INV_X1    g539(.A(new_n407), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n681), .A2(new_n726), .A3(new_n470), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n725), .A2(new_n607), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G119), .ZN(G21));
  NAND2_X1  g543(.A1(new_n713), .A2(new_n715), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n682), .B(new_n471), .C1(new_n630), .C2(new_n629), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n730), .A2(new_n470), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n560), .B1(new_n543), .B2(new_n306), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n551), .A2(new_n504), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n522), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n538), .B1(new_n540), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT112), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n738), .A3(new_n601), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n738), .B1(new_n737), .B2(new_n601), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n732), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G122), .ZN(G24));
  INV_X1    g557(.A(new_n736), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n612), .A2(new_n657), .A3(new_n699), .A4(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n713), .A2(new_n724), .A3(new_n715), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n366), .ZN(G27));
  NAND2_X1  g562(.A1(G469), .A2(G902), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(KEYINPUT113), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n308), .A2(new_n309), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n305), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n751), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(KEYINPUT114), .B1(new_n752), .B2(new_n305), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(new_n307), .A3(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n459), .A2(new_n472), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n757), .A2(new_n189), .A3(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n607), .A2(new_n601), .A3(new_n699), .A4(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT42), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n602), .B1(new_n684), .B2(new_n604), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n763), .A2(KEYINPUT42), .A3(new_n699), .A4(new_n759), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G131), .ZN(G33));
  NAND4_X1  g580(.A1(new_n607), .A2(new_n601), .A3(new_n671), .A4(new_n759), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G134), .ZN(G36));
  NAND2_X1  g582(.A1(new_n310), .A2(KEYINPUT45), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT45), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n308), .B2(new_n309), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(G469), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT115), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n772), .A2(G469), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n776), .A3(new_n769), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n751), .B1(new_n774), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n307), .B1(new_n778), .B2(KEYINPUT46), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT46), .ZN(new_n780));
  AOI211_X1 g594(.A(new_n780), .B(new_n751), .C1(new_n774), .C2(new_n777), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n189), .B(new_n692), .C1(new_n779), .C2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n626), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n402), .A3(new_n406), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n784), .A2(KEYINPUT116), .A3(KEYINPUT43), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT43), .B1(new_n784), .B2(KEYINPUT116), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n785), .A2(new_n786), .A3(new_n681), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT44), .B1(new_n614), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n782), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n536), .A2(new_n538), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n787), .B(KEYINPUT44), .C1(new_n733), .C2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n758), .B(KEYINPUT117), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n791), .A2(KEYINPUT118), .A3(new_n792), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n789), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G137), .ZN(G39));
  NAND4_X1  g612(.A1(new_n570), .A2(new_n602), .A3(new_n699), .A4(new_n758), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n774), .A2(new_n777), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n780), .B1(new_n801), .B2(new_n751), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n778), .A2(KEYINPUT46), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n307), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT47), .B1(new_n804), .B2(new_n189), .ZN(new_n805));
  OAI211_X1 g619(.A(KEYINPUT47), .B(new_n189), .C1(new_n779), .C2(new_n781), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n800), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G140), .ZN(G42));
  OAI21_X1  g623(.A(new_n307), .B1(new_n709), .B2(new_n711), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n810), .A2(KEYINPUT49), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n601), .A2(new_n189), .A3(new_n471), .ZN(new_n812));
  NOR4_X1   g626(.A1(new_n811), .A2(new_n680), .A3(new_n784), .A4(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n691), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n813), .B(new_n814), .C1(KEYINPUT49), .C2(new_n810), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n737), .A2(new_n601), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT112), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n739), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n785), .A2(new_n786), .A3(new_n463), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n730), .A2(new_n471), .A3(new_n680), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n821), .A2(KEYINPUT50), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n713), .A2(new_n715), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n758), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n463), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n823), .A2(KEYINPUT119), .A3(new_n758), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n733), .A2(new_n681), .A3(new_n736), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n785), .A2(new_n786), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n821), .A2(KEYINPUT50), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n822), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n805), .A2(new_n807), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n834), .B1(new_n189), .B2(new_n810), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n818), .A2(new_n792), .A3(new_n819), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n691), .A2(new_n602), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n828), .A2(new_n618), .A3(new_n626), .A4(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n833), .A2(KEYINPUT51), .A3(new_n837), .A4(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n828), .A2(new_n627), .A3(new_n838), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n818), .A2(new_n725), .A3(new_n819), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n841), .A2(new_n461), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n828), .A2(new_n763), .A3(new_n830), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n844), .A2(KEYINPUT48), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(KEYINPUT48), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n843), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT51), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n837), .A2(new_n839), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n822), .A2(new_n831), .A3(new_n832), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n840), .A2(new_n847), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n570), .A2(KEYINPUT107), .A3(new_n672), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n675), .B1(new_n674), .B2(new_n607), .ZN(new_n855));
  OAI22_X1  g669(.A1(new_n854), .A2(new_n855), .B1(new_n746), .B2(new_n745), .ZN(new_n856));
  INV_X1    g670(.A(new_n731), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n657), .A2(new_n190), .A3(new_n670), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(new_n757), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(new_n684), .B2(new_n690), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n570), .A2(KEYINPUT108), .A3(new_n700), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n702), .B1(new_n607), .B2(new_n703), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT52), .B1(new_n856), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n747), .B1(new_n673), .B2(new_n676), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n860), .B1(new_n701), .B2(new_n704), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT52), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n312), .A2(new_n601), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n402), .A2(new_n406), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n626), .ZN(new_n873));
  AND4_X1   g687(.A1(new_n726), .A2(new_n459), .A3(new_n473), .A4(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n612), .A2(new_n871), .A3(new_n874), .A4(new_n613), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n875), .A2(new_n659), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n717), .A2(new_n721), .A3(new_n728), .A4(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n470), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n823), .A2(new_n878), .A3(new_n857), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n879), .B1(new_n817), .B2(new_n739), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n829), .A2(new_n699), .A3(new_n759), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n758), .A2(new_n353), .A3(new_n657), .A4(new_n669), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n642), .A2(new_n406), .A3(new_n645), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n883), .A2(new_n616), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n607), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n767), .A2(new_n882), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(new_n762), .B2(new_n764), .ZN(new_n888));
  INV_X1    g702(.A(new_n475), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n570), .A2(KEYINPUT86), .A3(new_n602), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n608), .B1(new_n607), .B2(new_n601), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n881), .A2(new_n888), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n870), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n868), .B1(new_n866), .B2(new_n867), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n727), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n684), .B2(new_n604), .ZN(new_n900));
  AOI22_X1  g714(.A1(new_n763), .A2(new_n720), .B1(new_n900), .B2(new_n725), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n875), .A2(new_n659), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n763), .B2(new_n716), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n892), .A2(new_n901), .A3(new_n742), .A4(new_n903), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n767), .A2(new_n882), .A3(new_n886), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n765), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT53), .B1(new_n898), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n853), .B1(new_n895), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n894), .B1(new_n870), .B2(new_n893), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n898), .A2(KEYINPUT53), .A3(new_n907), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n910), .A2(new_n911), .A3(KEYINPUT54), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n852), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n460), .A2(new_n342), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT120), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n815), .B1(new_n913), .B2(new_n915), .ZN(G75));
  NOR2_X1   g730(.A1(new_n342), .A2(G952), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  AOI211_X1 g732(.A(new_n306), .B(new_n458), .C1(new_n910), .C2(new_n911), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n434), .B(new_n440), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT55), .ZN(new_n921));
  XNOR2_X1  g735(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n918), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n910), .A2(new_n911), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n925), .A2(G210), .A3(G902), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT56), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n924), .B1(new_n928), .B2(new_n921), .ZN(G51));
  XNOR2_X1  g743(.A(new_n750), .B(KEYINPUT122), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT57), .Z(new_n931));
  NAND3_X1  g745(.A1(new_n909), .A2(new_n912), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n304), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n925), .A2(G902), .A3(new_n801), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n917), .B1(new_n933), .B2(new_n934), .ZN(G54));
  AND2_X1   g749(.A1(KEYINPUT58), .A2(G475), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n925), .A2(G902), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n937), .A2(new_n393), .A3(new_n386), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n925), .A2(G902), .A3(new_n394), .A4(new_n936), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n938), .A2(new_n918), .A3(new_n939), .ZN(G60));
  NAND2_X1  g754(.A1(new_n620), .A2(new_n622), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n910), .A2(new_n911), .A3(KEYINPUT54), .ZN(new_n942));
  AOI21_X1  g756(.A(KEYINPUT54), .B1(new_n910), .B2(new_n911), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g758(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(new_n624), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n941), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n909), .A2(new_n941), .A3(new_n912), .A4(new_n946), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n918), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n947), .A2(new_n949), .ZN(G63));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n951));
  XNOR2_X1  g765(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n592), .A2(new_n306), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n955), .B1(new_n910), .B2(new_n911), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n918), .B1(new_n956), .B2(new_n589), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n925), .A2(new_n655), .A3(new_n954), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n951), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n925), .A2(new_n954), .ZN(new_n960));
  INV_X1    g774(.A(new_n589), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n956), .A2(new_n655), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n962), .A2(KEYINPUT61), .A3(new_n963), .A4(new_n918), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n959), .A2(new_n964), .ZN(G66));
  OAI22_X1  g779(.A1(new_n466), .A2(new_n467), .B1(G224), .B2(new_n342), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT125), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n877), .A2(new_n610), .A3(new_n880), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n967), .B1(new_n968), .B2(G953), .ZN(new_n969));
  OAI221_X1 g783(.A(new_n427), .B1(G898), .B2(new_n342), .C1(new_n433), .C2(new_n426), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(G69));
  AOI21_X1  g785(.A(new_n664), .B1(new_n192), .B2(G953), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n525), .A2(new_n526), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(new_n389), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n808), .A2(new_n797), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n866), .A2(new_n696), .A3(new_n705), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(KEYINPUT62), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT62), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n866), .A2(new_n978), .A3(new_n696), .A4(new_n705), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n758), .A2(new_n726), .A3(new_n873), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n693), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(new_n890), .B2(new_n891), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n975), .A2(new_n977), .A3(new_n979), .A4(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n974), .B1(new_n983), .B2(new_n342), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n763), .A2(new_n857), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n767), .B1(new_n985), .B2(new_n782), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n986), .B1(new_n762), .B2(new_n764), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n866), .A2(new_n705), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n975), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n664), .B1(new_n989), .B2(new_n342), .ZN(new_n990));
  INV_X1    g804(.A(new_n974), .ZN(new_n991));
  OAI22_X1  g805(.A1(new_n984), .A2(KEYINPUT126), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n984), .A2(KEYINPUT126), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n972), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OR2_X1    g808(.A1(new_n984), .A2(KEYINPUT126), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n984), .A2(KEYINPUT126), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n990), .A2(new_n991), .ZN(new_n997));
  INV_X1    g811(.A(new_n972), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n995), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n994), .A2(new_n999), .ZN(G72));
  NAND2_X1  g814(.A1(G472), .A2(G902), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT63), .Z(new_n1002));
  INV_X1    g816(.A(KEYINPUT127), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n531), .A2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(new_n564), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n925), .A2(new_n1002), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n686), .ZN(new_n1007));
  OR2_X1    g821(.A1(new_n983), .A2(new_n904), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1007), .B1(new_n1008), .B2(new_n1002), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n685), .A2(new_n522), .ZN(new_n1010));
  OR2_X1    g824(.A1(new_n989), .A2(new_n904), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1010), .B1(new_n1011), .B2(new_n1002), .ZN(new_n1012));
  NOR4_X1   g826(.A1(new_n1006), .A2(new_n1009), .A3(new_n1012), .A4(new_n917), .ZN(G57));
endmodule


