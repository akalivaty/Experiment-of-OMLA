

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745;

  INV_X1 U369 ( .A(n357), .ZN(n348) );
  INV_X1 U370 ( .A(n556), .ZN(n350) );
  NAND2_X1 U371 ( .A1(n419), .A2(n418), .ZN(n417) );
  NOR2_X1 U372 ( .A1(n665), .A2(n664), .ZN(n600) );
  XNOR2_X1 U373 ( .A(n560), .B(n559), .ZN(n665) );
  XNOR2_X1 U374 ( .A(n431), .B(n430), .ZN(n596) );
  XNOR2_X1 U375 ( .A(n441), .B(n439), .ZN(n563) );
  XNOR2_X1 U376 ( .A(n503), .B(n502), .ZN(n372) );
  XNOR2_X1 U377 ( .A(n500), .B(n499), .ZN(n503) );
  XNOR2_X1 U378 ( .A(n480), .B(G134), .ZN(n500) );
  NOR2_X2 U379 ( .A1(n635), .A2(n354), .ZN(n422) );
  NOR2_X1 U380 ( .A1(n349), .A2(n348), .ZN(n377) );
  INV_X1 U381 ( .A(n379), .ZN(n349) );
  NAND2_X1 U382 ( .A1(n653), .A2(n638), .ZN(n607) );
  XNOR2_X1 U383 ( .A(n602), .B(KEYINPUT31), .ZN(n653) );
  XNOR2_X2 U384 ( .A(n598), .B(KEYINPUT33), .ZN(n690) );
  INV_X1 U385 ( .A(n364), .ZN(n743) );
  NAND2_X1 U386 ( .A1(n362), .A2(n364), .ZN(n361) );
  XNOR2_X2 U387 ( .A(n428), .B(n350), .ZN(n364) );
  XNOR2_X1 U388 ( .A(G110), .B(G128), .ZN(n521) );
  NOR2_X1 U389 ( .A1(n564), .A2(n563), .ZN(n579) );
  XOR2_X1 U390 ( .A(n596), .B(KEYINPUT107), .Z(n351) );
  NOR2_X1 U391 ( .A1(n675), .A2(n603), .ZN(n602) );
  NOR2_X2 U392 ( .A1(n742), .A2(n642), .ZN(n385) );
  XNOR2_X2 U393 ( .A(n594), .B(KEYINPUT32), .ZN(n742) );
  NOR2_X2 U394 ( .A1(n680), .A2(n681), .ZN(n544) );
  AND2_X2 U395 ( .A1(n593), .A2(n398), .ZN(n594) );
  XNOR2_X2 U396 ( .A(n589), .B(n410), .ZN(n593) );
  XOR2_X1 U397 ( .A(KEYINPUT6), .B(n671), .Z(n597) );
  INV_X2 U398 ( .A(n606), .ZN(n671) );
  INV_X1 U399 ( .A(n745), .ZN(n362) );
  NAND2_X1 U400 ( .A1(n650), .A2(n654), .ZN(n686) );
  BUF_X1 U401 ( .A(n575), .Z(n415) );
  NOR2_X2 U402 ( .A1(n473), .A2(n563), .ZN(n647) );
  OR2_X1 U403 ( .A1(n626), .A2(G902), .ZN(n448) );
  NAND2_X1 U404 ( .A1(n377), .A2(n376), .ZN(n433) );
  NOR2_X1 U405 ( .A1(n717), .A2(n622), .ZN(n625) );
  NOR2_X1 U406 ( .A1(n671), .A2(n590), .ZN(n642) );
  XNOR2_X1 U407 ( .A(n561), .B(KEYINPUT111), .ZN(n739) );
  NOR2_X1 U408 ( .A1(n565), .A2(n680), .ZN(n555) );
  NOR2_X1 U409 ( .A1(n572), .A2(n415), .ZN(n558) );
  AND2_X1 U410 ( .A1(n592), .A2(n399), .ZN(n398) );
  NOR2_X1 U411 ( .A1(n591), .A2(n435), .ZN(n434) );
  NAND2_X1 U412 ( .A1(n600), .A2(n597), .ZN(n598) );
  XNOR2_X1 U413 ( .A(n551), .B(KEYINPUT98), .ZN(n604) );
  OR2_X1 U414 ( .A1(n557), .A2(n681), .ZN(n435) );
  XNOR2_X1 U415 ( .A(n472), .B(n471), .ZN(n712) );
  XNOR2_X1 U416 ( .A(n411), .B(n474), .ZN(n498) );
  XNOR2_X1 U417 ( .A(n382), .B(KEYINPUT3), .ZN(n411) );
  XNOR2_X1 U418 ( .A(n508), .B(G472), .ZN(n447) );
  INV_X1 U419 ( .A(G469), .ZN(n421) );
  XNOR2_X1 U420 ( .A(G113), .B(G101), .ZN(n474) );
  BUF_X1 U421 ( .A(n609), .Z(n352) );
  NOR2_X1 U422 ( .A1(G953), .A2(G237), .ZN(n505) );
  INV_X1 U423 ( .A(KEYINPUT72), .ZN(n412) );
  XNOR2_X1 U424 ( .A(KEYINPUT96), .B(KEYINPUT20), .ZN(n509) );
  XNOR2_X1 U425 ( .A(n437), .B(G116), .ZN(n478) );
  XNOR2_X1 U426 ( .A(G107), .B(G122), .ZN(n437) );
  INV_X1 U427 ( .A(KEYINPUT92), .ZN(n427) );
  AND2_X1 U428 ( .A1(n356), .A2(n570), .ZN(n369) );
  INV_X1 U429 ( .A(KEYINPUT83), .ZN(n424) );
  XNOR2_X1 U430 ( .A(n693), .B(n394), .ZN(n694) );
  XNOR2_X1 U431 ( .A(n395), .B(KEYINPUT118), .ZN(n394) );
  XNOR2_X1 U432 ( .A(n544), .B(KEYINPUT110), .ZN(n685) );
  XNOR2_X1 U433 ( .A(n387), .B(n386), .ZN(n552) );
  INV_X1 U434 ( .A(KEYINPUT30), .ZN(n386) );
  XNOR2_X1 U435 ( .A(n491), .B(n490), .ZN(n492) );
  INV_X1 U436 ( .A(KEYINPUT74), .ZN(n490) );
  XNOR2_X1 U437 ( .A(n498), .B(n507), .ZN(n406) );
  XNOR2_X1 U438 ( .A(n390), .B(n389), .ZN(n526) );
  INV_X1 U439 ( .A(KEYINPUT8), .ZN(n389) );
  XNOR2_X1 U440 ( .A(n469), .B(KEYINPUT9), .ZN(n438) );
  XOR2_X1 U441 ( .A(KEYINPUT104), .B(KEYINPUT7), .Z(n469) );
  NAND2_X1 U442 ( .A1(n621), .A2(n442), .ZN(n445) );
  NAND2_X1 U443 ( .A1(n619), .A2(n618), .ZN(n621) );
  NOR2_X1 U444 ( .A1(n661), .A2(n446), .ZN(n442) );
  XNOR2_X1 U445 ( .A(n531), .B(KEYINPUT25), .ZN(n430) );
  OR2_X1 U446 ( .A1(n715), .A2(G902), .ZN(n431) );
  INV_X1 U447 ( .A(KEYINPUT22), .ZN(n410) );
  XNOR2_X1 U448 ( .A(n440), .B(G478), .ZN(n439) );
  OR2_X1 U449 ( .A1(n712), .A2(G902), .ZN(n441) );
  INV_X1 U450 ( .A(KEYINPUT105), .ZN(n440) );
  BUF_X1 U451 ( .A(n733), .Z(n407) );
  XNOR2_X1 U452 ( .A(n413), .B(n477), .ZN(n375) );
  XNOR2_X1 U453 ( .A(n498), .B(n479), .ZN(n413) );
  XOR2_X1 U454 ( .A(KEYINPUT16), .B(KEYINPUT71), .Z(n476) );
  XNOR2_X1 U455 ( .A(n451), .B(n538), .ZN(n426) );
  NOR2_X1 U456 ( .A1(n407), .A2(G952), .ZN(n717) );
  OR2_X1 U457 ( .A1(n353), .A2(KEYINPUT121), .ZN(n378) );
  INV_X1 U458 ( .A(KEYINPUT46), .ZN(n371) );
  INV_X1 U459 ( .A(G125), .ZN(n453) );
  INV_X1 U460 ( .A(KEYINPUT52), .ZN(n395) );
  OR2_X1 U461 ( .A1(G237), .A2(G902), .ZN(n494) );
  XNOR2_X1 U462 ( .A(G116), .B(G146), .ZN(n504) );
  XOR2_X1 U463 ( .A(KEYINPUT12), .B(KEYINPUT102), .Z(n457) );
  XNOR2_X1 U464 ( .A(G104), .B(G143), .ZN(n456) );
  XOR2_X1 U465 ( .A(KEYINPUT11), .B(KEYINPUT101), .Z(n460) );
  XNOR2_X1 U466 ( .A(G122), .B(G113), .ZN(n462) );
  XNOR2_X1 U467 ( .A(n482), .B(n404), .ZN(n730) );
  XNOR2_X1 U468 ( .A(KEYINPUT10), .B(G140), .ZN(n404) );
  INV_X1 U469 ( .A(G137), .ZN(n499) );
  INV_X1 U470 ( .A(KEYINPUT48), .ZN(n429) );
  AND2_X1 U471 ( .A1(n571), .A2(n369), .ZN(n368) );
  XNOR2_X1 U472 ( .A(n611), .B(KEYINPUT45), .ZN(n612) );
  INV_X1 U473 ( .A(KEYINPUT80), .ZN(n611) );
  XNOR2_X1 U474 ( .A(KEYINPUT21), .B(n512), .ZN(n667) );
  XNOR2_X1 U475 ( .A(G119), .B(G137), .ZN(n527) );
  XNOR2_X1 U476 ( .A(n730), .B(n409), .ZN(n408) );
  INV_X1 U477 ( .A(KEYINPUT93), .ZN(n409) );
  XNOR2_X1 U478 ( .A(G104), .B(KEYINPUT87), .ZN(n475) );
  XNOR2_X1 U479 ( .A(G107), .B(G101), .ZN(n534) );
  XOR2_X1 U480 ( .A(G140), .B(G146), .Z(n535) );
  NOR2_X1 U481 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U482 ( .A(n546), .B(n545), .ZN(n663) );
  XNOR2_X1 U483 ( .A(n384), .B(n553), .ZN(n565) );
  NOR2_X1 U484 ( .A1(n552), .A2(n549), .ZN(n397) );
  XNOR2_X1 U485 ( .A(KEYINPUT66), .B(KEYINPUT19), .ZN(n496) );
  XNOR2_X1 U486 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U487 ( .A(n388), .B(n529), .ZN(n715) );
  XNOR2_X1 U488 ( .A(n408), .B(n525), .ZN(n529) );
  XNOR2_X1 U489 ( .A(n528), .B(n527), .ZN(n388) );
  XNOR2_X1 U490 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U491 ( .A(n438), .B(n478), .ZN(n470) );
  XNOR2_X1 U492 ( .A(n443), .B(n359), .ZN(n622) );
  NOR2_X1 U493 ( .A1(n445), .A2(n444), .ZN(n443) );
  INV_X1 U494 ( .A(G475), .ZN(n444) );
  XNOR2_X1 U495 ( .A(n375), .B(n489), .ZN(n702) );
  INV_X1 U496 ( .A(KEYINPUT35), .ZN(n416) );
  INV_X1 U497 ( .A(n599), .ZN(n418) );
  AND2_X1 U498 ( .A1(n400), .A2(n596), .ZN(n391) );
  AND2_X1 U499 ( .A1(n414), .A2(n383), .ZN(n635) );
  NOR2_X1 U500 ( .A1(n399), .A2(n351), .ZN(n383) );
  INV_X1 U501 ( .A(KEYINPUT82), .ZN(n392) );
  XNOR2_X1 U502 ( .A(n707), .B(n401), .ZN(n710) );
  INV_X1 U503 ( .A(KEYINPUT53), .ZN(n432) );
  XNOR2_X1 U504 ( .A(n495), .B(KEYINPUT89), .ZN(n681) );
  XNOR2_X1 U505 ( .A(KEYINPUT120), .B(n699), .ZN(n353) );
  INV_X1 U506 ( .A(n595), .ZN(n603) );
  AND2_X1 U507 ( .A1(n607), .A2(n686), .ZN(n354) );
  AND2_X1 U508 ( .A1(n657), .A2(n656), .ZN(n355) );
  BUF_X1 U509 ( .A(n665), .Z(n400) );
  INV_X1 U510 ( .A(n400), .ZN(n399) );
  NAND2_X1 U511 ( .A1(n543), .A2(n542), .ZN(n356) );
  AND2_X1 U512 ( .A1(n378), .A2(n582), .ZN(n357) );
  XNOR2_X1 U513 ( .A(KEYINPUT69), .B(KEYINPUT34), .ZN(n358) );
  XNOR2_X1 U514 ( .A(n466), .B(KEYINPUT59), .ZN(n359) );
  XOR2_X1 U515 ( .A(G902), .B(KEYINPUT15), .Z(n620) );
  NOR2_X1 U516 ( .A1(n375), .A2(n718), .ZN(n360) );
  NAND2_X1 U517 ( .A1(n361), .A2(n371), .ZN(n366) );
  NAND2_X1 U518 ( .A1(n366), .A2(n363), .ZN(n370) );
  NAND2_X1 U519 ( .A1(n365), .A2(n364), .ZN(n363) );
  NOR2_X1 U520 ( .A1(n745), .A2(n371), .ZN(n365) );
  XNOR2_X2 U521 ( .A(n367), .B(n429), .ZN(n436) );
  NAND2_X1 U522 ( .A1(n370), .A2(n368), .ZN(n367) );
  XNOR2_X1 U523 ( .A(n406), .B(n372), .ZN(n626) );
  XNOR2_X2 U524 ( .A(n372), .B(n427), .ZN(n729) );
  NAND2_X1 U525 ( .A1(n385), .A2(n373), .ZN(n609) );
  XNOR2_X1 U526 ( .A(n373), .B(n741), .ZN(G24) );
  XNOR2_X2 U527 ( .A(n417), .B(n416), .ZN(n373) );
  NOR2_X2 U528 ( .A1(n374), .A2(n587), .ZN(n405) );
  NOR2_X1 U529 ( .A1(n547), .A2(n374), .ZN(n648) );
  XNOR2_X1 U530 ( .A(n497), .B(n496), .ZN(n374) );
  OR2_X1 U531 ( .A1(n381), .A2(KEYINPUT121), .ZN(n376) );
  NAND2_X1 U532 ( .A1(n381), .A2(n380), .ZN(n379) );
  AND2_X1 U533 ( .A1(n353), .A2(KEYINPUT121), .ZN(n380) );
  XNOR2_X1 U534 ( .A(n662), .B(KEYINPUT79), .ZN(n381) );
  XNOR2_X2 U535 ( .A(G119), .B(KEYINPUT88), .ZN(n382) );
  XNOR2_X2 U536 ( .A(KEYINPUT42), .B(n548), .ZN(n745) );
  NOR2_X2 U537 ( .A1(n615), .A2(n616), .ZN(n661) );
  XNOR2_X1 U538 ( .A(n555), .B(n554), .ZN(n577) );
  INV_X1 U539 ( .A(n604), .ZN(n396) );
  NAND2_X1 U540 ( .A1(n396), .A2(n397), .ZN(n384) );
  NOR2_X1 U541 ( .A1(n606), .A2(n681), .ZN(n387) );
  NAND2_X1 U542 ( .A1(n733), .A2(G234), .ZN(n390) );
  NAND2_X1 U543 ( .A1(n593), .A2(n391), .ZN(n590) );
  NOR2_X2 U544 ( .A1(n663), .A2(n547), .ZN(n548) );
  XNOR2_X1 U545 ( .A(n420), .B(n358), .ZN(n419) );
  XNOR2_X1 U546 ( .A(n393), .B(n392), .ZN(n414) );
  NAND2_X1 U547 ( .A1(n593), .A2(n591), .ZN(n393) );
  XNOR2_X2 U548 ( .A(n566), .B(KEYINPUT38), .ZN(n680) );
  NAND2_X1 U549 ( .A1(n595), .A2(n588), .ZN(n589) );
  XNOR2_X2 U550 ( .A(n405), .B(KEYINPUT0), .ZN(n595) );
  NOR2_X2 U551 ( .A1(n631), .A2(n717), .ZN(n634) );
  XNOR2_X1 U552 ( .A(n709), .B(n708), .ZN(n401) );
  XNOR2_X1 U553 ( .A(n402), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U554 ( .A1(n705), .A2(n717), .ZN(n402) );
  NAND2_X1 U555 ( .A1(n403), .A2(n399), .ZN(n561) );
  XNOR2_X1 U556 ( .A(n558), .B(KEYINPUT36), .ZN(n403) );
  NAND2_X1 U557 ( .A1(n647), .A2(n434), .ZN(n572) );
  INV_X1 U558 ( .A(n620), .ZN(n446) );
  INV_X2 U559 ( .A(n445), .ZN(n706) );
  XNOR2_X1 U560 ( .A(n493), .B(n492), .ZN(n575) );
  XNOR2_X1 U561 ( .A(n425), .B(n424), .ZN(n423) );
  NOR2_X1 U562 ( .A1(n660), .A2(n661), .ZN(n662) );
  NOR2_X1 U563 ( .A1(n719), .A2(n731), .ZN(n659) );
  NAND2_X2 U564 ( .A1(n436), .A2(n355), .ZN(n731) );
  NAND2_X1 U565 ( .A1(n658), .A2(n614), .ZN(n615) );
  XNOR2_X2 U566 ( .A(n613), .B(n612), .ZN(n658) );
  XNOR2_X1 U567 ( .A(n731), .B(n412), .ZN(n617) );
  NOR2_X2 U568 ( .A1(n423), .A2(n610), .ZN(n613) );
  XNOR2_X2 U569 ( .A(G143), .B(G128), .ZN(n480) );
  NAND2_X1 U570 ( .A1(n690), .A2(n595), .ZN(n420) );
  XNOR2_X2 U571 ( .A(n539), .B(n421), .ZN(n560) );
  NAND2_X1 U572 ( .A1(n608), .A2(n422), .ZN(n425) );
  XNOR2_X2 U573 ( .A(n729), .B(n426), .ZN(n709) );
  NAND2_X1 U574 ( .A1(n577), .A2(n647), .ZN(n428) );
  XNOR2_X1 U575 ( .A(n433), .B(n432), .ZN(G75) );
  NAND2_X1 U576 ( .A1(n436), .A2(n657), .ZN(n616) );
  XNOR2_X2 U577 ( .A(n448), .B(n447), .ZN(n606) );
  XNOR2_X1 U578 ( .A(n630), .B(n629), .ZN(n631) );
  XOR2_X1 U579 ( .A(n701), .B(n700), .Z(n449) );
  AND2_X1 U580 ( .A1(n505), .A2(G210), .ZN(n450) );
  XOR2_X1 U581 ( .A(n537), .B(n536), .Z(n451) );
  XNOR2_X1 U582 ( .A(n506), .B(n450), .ZN(n507) );
  XNOR2_X1 U583 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U584 ( .A(n486), .B(n485), .ZN(n488) );
  XNOR2_X1 U585 ( .A(n538), .B(n476), .ZN(n477) );
  INV_X1 U586 ( .A(KEYINPUT41), .ZN(n545) );
  INV_X1 U587 ( .A(KEYINPUT73), .ZN(n553) );
  INV_X1 U588 ( .A(KEYINPUT63), .ZN(n632) );
  INV_X1 U589 ( .A(KEYINPUT60), .ZN(n623) );
  XNOR2_X1 U590 ( .A(n632), .B(KEYINPUT84), .ZN(n633) );
  XNOR2_X1 U591 ( .A(n623), .B(KEYINPUT67), .ZN(n624) );
  XOR2_X2 U592 ( .A(G953), .B(KEYINPUT64), .Z(n733) );
  INV_X1 U593 ( .A(G146), .ZN(n452) );
  NAND2_X1 U594 ( .A1(n452), .A2(G125), .ZN(n455) );
  NAND2_X1 U595 ( .A1(n453), .A2(G146), .ZN(n454) );
  NAND2_X1 U596 ( .A1(n455), .A2(n454), .ZN(n482) );
  XNOR2_X1 U597 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U598 ( .A(n730), .B(n458), .ZN(n465) );
  NAND2_X1 U599 ( .A1(n505), .A2(G214), .ZN(n459) );
  XNOR2_X1 U600 ( .A(n460), .B(n459), .ZN(n461) );
  XOR2_X1 U601 ( .A(n461), .B(G131), .Z(n463) );
  XNOR2_X1 U602 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U603 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U604 ( .A(KEYINPUT13), .B(G475), .ZN(n468) );
  NOR2_X1 U605 ( .A1(G902), .A2(n466), .ZN(n467) );
  XNOR2_X1 U606 ( .A(n468), .B(n467), .ZN(n564) );
  XNOR2_X1 U607 ( .A(n564), .B(KEYINPUT103), .ZN(n473) );
  XOR2_X1 U608 ( .A(n500), .B(n470), .Z(n472) );
  NAND2_X1 U609 ( .A1(G217), .A2(n526), .ZN(n471) );
  INV_X1 U610 ( .A(n647), .ZN(n650) );
  NAND2_X1 U611 ( .A1(n563), .A2(n473), .ZN(n654) );
  XNOR2_X1 U612 ( .A(n475), .B(G110), .ZN(n538) );
  INV_X1 U613 ( .A(n478), .ZN(n479) );
  XOR2_X1 U614 ( .A(KEYINPUT4), .B(KEYINPUT65), .Z(n501) );
  INV_X1 U615 ( .A(n480), .ZN(n481) );
  XOR2_X1 U616 ( .A(n501), .B(n481), .Z(n486) );
  NAND2_X1 U617 ( .A1(G224), .A2(n733), .ZN(n484) );
  INV_X1 U618 ( .A(n482), .ZN(n483) );
  XNOR2_X1 U619 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n487) );
  XNOR2_X1 U620 ( .A(n488), .B(n487), .ZN(n489) );
  NOR2_X1 U621 ( .A1(n702), .A2(n620), .ZN(n493) );
  NAND2_X1 U622 ( .A1(G210), .A2(n494), .ZN(n491) );
  NAND2_X1 U623 ( .A1(n494), .A2(G214), .ZN(n495) );
  NOR2_X1 U624 ( .A1(n575), .A2(n681), .ZN(n497) );
  XNOR2_X1 U625 ( .A(n501), .B(G131), .ZN(n502) );
  XNOR2_X1 U626 ( .A(n504), .B(KEYINPUT5), .ZN(n506) );
  XNOR2_X1 U627 ( .A(KEYINPUT70), .B(KEYINPUT99), .ZN(n508) );
  NAND2_X1 U628 ( .A1(n446), .A2(G234), .ZN(n510) );
  XNOR2_X1 U629 ( .A(n510), .B(n509), .ZN(n530) );
  NAND2_X1 U630 ( .A1(n530), .A2(G221), .ZN(n511) );
  XOR2_X1 U631 ( .A(KEYINPUT97), .B(n511), .Z(n512) );
  NAND2_X1 U632 ( .A1(G234), .A2(G237), .ZN(n513) );
  XNOR2_X1 U633 ( .A(n513), .B(KEYINPUT14), .ZN(n515) );
  NAND2_X1 U634 ( .A1(n515), .A2(G952), .ZN(n514) );
  XNOR2_X1 U635 ( .A(KEYINPUT90), .B(n514), .ZN(n695) );
  NOR2_X1 U636 ( .A1(G953), .A2(n695), .ZN(n581) );
  INV_X1 U637 ( .A(n407), .ZN(n516) );
  AND2_X1 U638 ( .A1(G902), .A2(n515), .ZN(n583) );
  NAND2_X1 U639 ( .A1(n516), .A2(n583), .ZN(n517) );
  NOR2_X1 U640 ( .A1(G900), .A2(n517), .ZN(n518) );
  NOR2_X1 U641 ( .A1(n581), .A2(n518), .ZN(n519) );
  XOR2_X1 U642 ( .A(KEYINPUT75), .B(n519), .Z(n549) );
  NOR2_X1 U643 ( .A1(n667), .A2(n549), .ZN(n520) );
  XNOR2_X1 U644 ( .A(KEYINPUT68), .B(n520), .ZN(n532) );
  XOR2_X1 U645 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n522) );
  XNOR2_X1 U646 ( .A(n522), .B(n521), .ZN(n524) );
  XOR2_X1 U647 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n523) );
  NAND2_X1 U648 ( .A1(n526), .A2(G221), .ZN(n528) );
  NAND2_X1 U649 ( .A1(G217), .A2(n530), .ZN(n531) );
  NAND2_X1 U650 ( .A1(n532), .A2(n596), .ZN(n557) );
  NOR2_X1 U651 ( .A1(n606), .A2(n557), .ZN(n533) );
  XNOR2_X1 U652 ( .A(KEYINPUT28), .B(n533), .ZN(n540) );
  XNOR2_X1 U653 ( .A(n535), .B(n534), .ZN(n537) );
  NAND2_X1 U654 ( .A1(G227), .A2(n733), .ZN(n536) );
  NOR2_X2 U655 ( .A1(G902), .A2(n709), .ZN(n539) );
  NAND2_X1 U656 ( .A1(n540), .A2(n560), .ZN(n547) );
  NAND2_X1 U657 ( .A1(n686), .A2(n648), .ZN(n541) );
  INV_X1 U658 ( .A(KEYINPUT47), .ZN(n562) );
  NAND2_X1 U659 ( .A1(n541), .A2(n562), .ZN(n543) );
  NAND2_X1 U660 ( .A1(n648), .A2(KEYINPUT47), .ZN(n542) );
  INV_X1 U661 ( .A(n415), .ZN(n566) );
  NAND2_X1 U662 ( .A1(n685), .A2(n579), .ZN(n546) );
  XNOR2_X1 U663 ( .A(KEYINPUT40), .B(KEYINPUT109), .ZN(n556) );
  NOR2_X1 U664 ( .A1(n667), .A2(n596), .ZN(n550) );
  NAND2_X1 U665 ( .A1(n550), .A2(n560), .ZN(n551) );
  INV_X1 U666 ( .A(KEYINPUT39), .ZN(n554) );
  INV_X1 U667 ( .A(n597), .ZN(n591) );
  INV_X1 U668 ( .A(KEYINPUT1), .ZN(n559) );
  XNOR2_X1 U669 ( .A(n739), .B(KEYINPUT81), .ZN(n571) );
  OR2_X1 U670 ( .A1(n562), .A2(n686), .ZN(n568) );
  NAND2_X1 U671 ( .A1(n564), .A2(n563), .ZN(n599) );
  NOR2_X1 U672 ( .A1(n565), .A2(n599), .ZN(n567) );
  NAND2_X1 U673 ( .A1(n567), .A2(n566), .ZN(n646) );
  NAND2_X1 U674 ( .A1(n568), .A2(n646), .ZN(n569) );
  XNOR2_X1 U675 ( .A(n569), .B(KEYINPUT77), .ZN(n570) );
  XOR2_X1 U676 ( .A(n572), .B(KEYINPUT108), .Z(n573) );
  NAND2_X1 U677 ( .A1(n573), .A2(n400), .ZN(n574) );
  XNOR2_X1 U678 ( .A(KEYINPUT43), .B(n574), .ZN(n576) );
  NAND2_X1 U679 ( .A1(n576), .A2(n415), .ZN(n657) );
  INV_X1 U680 ( .A(n654), .ZN(n643) );
  NAND2_X1 U681 ( .A1(n577), .A2(n643), .ZN(n656) );
  NAND2_X1 U682 ( .A1(KEYINPUT2), .A2(n656), .ZN(n578) );
  XOR2_X1 U683 ( .A(KEYINPUT76), .B(n578), .Z(n614) );
  INV_X1 U684 ( .A(n579), .ZN(n683) );
  NOR2_X1 U685 ( .A1(n667), .A2(n683), .ZN(n580) );
  XNOR2_X1 U686 ( .A(KEYINPUT106), .B(n580), .ZN(n588) );
  INV_X1 U687 ( .A(n581), .ZN(n585) );
  INV_X1 U688 ( .A(G953), .ZN(n582) );
  NOR2_X1 U689 ( .A1(G898), .A2(n582), .ZN(n718) );
  NAND2_X1 U690 ( .A1(n583), .A2(n718), .ZN(n584) );
  NAND2_X1 U691 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U692 ( .A(KEYINPUT91), .B(n586), .ZN(n587) );
  AND2_X1 U693 ( .A1(n351), .A2(n591), .ZN(n592) );
  OR2_X1 U694 ( .A1(n667), .A2(n596), .ZN(n664) );
  NAND2_X1 U695 ( .A1(n609), .A2(KEYINPUT44), .ZN(n608) );
  NAND2_X1 U696 ( .A1(n671), .A2(n600), .ZN(n601) );
  XNOR2_X1 U697 ( .A(n601), .B(KEYINPUT100), .ZN(n675) );
  NOR2_X1 U698 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U699 ( .A1(n606), .A2(n605), .ZN(n638) );
  NOR2_X1 U700 ( .A1(n352), .A2(KEYINPUT44), .ZN(n610) );
  NAND2_X1 U701 ( .A1(n658), .A2(n617), .ZN(n619) );
  INV_X1 U702 ( .A(KEYINPUT2), .ZN(n618) );
  XNOR2_X1 U703 ( .A(n625), .B(n624), .ZN(G60) );
  NAND2_X1 U704 ( .A1(n706), .A2(G472), .ZN(n630) );
  XOR2_X1 U705 ( .A(n626), .B(KEYINPUT112), .Z(n628) );
  XOR2_X1 U706 ( .A(KEYINPUT62), .B(KEYINPUT86), .Z(n627) );
  XNOR2_X1 U707 ( .A(n634), .B(n633), .ZN(G57) );
  XNOR2_X1 U708 ( .A(n635), .B(G101), .ZN(n636) );
  XNOR2_X1 U709 ( .A(n636), .B(KEYINPUT113), .ZN(G3) );
  NOR2_X1 U710 ( .A1(n650), .A2(n638), .ZN(n637) );
  XOR2_X1 U711 ( .A(G104), .B(n637), .Z(G6) );
  NOR2_X1 U712 ( .A1(n654), .A2(n638), .ZN(n640) );
  XNOR2_X1 U713 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n639) );
  XNOR2_X1 U714 ( .A(n640), .B(n639), .ZN(n641) );
  XNOR2_X1 U715 ( .A(G107), .B(n641), .ZN(G9) );
  XOR2_X1 U716 ( .A(n642), .B(G110), .Z(G12) );
  XOR2_X1 U717 ( .A(G128), .B(KEYINPUT29), .Z(n645) );
  NAND2_X1 U718 ( .A1(n648), .A2(n643), .ZN(n644) );
  XNOR2_X1 U719 ( .A(n645), .B(n644), .ZN(G30) );
  XNOR2_X1 U720 ( .A(G143), .B(n646), .ZN(G45) );
  NAND2_X1 U721 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U722 ( .A(n649), .B(G146), .ZN(G48) );
  NOR2_X1 U723 ( .A1(n650), .A2(n653), .ZN(n651) );
  XOR2_X1 U724 ( .A(KEYINPUT114), .B(n651), .Z(n652) );
  XNOR2_X1 U725 ( .A(G113), .B(n652), .ZN(G15) );
  NOR2_X1 U726 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U727 ( .A(G116), .B(n655), .Z(G18) );
  XNOR2_X1 U728 ( .A(G134), .B(n656), .ZN(G36) );
  XNOR2_X1 U729 ( .A(G140), .B(n657), .ZN(G42) );
  INV_X1 U730 ( .A(n658), .ZN(n719) );
  NOR2_X1 U731 ( .A1(n659), .A2(KEYINPUT2), .ZN(n660) );
  INV_X1 U732 ( .A(n663), .ZN(n679) );
  AND2_X1 U733 ( .A1(n690), .A2(n679), .ZN(n698) );
  XOR2_X1 U734 ( .A(KEYINPUT51), .B(KEYINPUT116), .Z(n677) );
  NAND2_X1 U735 ( .A1(n400), .A2(n664), .ZN(n666) );
  XNOR2_X1 U736 ( .A(KEYINPUT50), .B(n666), .ZN(n673) );
  XNOR2_X1 U737 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n669) );
  NAND2_X1 U738 ( .A1(n351), .A2(n667), .ZN(n668) );
  XOR2_X1 U739 ( .A(n669), .B(n668), .Z(n670) );
  NOR2_X1 U740 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U741 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U742 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U743 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U744 ( .A1(n679), .A2(n678), .ZN(n692) );
  AND2_X1 U745 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U746 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U747 ( .A(n684), .B(KEYINPUT117), .ZN(n688) );
  NAND2_X1 U748 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U749 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U750 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U751 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U752 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U753 ( .A(KEYINPUT119), .B(n696), .Z(n697) );
  NAND2_X1 U754 ( .A1(n706), .A2(G210), .ZN(n704) );
  XOR2_X1 U755 ( .A(KEYINPUT55), .B(KEYINPUT54), .Z(n701) );
  XNOR2_X1 U756 ( .A(KEYINPUT85), .B(KEYINPUT78), .ZN(n700) );
  XNOR2_X1 U757 ( .A(n702), .B(n449), .ZN(n703) );
  XNOR2_X1 U758 ( .A(n704), .B(n703), .ZN(n705) );
  XOR2_X1 U759 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n708) );
  NAND2_X1 U760 ( .A1(n706), .A2(G469), .ZN(n707) );
  NOR2_X1 U761 ( .A1(n717), .A2(n710), .ZN(G54) );
  NAND2_X1 U762 ( .A1(G478), .A2(n706), .ZN(n711) );
  XNOR2_X1 U763 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U764 ( .A1(n717), .A2(n713), .ZN(G63) );
  NAND2_X1 U765 ( .A1(G217), .A2(n706), .ZN(n714) );
  XNOR2_X1 U766 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U767 ( .A1(n717), .A2(n716), .ZN(G66) );
  NOR2_X1 U768 ( .A1(G953), .A2(n719), .ZN(n720) );
  XNOR2_X1 U769 ( .A(KEYINPUT125), .B(n720), .ZN(n727) );
  XOR2_X1 U770 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n722) );
  NAND2_X1 U771 ( .A1(G224), .A2(G953), .ZN(n721) );
  XNOR2_X1 U772 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U773 ( .A(KEYINPUT122), .B(n723), .ZN(n724) );
  NAND2_X1 U774 ( .A1(n724), .A2(G898), .ZN(n725) );
  XNOR2_X1 U775 ( .A(KEYINPUT124), .B(n725), .ZN(n726) );
  NAND2_X1 U776 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U777 ( .A(n360), .B(n728), .ZN(G69) );
  XNOR2_X1 U778 ( .A(n729), .B(n730), .ZN(n734) );
  XNOR2_X1 U779 ( .A(n731), .B(n734), .ZN(n732) );
  NAND2_X1 U780 ( .A1(n407), .A2(n732), .ZN(n738) );
  XNOR2_X1 U781 ( .A(G227), .B(n734), .ZN(n735) );
  NAND2_X1 U782 ( .A1(n735), .A2(G900), .ZN(n736) );
  NAND2_X1 U783 ( .A1(G953), .A2(n736), .ZN(n737) );
  NAND2_X1 U784 ( .A1(n738), .A2(n737), .ZN(G72) );
  XNOR2_X1 U785 ( .A(G125), .B(n739), .ZN(n740) );
  XNOR2_X1 U786 ( .A(n740), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U787 ( .A(G122), .B(KEYINPUT126), .ZN(n741) );
  XOR2_X1 U788 ( .A(n742), .B(G119), .Z(G21) );
  XNOR2_X1 U789 ( .A(G131), .B(KEYINPUT127), .ZN(n744) );
  XNOR2_X1 U790 ( .A(n744), .B(n743), .ZN(G33) );
  XOR2_X1 U791 ( .A(n745), .B(G137), .Z(G39) );
endmodule

