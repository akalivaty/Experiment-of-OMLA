//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1232, new_n1233, new_n1234, new_n1235, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1293,
    new_n1294, new_n1295;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT64), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G107), .ZN(new_n223));
  INV_X1    g0023(.A(G264), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n202), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n210), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n208), .ZN(new_n230));
  OAI21_X1  g0030(.A(G50), .B1(G58), .B2(G68), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI22_X1  g0032(.A1(new_n226), .A2(KEYINPUT1), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  AND3_X1   g0033(.A1(new_n214), .A2(new_n228), .A3(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  AOI21_X1  g0049(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n250));
  INV_X1    g0050(.A(G274), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n252));
  NOR3_X1   g0052(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G41), .ZN(new_n254));
  INV_X1    g0054(.A(G45), .ZN(new_n255));
  AOI21_X1  g0055(.A(G1), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n250), .A2(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(new_n257), .A2(G226), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT3), .B(G33), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G223), .A3(G1698), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G222), .ZN(new_n263));
  OAI221_X1 g0063(.A(new_n260), .B1(new_n202), .B2(new_n259), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  AOI211_X1 g0064(.A(new_n253), .B(new_n258), .C1(new_n264), .C2(new_n250), .ZN(new_n265));
  INV_X1    g0065(.A(G179), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G13), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n268), .A2(new_n208), .A3(G1), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n229), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n207), .A2(G20), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n272), .A2(G50), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n269), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G150), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n277), .B1(new_n201), .B2(new_n208), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n208), .A2(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT66), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT66), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(new_n208), .A3(G33), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT8), .B(G58), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n278), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n271), .ZN(new_n287));
  OAI221_X1 g0087(.A(new_n274), .B1(G50), .B2(new_n275), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n288), .B1(new_n265), .B2(G169), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n267), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n288), .B(KEYINPUT9), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n265), .A2(G190), .ZN(new_n292));
  INV_X1    g0092(.A(G200), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n291), .B(new_n292), .C1(new_n293), .C2(new_n265), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(KEYINPUT10), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT67), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(KEYINPUT10), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT68), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n297), .B(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n290), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n259), .A2(G226), .A3(new_n261), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n259), .A2(G232), .A3(G1698), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G97), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n250), .ZN(new_n306));
  INV_X1    g0106(.A(G33), .ZN(new_n307));
  OAI211_X1 g0107(.A(G1), .B(G13), .C1(new_n307), .C2(new_n254), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n308), .A2(G274), .A3(new_n256), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n252), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n309), .B1(new_n310), .B2(new_n217), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT13), .ZN(new_n313));
  AND3_X1   g0113(.A1(new_n306), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n313), .B1(new_n306), .B2(new_n312), .ZN(new_n315));
  OAI21_X1  g0115(.A(G169), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT14), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(KEYINPUT69), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT69), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n311), .B1(new_n250), .B2(new_n305), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(new_n320), .B2(new_n313), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n313), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n318), .A2(G179), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n317), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT72), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n316), .B2(KEYINPUT14), .ZN(new_n326));
  INV_X1    g0126(.A(new_n315), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n322), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT14), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n328), .A2(KEYINPUT72), .A3(new_n329), .A4(G169), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n324), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n272), .A2(G68), .A3(new_n273), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n207), .A2(new_n216), .A3(G13), .A4(G20), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n334), .B(KEYINPUT12), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(KEYINPUT70), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT70), .B1(new_n333), .B2(new_n335), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT11), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n280), .A2(G77), .A3(new_n282), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n276), .A2(G50), .B1(G20), .B2(new_n216), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n339), .B1(new_n342), .B2(new_n271), .ZN(new_n343));
  AOI211_X1 g0143(.A(KEYINPUT11), .B(new_n287), .C1(new_n340), .C2(new_n341), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n337), .A2(new_n338), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT71), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI221_X1 g0147(.A(KEYINPUT71), .B1(new_n343), .B2(new_n344), .C1(new_n337), .C2(new_n338), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n332), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n328), .A2(G200), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n318), .A2(G190), .A3(new_n321), .A4(new_n322), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n349), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n259), .A2(G223), .A3(new_n261), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n307), .A2(KEYINPUT3), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT3), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G33), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n357), .A2(new_n359), .A3(G226), .A4(G1698), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G33), .A2(G87), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n356), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n250), .ZN(new_n363));
  INV_X1    g0163(.A(G232), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n309), .B1(new_n310), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n363), .A2(new_n366), .A3(G179), .ZN(new_n367));
  INV_X1    g0167(.A(G169), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n363), .B2(new_n366), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT16), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT7), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(new_n259), .B2(G20), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n357), .A2(new_n359), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n374), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n216), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G58), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n377), .A2(new_n216), .ZN(new_n378));
  NOR2_X1   g0178(.A1(G58), .A2(G68), .ZN(new_n379));
  OAI21_X1  g0179(.A(G20), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n276), .A2(G159), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n371), .B1(new_n376), .B2(new_n382), .ZN(new_n383));
  NOR4_X1   g0183(.A1(new_n259), .A2(KEYINPUT74), .A3(new_n372), .A4(G20), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT74), .ZN(new_n385));
  AOI21_X1  g0185(.A(G20), .B1(new_n357), .B2(new_n359), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n385), .B1(new_n386), .B2(KEYINPUT7), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT73), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n374), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n357), .A2(new_n359), .A3(KEYINPUT73), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(new_n208), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n372), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n216), .B1(new_n388), .B2(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n382), .A2(new_n371), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n271), .B(new_n383), .C1(new_n394), .C2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n272), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n285), .A2(new_n273), .ZN(new_n399));
  OAI22_X1  g0199(.A1(new_n398), .A2(new_n399), .B1(new_n275), .B2(new_n285), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n370), .B1(new_n397), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n402), .B(KEYINPUT18), .ZN(new_n403));
  INV_X1    g0203(.A(G190), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n363), .A2(new_n366), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n365), .B1(new_n250), .B2(new_n362), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n405), .B1(G200), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n388), .A2(new_n393), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n396), .B1(new_n408), .B2(G68), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n383), .A2(new_n271), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n407), .B(new_n401), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  XNOR2_X1  g0211(.A(new_n411), .B(KEYINPUT17), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n403), .A2(new_n412), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n285), .A2(new_n276), .B1(G20), .B2(G77), .ZN(new_n414));
  OR2_X1    g0214(.A1(new_n218), .A2(KEYINPUT15), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n218), .A2(KEYINPUT15), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n414), .B1(new_n279), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n271), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n272), .A2(G77), .A3(new_n273), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n420), .B(new_n421), .C1(G77), .C2(new_n275), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n374), .A2(G107), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n259), .A2(G1698), .ZN(new_n424));
  OAI221_X1 g0224(.A(new_n423), .B1(new_n262), .B2(new_n364), .C1(new_n217), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n250), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n253), .B1(G244), .B2(new_n257), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n422), .B1(new_n429), .B2(G169), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n428), .A2(G179), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n422), .B1(new_n429), .B2(G190), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n428), .A2(G200), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  NOR4_X1   g0237(.A1(new_n301), .A2(new_n355), .A3(new_n413), .A4(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT77), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n259), .A2(new_n208), .A3(G68), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT19), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n208), .B1(new_n304), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(G87), .B2(new_n205), .ZN(new_n443));
  INV_X1    g0243(.A(G97), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n441), .B1(new_n279), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n440), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n446), .A2(new_n271), .B1(new_n269), .B2(new_n418), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n307), .A2(G1), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n269), .A2(new_n271), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G87), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n222), .A2(G1698), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n259), .B(new_n452), .C1(G238), .C2(G1698), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G116), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n250), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n255), .A2(G1), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(new_n219), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n308), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n308), .A2(G274), .ZN(new_n460));
  INV_X1    g0260(.A(new_n457), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n293), .B1(new_n456), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n439), .B1(new_n451), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n308), .B1(new_n453), .B2(new_n454), .ZN(new_n466));
  OAI21_X1  g0266(.A(G200), .B1(new_n466), .B2(new_n462), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n467), .A2(new_n447), .A3(KEYINPUT77), .A4(new_n450), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n466), .A2(new_n462), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G190), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n465), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n449), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT76), .ZN(new_n473));
  XNOR2_X1  g0273(.A(new_n417), .B(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n447), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n469), .A2(new_n266), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n368), .B1(new_n466), .B2(new_n462), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n471), .A2(KEYINPUT78), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT78), .B1(new_n471), .B2(new_n478), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT75), .ZN(new_n483));
  XNOR2_X1  g0283(.A(KEYINPUT5), .B(G41), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n250), .B1(new_n457), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G257), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n484), .A2(new_n308), .A3(G274), .A4(new_n457), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n259), .A2(G244), .A3(new_n261), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n259), .A2(KEYINPUT4), .A3(G244), .A4(new_n261), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n259), .A2(G250), .A3(G1698), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G283), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n491), .A2(new_n492), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n488), .B1(new_n495), .B2(new_n250), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n266), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT6), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n444), .A2(new_n223), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n498), .B1(new_n499), .B2(new_n204), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n223), .A2(KEYINPUT6), .A3(G97), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n502), .A2(G20), .B1(G77), .B2(new_n276), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n259), .A2(new_n372), .A3(G20), .ZN(new_n504));
  AOI21_X1  g0304(.A(KEYINPUT7), .B1(new_n374), .B2(new_n208), .ZN(new_n505));
  OAI21_X1  g0305(.A(G107), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n271), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n275), .A2(G97), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n509), .B1(new_n449), .B2(G97), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n497), .B(new_n511), .C1(G169), .C2(new_n496), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n495), .A2(new_n250), .ZN(new_n513));
  INV_X1    g0313(.A(new_n488), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G200), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n496), .A2(G190), .ZN(new_n517));
  INV_X1    g0317(.A(new_n510), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n518), .B1(new_n507), .B2(new_n271), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n483), .B1(new_n512), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n259), .A2(new_n208), .A3(G87), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT22), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT22), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n259), .A2(new_n524), .A3(new_n208), .A4(G87), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g0326(.A(KEYINPUT80), .B(KEYINPUT24), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n454), .A2(G20), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT23), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n208), .B2(G107), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n223), .A2(KEYINPUT23), .A3(G20), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n526), .A2(new_n527), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n527), .B1(new_n526), .B2(new_n532), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n271), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT25), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n275), .B2(G107), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n269), .A2(KEYINPUT25), .A3(new_n223), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n537), .A2(new_n538), .B1(new_n449), .B2(G107), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n259), .A2(G257), .A3(G1698), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G33), .A2(G294), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n540), .B(new_n541), .C1(new_n262), .C2(new_n219), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n542), .A2(new_n250), .B1(new_n485), .B2(G264), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(G190), .A3(new_n487), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n250), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n485), .A2(G264), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n487), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(G200), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n535), .A2(new_n539), .A3(new_n544), .A4(new_n548), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n535), .A2(new_n539), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n547), .A2(new_n368), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(G179), .B2(new_n547), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n549), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n521), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n484), .A2(new_n457), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n555), .A2(G270), .A3(new_n308), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n487), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n259), .A2(G257), .A3(new_n261), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n374), .A2(G303), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n559), .B(new_n560), .C1(new_n424), .C2(new_n224), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n250), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n449), .A2(G116), .ZN(new_n564));
  INV_X1    g0364(.A(G116), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n269), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n270), .A2(new_n229), .B1(G20), .B2(new_n565), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n494), .B(new_n208), .C1(G33), .C2(new_n444), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT20), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n567), .A2(KEYINPUT20), .A3(new_n568), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n564), .B(new_n566), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n563), .A2(G169), .A3(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT21), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(KEYINPUT79), .A3(new_n573), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n558), .A2(new_n562), .A3(G179), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n571), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n558), .A2(new_n562), .A3(G190), .ZN(new_n577));
  INV_X1    g0377(.A(new_n571), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n557), .B1(new_n250), .B2(new_n561), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n577), .B(new_n578), .C1(new_n579), .C2(new_n293), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n573), .A2(KEYINPUT79), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n563), .A2(G169), .A3(new_n581), .A4(new_n571), .ZN(new_n582));
  AND4_X1   g0382(.A1(new_n574), .A2(new_n576), .A3(new_n580), .A4(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n512), .A2(new_n483), .A3(new_n520), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AND4_X1   g0385(.A1(new_n438), .A2(new_n482), .A3(new_n554), .A4(new_n585), .ZN(G372));
  INV_X1    g0386(.A(new_n403), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n317), .A2(new_n323), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(new_n326), .B2(new_n330), .ZN(new_n589));
  INV_X1    g0389(.A(new_n354), .ZN(new_n590));
  OAI22_X1  g0390(.A1(new_n589), .A2(new_n349), .B1(new_n590), .B2(new_n433), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n587), .B1(new_n591), .B2(new_n412), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(new_n296), .B2(new_n299), .ZN(new_n593));
  OR3_X1    g0393(.A1(new_n593), .A2(KEYINPUT82), .A3(new_n290), .ZN(new_n594));
  OAI21_X1  g0394(.A(KEYINPUT82), .B1(new_n593), .B2(new_n290), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n471), .A2(new_n478), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT78), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n512), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n599), .A2(new_n600), .A3(KEYINPUT26), .A4(new_n479), .ZN(new_n601));
  OR2_X1    g0401(.A1(new_n601), .A2(KEYINPUT81), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT26), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n470), .A2(new_n447), .A3(new_n467), .A4(new_n450), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n478), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n603), .B1(new_n512), .B2(new_n605), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n606), .A2(KEYINPUT81), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n601), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n550), .A2(new_n552), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n574), .A2(new_n576), .A3(new_n582), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n512), .A2(new_n549), .A3(new_n520), .A4(new_n604), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n602), .A2(new_n478), .A3(new_n608), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n438), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n596), .A2(new_n615), .ZN(G369));
  NAND3_X1  g0416(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n617));
  OR2_X1    g0417(.A1(new_n617), .A2(KEYINPUT27), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(KEYINPUT27), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(G213), .A3(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(G343), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n578), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n610), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n583), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n625), .B1(new_n626), .B2(new_n624), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(G330), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n628), .A2(KEYINPUT83), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(KEYINPUT83), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n553), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n550), .B2(new_n623), .ZN(new_n634));
  INV_X1    g0434(.A(new_n609), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n634), .B1(new_n635), .B2(new_n623), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n610), .A2(new_n623), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n633), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n622), .B(KEYINPUT84), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n609), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n638), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g0445(.A(new_n645), .B(KEYINPUT85), .ZN(G399));
  INV_X1    g0446(.A(new_n211), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n647), .A2(G41), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(G1), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n231), .B2(new_n649), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n652), .B(KEYINPUT28), .ZN(new_n653));
  INV_X1    g0453(.A(G330), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n513), .A2(new_n514), .A3(new_n543), .A4(new_n469), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n579), .A2(G179), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT30), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n543), .A2(new_n469), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT30), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n658), .A2(new_n575), .A3(new_n659), .A4(new_n496), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n579), .A2(G179), .A3(new_n469), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n662), .A2(new_n515), .A3(new_n547), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT31), .B1(new_n664), .B2(new_n622), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT31), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n642), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n665), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n482), .A2(new_n585), .A3(new_n554), .A4(new_n642), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n654), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT29), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT86), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n614), .A2(new_n672), .A3(new_n642), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n672), .B1(new_n614), .B2(new_n642), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n671), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n478), .B1(new_n611), .B2(new_n612), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n512), .A2(new_n605), .A3(new_n603), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT87), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n599), .A2(new_n479), .A3(new_n600), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n603), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n676), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n622), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(KEYINPUT29), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n670), .B1(new_n675), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n653), .B1(new_n685), .B2(G1), .ZN(G364));
  NOR2_X1   g0486(.A1(new_n268), .A2(G20), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n207), .B1(new_n687), .B2(G45), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n648), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OAI211_X1 g0491(.A(new_n631), .B(new_n691), .C1(G330), .C2(new_n627), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n647), .A2(new_n374), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G355), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(G116), .B2(new_n211), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n357), .A2(new_n359), .A3(KEYINPUT73), .ZN(new_n696));
  AOI21_X1  g0496(.A(KEYINPUT73), .B1(new_n357), .B2(new_n359), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(new_n647), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n701), .B1(new_n255), .B2(new_n232), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n245), .A2(new_n255), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n695), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(G13), .A2(G33), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G20), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n229), .B1(G20), .B2(new_n368), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n690), .B1(new_n704), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n208), .A2(G179), .ZN(new_n712));
  NOR2_X1   g0512(.A1(G190), .A2(G200), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n714), .A2(KEYINPUT89), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(KEYINPUT89), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G329), .ZN(new_n719));
  INV_X1    g0519(.A(G283), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n712), .A2(new_n404), .A3(G200), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n712), .A2(G190), .A3(G200), .ZN(new_n722));
  INV_X1    g0522(.A(G303), .ZN(new_n723));
  OAI22_X1  g0523(.A1(new_n720), .A2(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n208), .A2(new_n266), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G200), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G190), .ZN(new_n727));
  XNOR2_X1  g0527(.A(KEYINPUT33), .B(G317), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n724), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n725), .A2(new_n713), .ZN(new_n730));
  INV_X1    g0530(.A(G311), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n374), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n725), .A2(G190), .A3(new_n293), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n732), .B1(G322), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n726), .A2(new_n404), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n266), .A2(new_n293), .A3(G190), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  AOI22_X1  g0538(.A1(new_n736), .A2(G326), .B1(G294), .B2(new_n738), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n719), .A2(new_n729), .A3(new_n735), .A4(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G159), .ZN(new_n741));
  OR3_X1    g0541(.A1(new_n717), .A2(KEYINPUT32), .A3(new_n741), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n738), .B(KEYINPUT90), .Z(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G97), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n722), .A2(new_n218), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n721), .A2(new_n223), .ZN(new_n746));
  AOI211_X1 g0546(.A(new_n745), .B(new_n746), .C1(G68), .C2(new_n727), .ZN(new_n747));
  OAI21_X1  g0547(.A(KEYINPUT32), .B1(new_n717), .B2(new_n741), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n742), .A2(new_n744), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n733), .A2(new_n377), .B1(new_n730), .B2(new_n202), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n750), .A2(KEYINPUT88), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(KEYINPUT88), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n374), .B1(new_n736), .B2(G50), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n751), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n740), .B1(new_n749), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT91), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n708), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(new_n755), .B2(new_n756), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n711), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n707), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n760), .B1(new_n627), .B2(new_n761), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n692), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(G396));
  NOR2_X1   g0564(.A1(new_n708), .A2(new_n705), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n730), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n734), .A2(G143), .B1(new_n767), .B2(G159), .ZN(new_n768));
  INV_X1    g0568(.A(new_n727), .ZN(new_n769));
  INV_X1    g0569(.A(G150), .ZN(new_n770));
  INV_X1    g0570(.A(G137), .ZN(new_n771));
  INV_X1    g0571(.A(new_n736), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n768), .B1(new_n769), .B2(new_n770), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT34), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n721), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n698), .B1(G68), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n722), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n778), .A2(G50), .B1(new_n738), .B2(G58), .ZN(new_n779));
  INV_X1    g0579(.A(G132), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n777), .B(new_n779), .C1(new_n780), .C2(new_n717), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n775), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n773), .A2(new_n774), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n769), .A2(new_n720), .B1(new_n721), .B2(new_n218), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n717), .A2(new_n731), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n772), .A2(new_n723), .B1(new_n722), .B2(new_n223), .ZN(new_n786));
  INV_X1    g0586(.A(G294), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n374), .B1(new_n730), .B2(new_n565), .C1(new_n787), .C2(new_n733), .ZN(new_n788));
  NOR4_X1   g0588(.A1(new_n784), .A2(new_n785), .A3(new_n786), .A4(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n782), .A2(new_n783), .B1(new_n789), .B2(new_n744), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n690), .B1(G77), .B2(new_n766), .C1(new_n790), .C2(new_n758), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT92), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n432), .A2(new_n623), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n422), .A2(new_n622), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n436), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n793), .B1(new_n795), .B2(new_n432), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n792), .B1(new_n706), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n796), .B1(new_n673), .B2(new_n674), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n614), .A2(new_n642), .A3(new_n797), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n670), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(KEYINPUT93), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n690), .B1(new_n801), .B2(new_n670), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n802), .A2(KEYINPUT93), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n798), .B1(new_n805), .B2(new_n806), .ZN(G384));
  OR2_X1    g0607(.A1(new_n502), .A2(KEYINPUT35), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n502), .A2(KEYINPUT35), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n808), .A2(G116), .A3(new_n230), .A4(new_n809), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT36), .Z(new_n811));
  OAI211_X1 g0611(.A(new_n232), .B(G77), .C1(new_n377), .C2(new_n216), .ZN(new_n812));
  INV_X1    g0612(.A(G50), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G68), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n207), .B(G13), .C1(new_n812), .C2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n675), .A2(new_n438), .A3(new_n684), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n596), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT99), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n350), .A2(new_n622), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n354), .B(new_n820), .C1(new_n589), .C2(new_n349), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n350), .B(new_n622), .C1(new_n332), .C2(new_n590), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(new_n800), .B2(new_n793), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT38), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT94), .ZN(new_n827));
  AOI21_X1  g0627(.A(KEYINPUT7), .B1(new_n698), .B2(new_n208), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n375), .A2(KEYINPUT74), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n386), .A2(new_n385), .A3(KEYINPUT7), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(G68), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n395), .ZN(new_n833));
  OAI21_X1  g0633(.A(G68), .B1(new_n504), .B2(new_n505), .ZN(new_n834));
  INV_X1    g0634(.A(new_n382), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n287), .B1(new_n836), .B2(new_n371), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n400), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n411), .B1(new_n838), .B2(new_n370), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT37), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n838), .B2(new_n620), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n827), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n401), .B1(new_n409), .B2(new_n410), .ZN(new_n843));
  INV_X1    g0643(.A(new_n620), .ZN(new_n844));
  AOI21_X1  g0644(.A(KEYINPUT37), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n370), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n845), .A2(KEYINPUT94), .A3(new_n847), .A4(new_n411), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n842), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n287), .B1(new_n832), .B2(new_n395), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n371), .B1(new_n394), .B2(new_n382), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n400), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n411), .B1(new_n852), .B2(new_n620), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n852), .A2(new_n370), .ZN(new_n854));
  OAI21_X1  g0654(.A(KEYINPUT37), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n849), .A2(KEYINPUT95), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT16), .B1(new_n832), .B2(new_n835), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n271), .B1(new_n394), .B2(new_n396), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n401), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n844), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n413), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n856), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT95), .B1(new_n849), .B2(new_n855), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n826), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n849), .A2(new_n855), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT95), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n868), .A2(KEYINPUT38), .A3(new_n862), .A4(new_n856), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n865), .A2(KEYINPUT96), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT96), .B1(new_n865), .B2(new_n869), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n825), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT39), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n860), .B1(new_n403), .B2(new_n412), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n859), .A2(new_n846), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n875), .A2(new_n860), .A3(new_n411), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n842), .A2(new_n848), .B1(new_n876), .B2(KEYINPUT37), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n874), .B1(new_n877), .B2(KEYINPUT95), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT97), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n878), .A2(new_n879), .A3(KEYINPUT38), .A4(new_n868), .ZN(new_n880));
  NOR3_X1   g0680(.A1(new_n863), .A2(new_n826), .A3(new_n864), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n838), .A2(new_n620), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT37), .B1(new_n839), .B2(new_n882), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n413), .A2(new_n882), .B1(new_n849), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT97), .B1(new_n884), .B2(KEYINPUT38), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n873), .B(new_n880), .C1(new_n881), .C2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n351), .A2(new_n622), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n865), .A2(KEYINPUT39), .A3(new_n869), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n587), .A2(new_n620), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n872), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT98), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT98), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n872), .A2(new_n889), .A3(new_n893), .A4(new_n890), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n819), .B(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n796), .B1(new_n821), .B2(new_n822), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n666), .B(new_n623), .C1(new_n661), .C2(new_n663), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n665), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n669), .A2(new_n899), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n897), .A2(new_n900), .A3(KEYINPUT40), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n901), .B(new_n880), .C1(new_n881), .C2(new_n885), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT100), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n902), .B(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n897), .A2(new_n900), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT96), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT38), .B1(new_n878), .B2(new_n868), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n906), .B1(new_n881), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n865), .A2(KEYINPUT96), .A3(new_n869), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n904), .B1(KEYINPUT40), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n438), .A2(new_n900), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n912), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n913), .A2(G330), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n896), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n207), .B2(new_n687), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n896), .A2(new_n915), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n816), .B1(new_n917), .B2(new_n918), .ZN(G367));
  NAND2_X1  g0719(.A1(new_n700), .A2(new_n241), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n710), .B1(new_n647), .B2(new_n417), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n691), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n451), .A2(new_n622), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n478), .A2(new_n923), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n924), .A2(KEYINPUT101), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n604), .A2(new_n478), .A3(new_n923), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(KEYINPUT101), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n721), .A2(new_n444), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n738), .A2(G107), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n772), .B2(new_n731), .ZN(new_n931));
  AOI211_X1 g0731(.A(new_n929), .B(new_n931), .C1(G294), .C2(new_n727), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n733), .A2(new_n723), .B1(new_n730), .B2(new_n720), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n699), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n718), .A2(G317), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n778), .A2(G116), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT46), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n932), .A2(new_n934), .A3(new_n935), .A4(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n743), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n939), .A2(new_n216), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n769), .A2(new_n741), .B1(new_n722), .B2(new_n377), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n717), .A2(new_n771), .ZN(new_n942));
  INV_X1    g0742(.A(G143), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n772), .A2(new_n943), .B1(new_n721), .B2(new_n202), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n259), .B1(new_n730), .B2(new_n813), .C1(new_n770), .C2(new_n733), .ZN(new_n945));
  OR4_X1    g0745(.A1(new_n941), .A2(new_n942), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n938), .B1(new_n940), .B2(new_n946), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n947), .B(KEYINPUT47), .Z(new_n948));
  OAI221_X1 g0748(.A(new_n922), .B1(new_n761), .B2(new_n928), .C1(new_n948), .C2(new_n758), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n648), .B(KEYINPUT41), .Z(new_n950));
  NAND2_X1  g0750(.A1(new_n600), .A2(new_n641), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n512), .B(new_n520), .C1(new_n519), .C2(new_n642), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n644), .A2(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT44), .Z(new_n955));
  NOR2_X1   g0755(.A1(new_n644), .A2(new_n953), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT45), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(new_n638), .B2(KEYINPUT106), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT106), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n637), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n958), .A2(new_n960), .A3(new_n637), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n640), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(KEYINPUT104), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n636), .A2(new_n639), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n965), .A2(KEYINPUT104), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n632), .B2(KEYINPUT105), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n632), .A2(KEYINPUT105), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n970), .B(new_n971), .Z(new_n972));
  NAND3_X1  g0772(.A1(new_n964), .A2(new_n685), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n950), .B1(new_n973), .B2(new_n685), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(new_n689), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n953), .A2(new_n640), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT42), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n512), .B1(new_n635), .B2(new_n952), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n642), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT102), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n928), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT103), .Z(new_n986));
  AND2_X1   g0786(.A1(new_n928), .A2(KEYINPUT43), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n986), .B1(new_n980), .B2(new_n988), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n637), .A2(new_n953), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n989), .B(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n949), .B1(new_n975), .B2(new_n991), .ZN(G387));
  INV_X1    g0792(.A(new_n650), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n693), .A2(new_n993), .B1(new_n223), .B2(new_n647), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n238), .A2(new_n255), .ZN(new_n995));
  AOI21_X1  g0795(.A(G45), .B1(G68), .B2(G77), .ZN(new_n996));
  AND3_X1   g0796(.A1(new_n285), .A2(KEYINPUT50), .A3(new_n813), .ZN(new_n997));
  AOI21_X1  g0797(.A(KEYINPUT50), .B1(new_n285), .B2(new_n813), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n650), .B(new_n996), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n700), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n994), .B1(new_n995), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n709), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n690), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n636), .A2(new_n761), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n741), .A2(new_n772), .B1(new_n769), .B2(new_n284), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n929), .B(new_n1005), .C1(G77), .C2(new_n778), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n474), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n743), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n718), .A2(G150), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n733), .A2(new_n813), .B1(new_n730), .B2(new_n216), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1010), .A2(new_n698), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1006), .A2(new_n1008), .A3(new_n1009), .A4(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n734), .A2(G317), .B1(new_n767), .B2(G303), .ZN(new_n1013));
  INV_X1    g0813(.A(G322), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1013), .B1(new_n769), .B2(new_n731), .C1(new_n1014), .C2(new_n772), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT48), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n778), .A2(G294), .B1(new_n738), .B2(G283), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT49), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1022), .A2(KEYINPUT107), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n698), .B1(new_n565), .B2(new_n721), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(new_n718), .B2(G326), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT107), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1025), .B1(new_n1021), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1012), .B1(new_n1023), .B2(new_n1027), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1003), .B(new_n1004), .C1(new_n708), .C2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n972), .B2(new_n689), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n972), .A2(new_n685), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n648), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n972), .A2(new_n685), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1030), .B1(new_n1032), .B2(new_n1033), .ZN(G393));
  NAND3_X1  g0834(.A1(new_n1031), .A2(new_n963), .A3(new_n962), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1035), .A2(new_n648), .A3(new_n973), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n953), .A2(new_n707), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n709), .B1(new_n444), .B2(new_n211), .C1(new_n701), .C2(new_n248), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT108), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1040), .A2(new_n690), .A3(new_n1041), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n699), .B1(new_n284), .B2(new_n730), .C1(new_n717), .C2(new_n943), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n722), .A2(new_n216), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n769), .A2(new_n813), .B1(new_n721), .B2(new_n218), .ZN(new_n1045));
  NOR3_X1   g0845(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n772), .A2(new_n770), .B1(new_n741), .B2(new_n733), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT51), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n743), .A2(G77), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1046), .A2(new_n1049), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n259), .B(new_n746), .C1(G283), .C2(new_n778), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n1014), .B2(new_n717), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT109), .Z(new_n1055));
  AOI22_X1  g0855(.A1(new_n767), .A2(G294), .B1(G116), .B2(new_n738), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n723), .B2(new_n769), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT110), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G317), .A2(new_n736), .B1(new_n734), .B2(G311), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT52), .Z(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1052), .B1(new_n1055), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1042), .B1(new_n1062), .B2(new_n708), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n964), .A2(new_n689), .B1(new_n1037), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1036), .A2(new_n1064), .ZN(G390));
  XNOR2_X1  g0865(.A(KEYINPUT54), .B(G143), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n727), .A2(G137), .B1(new_n767), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT114), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n743), .A2(G159), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n1069), .B2(new_n1068), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT115), .ZN(new_n1072));
  OAI21_X1  g0872(.A(KEYINPUT53), .B1(new_n722), .B2(new_n770), .ZN(new_n1073));
  OR3_X1    g0873(.A1(new_n722), .A2(KEYINPUT53), .A3(new_n770), .ZN(new_n1074));
  INV_X1    g0874(.A(G125), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1073), .B(new_n1074), .C1(new_n717), .C2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(G128), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n259), .B1(new_n780), .B2(new_n733), .C1(new_n772), .C2(new_n1077), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1076), .B(new_n1078), .C1(G50), .C2(new_n776), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1072), .A2(new_n1079), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n223), .A2(new_n769), .B1(new_n772), .B2(new_n720), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n745), .B(new_n1081), .C1(G68), .C2(new_n776), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n718), .A2(G294), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n374), .B1(new_n733), .B2(new_n565), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G97), .B2(new_n767), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1082), .A2(new_n1050), .A3(new_n1083), .A4(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n758), .B1(new_n1080), .B2(new_n1086), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n691), .B(new_n1087), .C1(new_n284), .C2(new_n765), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n886), .A2(new_n888), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1088), .B1(new_n1090), .B2(new_n706), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1089), .B1(new_n825), .B2(new_n887), .ZN(new_n1092));
  OR2_X1    g0892(.A1(new_n682), .A2(new_n622), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n795), .A2(new_n432), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n793), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n823), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n887), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n881), .A2(new_n885), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .A4(new_n880), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n654), .B1(new_n669), .B2(new_n899), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n897), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1101), .A2(KEYINPUT111), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n670), .A2(new_n797), .A3(new_n823), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  AND3_X1   g0905(.A1(new_n1092), .A2(new_n1099), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1101), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1092), .A2(new_n1099), .B1(KEYINPUT111), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1091), .B1(new_n1109), .B2(new_n688), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n438), .A2(new_n1100), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n817), .A2(new_n596), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n670), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n824), .B1(new_n1113), .B2(new_n796), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1114), .A2(new_n1101), .B1(new_n793), .B2(new_n800), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1100), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n824), .B1(new_n1116), .B2(new_n796), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n1103), .ZN(new_n1118));
  OAI21_X1  g0918(.A(KEYINPUT112), .B1(new_n1118), .B2(new_n1095), .ZN(new_n1119));
  NOR3_X1   g0919(.A1(new_n682), .A2(new_n622), .A3(new_n1094), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n793), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT112), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1122), .A2(new_n1123), .A3(new_n1117), .A4(new_n1103), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1115), .B1(new_n1119), .B2(new_n1124), .ZN(new_n1125));
  OR2_X1    g0925(.A1(new_n1112), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1109), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1112), .A2(new_n1125), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1127), .A2(new_n648), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(KEYINPUT113), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT113), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1127), .A2(new_n1132), .A3(new_n648), .A4(new_n1129), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1110), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(G378));
  OAI21_X1  g0935(.A(G330), .B1(new_n910), .B2(KEYINPUT40), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n902), .B(KEYINPUT100), .ZN(new_n1137));
  XOR2_X1   g0937(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n288), .A2(new_n844), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT116), .Z(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n300), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n300), .A2(new_n1142), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1139), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1145), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1147), .A2(new_n1138), .A3(new_n1143), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NOR3_X1   g0949(.A1(new_n1136), .A2(new_n1137), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1149), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n905), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n870), .B2(new_n871), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT40), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n654), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1151), .B1(new_n1155), .B2(new_n904), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n894), .B(new_n892), .C1(new_n1150), .C2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT118), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n892), .A2(new_n894), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1155), .A2(new_n904), .A3(new_n1151), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1149), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1157), .A2(new_n1158), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1159), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(KEYINPUT118), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1163), .A2(new_n1165), .A3(new_n689), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n733), .A2(new_n1077), .B1(new_n730), .B2(new_n771), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G132), .B2(new_n727), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n736), .A2(G125), .B1(new_n778), .B2(new_n1067), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1168), .B(new_n1169), .C1(new_n939), .C2(new_n770), .ZN(new_n1170));
  OR2_X1    g0970(.A1(new_n1170), .A2(KEYINPUT59), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(KEYINPUT59), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n307), .B(new_n254), .C1(new_n721), .C2(new_n741), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n718), .B2(G124), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1171), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  AOI211_X1 g0975(.A(G41), .B(new_n699), .C1(G107), .C2(new_n734), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1176), .B1(new_n720), .B2(new_n717), .C1(new_n474), .C2(new_n730), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n377), .A2(new_n721), .B1(new_n722), .B2(new_n202), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n444), .A2(new_n769), .B1(new_n772), .B2(new_n565), .ZN(new_n1179));
  NOR4_X1   g0979(.A1(new_n1177), .A2(new_n940), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1180), .A2(KEYINPUT58), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(KEYINPUT58), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n254), .B1(new_n698), .B2(new_n307), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n813), .ZN(new_n1184));
  AND4_X1   g0984(.A1(new_n1175), .A2(new_n1181), .A3(new_n1182), .A4(new_n1184), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n690), .B1(G50), .B2(new_n766), .C1(new_n1185), .C2(new_n758), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n1149), .B2(new_n705), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT117), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1166), .A2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1112), .B(KEYINPUT119), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1129), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1162), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1192), .B(KEYINPUT57), .C1(new_n1193), .C2(new_n1164), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n648), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1163), .A2(new_n1165), .A3(new_n1192), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT57), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT120), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1195), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1196), .A2(KEYINPUT120), .A3(new_n1197), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1190), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(G375));
  OAI21_X1  g1003(.A(new_n690), .B1(G68), .B2(new_n766), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n1204), .B(KEYINPUT121), .Z(new_n1205));
  AOI22_X1  g1005(.A1(new_n727), .A2(G116), .B1(new_n736), .B2(G294), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n734), .A2(G283), .B1(new_n767), .B2(G107), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(new_n444), .C2(new_n722), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G303), .B2(new_n718), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n374), .B1(new_n721), .B2(new_n202), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT122), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1209), .A2(new_n1008), .A3(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT123), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n769), .A2(new_n1066), .B1(new_n721), .B2(new_n377), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n772), .A2(new_n780), .B1(new_n722), .B2(new_n741), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n743), .A2(G50), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n718), .A2(G128), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n733), .A2(new_n771), .B1(new_n730), .B2(new_n770), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1220), .A2(new_n698), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .A4(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1214), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1205), .B1(new_n758), .B2(new_n1224), .C1(new_n823), .C2(new_n706), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n1125), .B2(new_n688), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1128), .A2(new_n950), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1112), .A2(new_n1125), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1227), .B1(new_n1228), .B2(new_n1230), .ZN(G381));
  OR4_X1    g1031(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1110), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1130), .A2(new_n1233), .ZN(new_n1234));
  NOR4_X1   g1034(.A1(new_n1232), .A2(G387), .A3(G381), .A4(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n1202), .ZN(G407));
  INV_X1    g1036(.A(new_n1234), .ZN(new_n1237));
  INV_X1    g1037(.A(G213), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1238), .A2(G343), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1202), .A2(new_n1237), .A3(new_n1239), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT124), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1241), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1042(.A(new_n1239), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1112), .A2(new_n1125), .A3(KEYINPUT60), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n648), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1126), .A2(KEYINPUT60), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1245), .B1(new_n1246), .B2(new_n1229), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1247), .A2(new_n1226), .ZN(new_n1248));
  OR2_X1    g1048(.A1(new_n1248), .A2(G384), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(G384), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n1134), .B(new_n1190), .C1(new_n1200), .C2(new_n1201), .ZN(new_n1252));
  OR2_X1    g1052(.A1(new_n1196), .A2(new_n950), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1157), .A2(new_n1162), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1188), .B1(new_n1254), .B2(new_n689), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1234), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1243), .B(new_n1251), .C1(new_n1252), .C2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(KEYINPUT62), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT61), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1256), .B1(new_n1202), .B2(G378), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT125), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1249), .A2(new_n1261), .A3(new_n1250), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1239), .A2(G2897), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1261), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n1260), .A2(new_n1239), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1269), .A2(new_n648), .A3(new_n1201), .A4(new_n1194), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1190), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1270), .A2(G378), .A3(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1256), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT62), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1274), .A2(new_n1275), .A3(new_n1243), .A4(new_n1251), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1258), .A2(new_n1259), .A3(new_n1268), .A4(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(G390), .ZN(new_n1278));
  AND2_X1   g1078(.A1(G387), .A2(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(G387), .A2(new_n1278), .ZN(new_n1280));
  OAI21_X1  g1080(.A(KEYINPUT126), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(G393), .B(new_n763), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1282), .ZN(new_n1284));
  OAI211_X1 g1084(.A(KEYINPUT126), .B(new_n1284), .C1(new_n1279), .C2(new_n1280), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1277), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT63), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1286), .B1(new_n1257), .B2(new_n1288), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1274), .A2(KEYINPUT63), .A3(new_n1243), .A4(new_n1251), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1289), .A2(new_n1259), .A3(new_n1290), .A4(new_n1268), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1287), .A2(new_n1291), .ZN(G405));
  NAND2_X1  g1092(.A1(new_n1251), .A2(KEYINPUT127), .ZN(new_n1293));
  XNOR2_X1  g1093(.A(new_n1286), .B(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1252), .B1(G375), .B2(new_n1237), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1294), .B(new_n1295), .ZN(G402));
endmodule


