//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 1 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G221), .ZN(new_n188));
  INV_X1    g002(.A(G234), .ZN(new_n189));
  NOR3_X1   g003(.A1(new_n188), .A2(new_n189), .A3(G953), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n187), .B(new_n190), .Z(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT78), .ZN(new_n193));
  AND3_X1   g007(.A1(KEYINPUT77), .A2(G125), .A3(G140), .ZN(new_n194));
  AOI21_X1  g008(.A(G140), .B1(KEYINPUT77), .B2(G125), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n193), .B(KEYINPUT16), .C1(new_n194), .C2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT16), .ZN(new_n197));
  NAND2_X1  g011(.A1(KEYINPUT77), .A2(G125), .ZN(new_n198));
  INV_X1    g012(.A(G140), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(KEYINPUT77), .A2(G125), .A3(G140), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n197), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(G125), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT78), .B1(new_n203), .B2(KEYINPUT16), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n196), .B1(new_n202), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G146), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  INV_X1    g021(.A(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G140), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT80), .ZN(new_n210));
  AND3_X1   g024(.A1(new_n203), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n210), .B1(new_n203), .B2(new_n209), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n207), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n206), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT79), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT24), .B(G110), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT76), .ZN(new_n218));
  INV_X1    g032(.A(G119), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G128), .ZN(new_n220));
  INV_X1    g034(.A(G128), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G119), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n218), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n220), .A2(new_n222), .A3(new_n218), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n217), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n221), .A2(KEYINPUT23), .A3(G119), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n219), .A2(G128), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n220), .B(new_n227), .C1(new_n228), .C2(KEYINPUT23), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(G110), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n215), .B1(new_n226), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n230), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n220), .A2(new_n222), .A3(new_n218), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n216), .B1(new_n233), .B2(new_n223), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n232), .A2(KEYINPUT79), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n214), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n224), .A2(new_n225), .A3(new_n217), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n229), .A2(G110), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n196), .B(new_n207), .C1(new_n202), .C2(new_n204), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n239), .B1(new_n240), .B2(new_n206), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n192), .B1(new_n236), .B2(new_n241), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n206), .A2(new_n213), .ZN(new_n243));
  NOR3_X1   g057(.A1(new_n226), .A2(new_n230), .A3(new_n215), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT79), .B1(new_n232), .B2(new_n234), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n206), .A2(new_n240), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(new_n237), .A3(new_n238), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n246), .A2(new_n248), .A3(new_n191), .ZN(new_n249));
  INV_X1    g063(.A(G902), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n242), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT81), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT25), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n251), .A2(KEYINPUT81), .A3(KEYINPUT25), .ZN(new_n255));
  OAI21_X1  g069(.A(G217), .B1(new_n189), .B2(G902), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n256), .B(KEYINPUT75), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n254), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n242), .A2(new_n249), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n257), .A2(G902), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n219), .A2(G116), .ZN(new_n264));
  INV_X1    g078(.A(G116), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G119), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT2), .B(G113), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n264), .A2(new_n266), .A3(KEYINPUT72), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  OR2_X1    g086(.A1(new_n267), .A2(new_n270), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n207), .A2(G143), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT64), .ZN(new_n277));
  NOR3_X1   g091(.A1(new_n277), .A2(new_n207), .A3(G143), .ZN(new_n278));
  INV_X1    g092(.A(G143), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT64), .B1(new_n279), .B2(G146), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n276), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  AND2_X1   g095(.A1(KEYINPUT0), .A2(G128), .ZN(new_n282));
  NOR2_X1   g096(.A1(KEYINPUT0), .A2(G128), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n279), .A2(G146), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT65), .B1(new_n207), .B2(G143), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT65), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(new_n279), .A3(G146), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n285), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n281), .A2(new_n284), .B1(new_n289), .B2(new_n282), .ZN(new_n290));
  XNOR2_X1  g104(.A(KEYINPUT67), .B(G137), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT11), .ZN(new_n292));
  INV_X1    g106(.A(G134), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n291), .A2(new_n294), .B1(new_n293), .B2(G137), .ZN(new_n295));
  INV_X1    g109(.A(G131), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n292), .B1(new_n293), .B2(G137), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT66), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT66), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n299), .B(new_n292), .C1(new_n293), .C2(G137), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n295), .A2(new_n296), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n296), .B1(new_n295), .B2(new_n301), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n290), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n295), .A2(new_n301), .A3(new_n296), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT69), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT68), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n307), .B1(new_n293), .B2(G137), .ZN(new_n308));
  INV_X1    g122(.A(G137), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(KEYINPUT68), .A3(G134), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n308), .B(new_n310), .C1(new_n291), .C2(G134), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n306), .B1(new_n311), .B2(G131), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n309), .A2(KEYINPUT67), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT67), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G137), .ZN(new_n315));
  AOI21_X1  g129(.A(G134), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n308), .A2(new_n310), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n306), .B(G131), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n305), .B1(new_n312), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT71), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n287), .B1(new_n279), .B2(G146), .ZN(new_n322));
  NOR3_X1   g136(.A1(new_n207), .A2(KEYINPUT65), .A3(G143), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n276), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AND2_X1   g138(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n325));
  NOR2_X1   g139(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G128), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n321), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  NOR3_X1   g143(.A1(new_n325), .A2(new_n326), .A3(new_n221), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n289), .A2(KEYINPUT71), .A3(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(G128), .B1(new_n327), .B2(new_n285), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n329), .A2(new_n331), .B1(new_n281), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n304), .B1(new_n320), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT30), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n332), .A2(new_n281), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n289), .A2(KEYINPUT71), .A3(new_n330), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT71), .B1(new_n289), .B2(new_n330), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(G131), .B1(new_n316), .B2(new_n317), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT69), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n318), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n339), .A2(new_n342), .A3(new_n305), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT30), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n344), .A3(new_n304), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n275), .B1(new_n335), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n275), .A3(new_n304), .ZN(new_n347));
  NOR2_X1   g161(.A1(G237), .A2(G953), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G210), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n349), .B(KEYINPUT27), .ZN(new_n350));
  XNOR2_X1  g164(.A(KEYINPUT26), .B(G101), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n350), .B(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT31), .B1(new_n346), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT28), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n347), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n334), .A2(new_n274), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n343), .A2(KEYINPUT28), .A3(new_n275), .A4(new_n304), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n352), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n343), .A2(new_n344), .A3(new_n304), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n344), .B1(new_n343), .B2(new_n304), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n274), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT31), .ZN(new_n365));
  INV_X1    g179(.A(new_n353), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n354), .A2(new_n361), .A3(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(G472), .A2(G902), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n368), .A2(KEYINPUT32), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(KEYINPUT32), .B1(new_n368), .B2(new_n369), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT29), .ZN(new_n373));
  INV_X1    g187(.A(new_n347), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n346), .A2(new_n374), .A3(new_n352), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n275), .B1(new_n343), .B2(new_n304), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n376), .B1(new_n355), .B2(new_n347), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n360), .B1(new_n377), .B2(new_n358), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n373), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n250), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n352), .A2(KEYINPUT29), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT73), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n357), .A2(new_n382), .A3(new_n347), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n334), .A2(KEYINPUT73), .A3(new_n274), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(KEYINPUT28), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT74), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(new_n356), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n383), .A2(KEYINPUT74), .A3(KEYINPUT28), .A4(new_n384), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n381), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(G472), .B1(new_n380), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n263), .B1(new_n372), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT10), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n221), .B1(new_n276), .B2(KEYINPUT1), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n289), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n394), .B1(new_n329), .B2(new_n331), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT83), .ZN(new_n396));
  INV_X1    g210(.A(G107), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n396), .B1(new_n397), .B2(G104), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(G104), .ZN(new_n399));
  INV_X1    g213(.A(G104), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(KEYINPUT83), .A3(G107), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n398), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G101), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n397), .A2(G104), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G101), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n397), .A2(KEYINPUT3), .A3(G104), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT3), .B1(new_n397), .B2(G104), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n405), .B(new_n406), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n392), .B1(new_n395), .B2(new_n410), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n403), .A2(new_n409), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n339), .A2(KEYINPUT10), .A3(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n302), .A2(new_n303), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT3), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n416), .B1(new_n400), .B2(G107), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n397), .A2(KEYINPUT3), .A3(G104), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n404), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n415), .B1(new_n419), .B2(new_n406), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G101), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(new_n415), .A3(G101), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n290), .A3(new_n424), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n411), .A2(new_n413), .A3(new_n414), .A4(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT12), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n289), .A2(new_n393), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n428), .B1(new_n337), .B2(new_n338), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n412), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n336), .B(new_n410), .C1(new_n337), .C2(new_n338), .ZN(new_n431));
  AOI211_X1 g245(.A(new_n427), .B(new_n414), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n431), .B1(new_n395), .B2(new_n410), .ZN(new_n433));
  INV_X1    g247(.A(new_n414), .ZN(new_n434));
  AOI21_X1  g248(.A(KEYINPUT12), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n426), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(G110), .B(G140), .ZN(new_n437));
  INV_X1    g251(.A(G227), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n438), .A2(G953), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n437), .B(new_n439), .ZN(new_n440));
  XOR2_X1   g254(.A(new_n440), .B(KEYINPUT82), .Z(new_n441));
  INV_X1    g255(.A(new_n440), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n426), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n412), .A2(KEYINPUT10), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n425), .B1(new_n333), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT10), .B1(new_n429), .B2(new_n412), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n434), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n436), .A2(new_n441), .B1(new_n443), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(G469), .B1(new_n448), .B2(G902), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT84), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n447), .A2(new_n426), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n440), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n426), .B(new_n442), .C1(new_n432), .C2(new_n435), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G469), .ZN(new_n455));
  AND4_X1   g269(.A1(new_n450), .A2(new_n454), .A3(new_n455), .A4(new_n250), .ZN(new_n456));
  AOI21_X1  g270(.A(G902), .B1(new_n452), .B2(new_n453), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n450), .B1(new_n457), .B2(new_n455), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n449), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT9), .B(G234), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n188), .B1(new_n461), .B2(new_n250), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G237), .ZN(new_n464));
  INV_X1    g278(.A(G953), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n464), .A2(new_n465), .A3(G214), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT90), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n467), .A2(G143), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n348), .B(G214), .C1(new_n467), .C2(G143), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(G131), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT17), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n469), .A2(new_n470), .A3(new_n296), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n296), .B1(new_n469), .B2(new_n470), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT17), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n475), .A2(new_n240), .A3(new_n206), .A4(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT92), .B1(new_n194), .B2(new_n195), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT92), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n200), .A2(new_n480), .A3(new_n201), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n479), .A2(new_n481), .A3(KEYINPUT93), .A4(G146), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT18), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n469), .B(new_n470), .C1(KEYINPUT91), .C2(new_n483), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n483), .A2(KEYINPUT91), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n469), .A2(new_n470), .A3(new_n296), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n486), .B1(new_n487), .B2(new_n476), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT93), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n479), .A2(new_n481), .A3(G146), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n213), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n485), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(G113), .B(G122), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(new_n400), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n478), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n472), .A2(new_n474), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n479), .A2(new_n481), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT19), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n203), .A2(new_n209), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT80), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n203), .A2(new_n209), .A3(new_n210), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT19), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(G146), .B1(new_n498), .B2(new_n503), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n206), .B(new_n496), .C1(new_n504), .C2(KEYINPUT94), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT19), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n502), .B1(new_n479), .B2(new_n481), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n207), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT94), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n492), .B1(new_n505), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n494), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n495), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(G475), .A2(G902), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(KEYINPUT20), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT20), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n504), .A2(KEYINPUT94), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n508), .A2(new_n509), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n518), .A2(new_n519), .A3(new_n206), .A4(new_n496), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n494), .B1(new_n520), .B2(new_n492), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n517), .B(new_n514), .C1(new_n521), .C2(new_n495), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n494), .B1(new_n478), .B2(new_n492), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n250), .B1(new_n495), .B2(new_n524), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n525), .A2(G475), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(G122), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT95), .B1(new_n529), .B2(G116), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT95), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(new_n265), .A3(G122), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n533), .A2(KEYINPUT14), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n533), .A2(KEYINPUT14), .B1(G116), .B2(new_n529), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n397), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n529), .A2(G116), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n533), .A2(new_n397), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(KEYINPUT96), .B1(new_n279), .B2(G128), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT96), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n540), .A2(new_n221), .A3(G143), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n279), .A2(G128), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n542), .A2(new_n293), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n293), .B1(new_n542), .B2(new_n543), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n538), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT13), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n542), .B(new_n543), .C1(new_n547), .C2(new_n293), .ZN(new_n548));
  INV_X1    g362(.A(new_n538), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n397), .B1(new_n533), .B2(new_n537), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n542), .A2(new_n547), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n545), .A2(new_n552), .ZN(new_n553));
  OAI22_X1  g367(.A1(new_n536), .A2(new_n546), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n461), .A2(G217), .A3(new_n465), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n555), .ZN(new_n557));
  OAI221_X1 g371(.A(new_n557), .B1(new_n551), .B2(new_n553), .C1(new_n536), .C2(new_n546), .ZN(new_n558));
  AOI21_X1  g372(.A(G902), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(G478), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n560), .A2(KEYINPUT15), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n559), .A2(new_n562), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(G234), .A2(G237), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(G952), .A3(new_n465), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT21), .B(G898), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(G902), .A3(G953), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n528), .A2(new_n565), .A3(new_n572), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n459), .A2(new_n463), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(G214), .B1(G237), .B2(G902), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT85), .ZN(new_n576));
  OAI21_X1  g390(.A(G210), .B1(G237), .B2(G902), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n281), .A2(new_n284), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n289), .A2(new_n282), .ZN(new_n580));
  OAI21_X1  g394(.A(G125), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n581), .B1(new_n339), .B2(G125), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n465), .A2(G224), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT87), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n582), .B(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n423), .A2(new_n274), .A3(new_n424), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n264), .A2(new_n266), .A3(KEYINPUT72), .ZN(new_n587));
  AOI21_X1  g401(.A(KEYINPUT72), .B1(new_n264), .B2(new_n266), .ZN(new_n588));
  OAI21_X1  g402(.A(KEYINPUT5), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(G113), .B1(new_n264), .B2(KEYINPUT5), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n592), .A2(new_n412), .A3(new_n273), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT6), .ZN(new_n595));
  XNOR2_X1  g409(.A(G110), .B(G122), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n586), .A2(new_n593), .A3(new_n596), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(KEYINPUT6), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n596), .B1(new_n586), .B2(new_n593), .ZN(new_n601));
  OAI211_X1 g415(.A(KEYINPUT86), .B(new_n598), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n601), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT86), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n603), .A2(new_n604), .A3(KEYINPUT6), .A4(new_n599), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n585), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n584), .A2(KEYINPUT7), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n582), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n607), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n581), .B(new_n609), .C1(new_n339), .C2(G125), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n592), .A2(new_n273), .A3(new_n410), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n264), .A2(new_n266), .A3(KEYINPUT5), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n273), .B1(new_n612), .B2(new_n590), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n412), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n596), .B(KEYINPUT8), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n611), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n608), .A2(new_n599), .A3(new_n610), .A4(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n250), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n578), .B1(new_n606), .B2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT88), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OAI211_X1 g435(.A(KEYINPUT88), .B(new_n578), .C1(new_n606), .C2(new_n618), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n602), .A2(new_n605), .ZN(new_n624));
  INV_X1    g438(.A(new_n585), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n618), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n577), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT89), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n606), .A2(new_n578), .A3(new_n618), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT89), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n576), .B1(new_n623), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n391), .A2(new_n574), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G101), .ZN(G3));
  NAND2_X1  g450(.A1(new_n459), .A2(new_n463), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n368), .A2(new_n250), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT97), .ZN(new_n639));
  INV_X1    g453(.A(G472), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n368), .B(new_n250), .C1(new_n639), .C2(new_n640), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n262), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n637), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT98), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n577), .B1(new_n626), .B2(new_n627), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n575), .B1(new_n647), .B2(new_n630), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n556), .A2(new_n558), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(KEYINPUT33), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT33), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n556), .A2(new_n558), .A3(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n650), .A2(new_n652), .A3(G478), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n560), .A2(new_n250), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n654), .B1(new_n559), .B2(new_n560), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n528), .A2(new_n657), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n648), .A2(new_n658), .A3(new_n572), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n646), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT34), .B(G104), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G6));
  AOI21_X1  g476(.A(new_n526), .B1(new_n563), .B2(new_n564), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT99), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n516), .A2(new_n664), .A3(new_n522), .ZN(new_n665));
  OAI211_X1 g479(.A(KEYINPUT99), .B(KEYINPUT20), .C1(new_n513), .C2(new_n515), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n648), .A2(new_n667), .A3(new_n572), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n646), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT35), .B(G107), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G9));
  INV_X1    g485(.A(new_n260), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n236), .A2(new_n241), .A3(KEYINPUT100), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT100), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n246), .B2(new_n248), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n192), .A2(KEYINPUT36), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n674), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  OAI22_X1  g493(.A1(new_n673), .A2(new_n676), .B1(KEYINPUT36), .B2(new_n192), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n672), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n258), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n642), .A2(new_n643), .A3(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT101), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n642), .A2(new_n683), .A3(new_n643), .A4(KEYINPUT101), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n574), .A2(new_n686), .A3(new_n634), .A4(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(KEYINPUT37), .B(G110), .Z(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G12));
  OR2_X1    g504(.A1(new_n570), .A2(G900), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n567), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n663), .A2(new_n665), .A3(new_n666), .A4(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n575), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n695), .B1(new_n628), .B2(new_n619), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n694), .A2(KEYINPUT102), .A3(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT102), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n698), .B1(new_n648), .B2(new_n693), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n257), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n701), .B1(new_n252), .B2(new_n253), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n681), .B1(new_n702), .B2(new_n255), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n703), .B1(new_n372), .B2(new_n390), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n454), .A2(new_n455), .A3(new_n250), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(KEYINPUT84), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n457), .A2(new_n450), .A3(new_n455), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n462), .B1(new_n708), .B2(new_n449), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n700), .A2(new_n704), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G128), .ZN(G30));
  NAND2_X1  g525(.A1(new_n368), .A2(new_n369), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT32), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n368), .A2(KEYINPUT32), .A3(new_n369), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n383), .A2(new_n384), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n250), .B1(new_n716), .B2(new_n352), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n352), .B1(new_n346), .B2(new_n374), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(G472), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n714), .A2(new_n715), .A3(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n528), .A2(new_n565), .ZN(new_n723));
  NOR4_X1   g537(.A1(new_n722), .A2(new_n695), .A3(new_n683), .A4(new_n723), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n618), .B1(new_n624), .B2(new_n625), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n631), .B1(new_n725), .B2(new_n577), .ZN(new_n726));
  NOR4_X1   g540(.A1(new_n606), .A2(KEYINPUT89), .A3(new_n618), .A4(new_n578), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n621), .B(new_n622), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n729));
  XOR2_X1   g543(.A(new_n728), .B(new_n729), .Z(new_n730));
  NAND3_X1  g544(.A1(new_n724), .A2(new_n730), .A3(KEYINPUT104), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n692), .B(KEYINPUT39), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n637), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(KEYINPUT40), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n724), .A2(new_n730), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n736), .B1(KEYINPUT104), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G143), .ZN(G45));
  NAND3_X1  g553(.A1(new_n528), .A2(new_n657), .A3(new_n692), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT105), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n526), .B1(new_n516), .B2(new_n522), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n656), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(KEYINPUT105), .A3(new_n692), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n742), .A2(new_n745), .A3(new_n696), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT106), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT106), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n742), .A2(new_n745), .A3(new_n748), .A4(new_n696), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n747), .A2(new_n709), .A3(new_n704), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G146), .ZN(G48));
  NAND2_X1  g565(.A1(new_n372), .A2(new_n390), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n457), .A2(new_n455), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n463), .B(new_n753), .C1(new_n456), .C2(new_n458), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n752), .A2(new_n659), .A3(new_n755), .A4(new_n262), .ZN(new_n756));
  XNOR2_X1  g570(.A(KEYINPUT41), .B(G113), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n756), .B(new_n757), .ZN(G15));
  NAND4_X1  g572(.A1(new_n752), .A2(new_n668), .A3(new_n755), .A4(new_n262), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G116), .ZN(G18));
  NOR2_X1   g574(.A1(new_n754), .A2(new_n648), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n761), .A2(new_n752), .A3(new_n573), .A4(new_n683), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G119), .ZN(G21));
  NOR2_X1   g577(.A1(new_n648), .A2(new_n723), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n755), .A2(new_n764), .A3(new_n571), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n638), .A2(G472), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT107), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n387), .A2(new_n388), .A3(new_n360), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n354), .A2(new_n367), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n369), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n638), .A2(new_n772), .A3(G472), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n767), .A2(new_n771), .A3(new_n262), .A4(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(KEYINPUT108), .B1(new_n765), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n772), .B1(new_n638), .B2(G472), .ZN(new_n776));
  AOI211_X1 g590(.A(KEYINPUT107), .B(new_n640), .C1(new_n368), .C2(new_n250), .ZN(new_n777));
  INV_X1    g591(.A(new_n369), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n778), .B1(new_n768), .B2(new_n769), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  AOI22_X1  g594(.A1(new_n523), .A2(new_n527), .B1(new_n563), .B2(new_n564), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n696), .A2(new_n571), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n754), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT108), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n780), .A2(new_n783), .A3(new_n784), .A4(new_n262), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n775), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G122), .ZN(G24));
  AOI21_X1  g601(.A(KEYINPUT105), .B1(new_n744), .B2(new_n692), .ZN(new_n788));
  INV_X1    g602(.A(new_n692), .ZN(new_n789));
  NOR4_X1   g603(.A1(new_n743), .A2(new_n656), .A3(new_n741), .A4(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n780), .A2(new_n791), .A3(new_n761), .A4(new_n683), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G125), .ZN(G27));
  NOR2_X1   g607(.A1(new_n728), .A2(new_n695), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n391), .A2(new_n709), .A3(new_n791), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n623), .A2(new_n575), .A3(new_n633), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n798), .A2(new_n637), .ZN(new_n799));
  XNOR2_X1  g613(.A(KEYINPUT109), .B(KEYINPUT42), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n799), .A2(new_n391), .A3(new_n791), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G131), .ZN(G33));
  XOR2_X1   g617(.A(new_n693), .B(KEYINPUT110), .Z(new_n804));
  NAND3_X1  g618(.A1(new_n799), .A2(new_n391), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G134), .ZN(G36));
  AND2_X1   g620(.A1(new_n448), .A2(KEYINPUT45), .ZN(new_n807));
  OAI21_X1  g621(.A(G469), .B1(new_n448), .B2(KEYINPUT45), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT111), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n455), .A2(new_n250), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n812), .A2(KEYINPUT46), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n708), .B1(new_n812), .B2(KEYINPUT46), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n463), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n657), .A2(new_n743), .ZN(new_n816));
  XOR2_X1   g630(.A(new_n816), .B(KEYINPUT43), .Z(new_n817));
  NAND2_X1  g631(.A1(new_n642), .A2(new_n643), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n817), .A2(new_n818), .A3(new_n683), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n798), .B1(new_n819), .B2(KEYINPUT44), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n820), .B1(KEYINPUT44), .B2(new_n819), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n815), .A2(new_n821), .A3(new_n733), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(new_n309), .ZN(G39));
  INV_X1    g637(.A(KEYINPUT47), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n815), .B(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n791), .ZN(new_n826));
  NOR4_X1   g640(.A1(new_n826), .A2(new_n752), .A3(new_n798), .A4(new_n262), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(G140), .ZN(G42));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n704), .A2(new_n749), .A3(new_n709), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n748), .B1(new_n791), .B2(new_n696), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n710), .B(new_n792), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n696), .A2(new_n703), .A3(new_n692), .A4(new_n781), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n637), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT113), .B1(new_n836), .B2(new_n721), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n258), .A2(new_n682), .A3(new_n692), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n648), .A2(new_n838), .A3(new_n723), .ZN(new_n839));
  AND4_X1   g653(.A1(KEYINPUT113), .A2(new_n839), .A3(new_n709), .A4(new_n721), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n831), .B1(new_n834), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n710), .A2(new_n792), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n839), .A2(new_n709), .A3(new_n721), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n836), .A2(KEYINPUT113), .A3(new_n721), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n843), .A2(KEYINPUT52), .A3(new_n750), .A4(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n842), .A2(new_n849), .A3(KEYINPUT114), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT114), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n851), .B(new_n831), .C1(new_n834), .C2(new_n841), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT112), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n634), .A2(new_n854), .A3(new_n571), .A4(new_n744), .ZN(new_n855));
  INV_X1    g669(.A(new_n576), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n728), .A2(new_n856), .A3(new_n571), .A4(new_n744), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(KEYINPUT112), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n855), .A2(new_n645), .A3(new_n858), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n728), .A2(new_n856), .A3(new_n571), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n663), .A2(new_n523), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n645), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n859), .A2(new_n635), .A3(new_n688), .A4(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n762), .A2(new_n756), .A3(new_n759), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n866), .B1(new_n785), .B2(new_n775), .ZN(new_n867));
  NOR4_X1   g681(.A1(new_n777), .A2(new_n776), .A3(new_n779), .A4(new_n703), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n868), .A2(new_n799), .A3(new_n791), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n665), .A2(new_n666), .ZN(new_n870));
  NOR4_X1   g684(.A1(new_n870), .A2(new_n526), .A3(new_n565), .A4(new_n789), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n704), .A2(new_n709), .A3(new_n794), .A4(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n869), .A2(new_n805), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n865), .A2(new_n867), .A3(new_n802), .A4(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n830), .B1(new_n853), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n842), .A2(new_n849), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n855), .A2(new_n645), .A3(new_n858), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n863), .A2(new_n688), .A3(new_n635), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n873), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n877), .A2(new_n802), .A3(new_n867), .A4(new_n880), .ZN(new_n881));
  XNOR2_X1  g695(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n876), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT116), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n884), .A3(KEYINPUT54), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n842), .A2(new_n849), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n886), .A2(new_n875), .ZN(new_n887));
  INV_X1    g701(.A(new_n882), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n797), .A2(new_n801), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n762), .A2(new_n756), .A3(new_n759), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n786), .ZN(new_n891));
  OAI21_X1  g705(.A(KEYINPUT117), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n864), .A2(new_n830), .A3(new_n873), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT117), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n802), .A2(new_n894), .A3(new_n786), .A4(new_n890), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  OAI22_X1  g710(.A1(new_n887), .A2(new_n888), .B1(new_n853), .B2(new_n896), .ZN(new_n897));
  OR2_X1    g711(.A1(new_n897), .A2(KEYINPUT54), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n885), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n884), .B1(new_n883), .B2(KEYINPUT54), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n567), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n817), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n774), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n708), .A2(new_n753), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n907), .A2(new_n463), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n794), .B(new_n906), .C1(new_n825), .C2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n798), .A2(new_n754), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n910), .A2(new_n262), .A3(new_n902), .A4(new_n722), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n911), .A2(new_n528), .A3(new_n657), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n903), .A2(new_n910), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n912), .B1(new_n868), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT51), .ZN(new_n916));
  NOR4_X1   g730(.A1(new_n905), .A2(new_n575), .A3(new_n730), .A4(new_n754), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n917), .A2(KEYINPUT50), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(KEYINPUT50), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n909), .A2(new_n915), .A3(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT119), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n914), .A2(new_n391), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT48), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n465), .A2(G952), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n911), .A2(new_n658), .ZN(new_n926));
  AOI211_X1 g740(.A(new_n925), .B(new_n926), .C1(new_n761), .C2(new_n906), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n918), .A2(new_n919), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n929), .A2(KEYINPUT118), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(KEYINPUT118), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n930), .A2(new_n909), .A3(new_n915), .A4(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n928), .B1(new_n932), .B2(new_n916), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n901), .A2(new_n922), .A3(new_n933), .ZN(new_n934));
  OR2_X1    g748(.A1(G952), .A2(G953), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n730), .ZN(new_n937));
  NOR4_X1   g751(.A1(new_n263), .A2(new_n816), .A3(new_n576), .A4(new_n462), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n907), .B(KEYINPUT49), .Z(new_n939));
  NAND4_X1  g753(.A1(new_n937), .A2(new_n722), .A3(new_n938), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n936), .A2(new_n940), .ZN(G75));
  AND2_X1   g755(.A1(new_n850), .A2(new_n852), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n943));
  AOI22_X1  g757(.A1(new_n942), .A2(new_n943), .B1(new_n881), .B2(new_n882), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n944), .A2(new_n250), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(G210), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n624), .A2(new_n625), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n947), .A2(new_n606), .ZN(new_n948));
  XNOR2_X1  g762(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(new_n950));
  XNOR2_X1  g764(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n946), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT122), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n465), .A2(G952), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT56), .B1(new_n945), .B2(G210), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n955), .B1(new_n956), .B2(new_n950), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n953), .A2(new_n957), .ZN(G51));
  XNOR2_X1  g772(.A(new_n897), .B(KEYINPUT54), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n811), .B(KEYINPUT57), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n454), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n945), .A2(new_n810), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n954), .B1(new_n962), .B2(new_n963), .ZN(G54));
  NAND3_X1  g778(.A1(new_n945), .A2(KEYINPUT58), .A3(G475), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n965), .A2(new_n513), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n965), .A2(new_n513), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n966), .A2(new_n967), .A3(new_n954), .ZN(G60));
  NAND2_X1  g782(.A1(new_n650), .A2(new_n652), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n654), .B(KEYINPUT59), .Z(new_n970));
  AND3_X1   g784(.A1(new_n959), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n969), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n970), .B1(new_n899), .B2(new_n900), .ZN(new_n973));
  AOI211_X1 g787(.A(new_n954), .B(new_n971), .C1(new_n972), .C2(new_n973), .ZN(G63));
  NAND2_X1  g788(.A1(G217), .A2(G902), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT60), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n880), .A2(new_n895), .A3(KEYINPUT53), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n977), .A2(new_n852), .A3(new_n850), .A4(new_n892), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n881), .A2(new_n882), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n976), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n679), .A2(new_n680), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n259), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n983), .B1(new_n944), .B2(new_n976), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n982), .A2(new_n984), .A3(KEYINPUT61), .A4(new_n955), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT61), .ZN(new_n986));
  OAI211_X1 g800(.A(KEYINPUT123), .B(new_n955), .C1(new_n980), .C2(new_n259), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n982), .ZN(new_n988));
  AOI21_X1  g802(.A(KEYINPUT123), .B1(new_n984), .B2(new_n955), .ZN(new_n989));
  OAI211_X1 g803(.A(KEYINPUT124), .B(new_n986), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT123), .ZN(new_n992));
  INV_X1    g806(.A(new_n976), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n259), .B1(new_n897), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n992), .B1(new_n994), .B2(new_n954), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n995), .A2(new_n987), .A3(new_n982), .ZN(new_n996));
  AOI21_X1  g810(.A(KEYINPUT124), .B1(new_n996), .B2(new_n986), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n985), .B1(new_n991), .B2(new_n997), .ZN(G66));
  INV_X1    g812(.A(G224), .ZN(new_n999));
  OAI21_X1  g813(.A(G953), .B1(new_n568), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n891), .A2(new_n864), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n1000), .B1(new_n1001), .B2(G953), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n602), .B(new_n605), .C1(G898), .C2(new_n465), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1002), .B(new_n1003), .ZN(G69));
  AOI21_X1  g818(.A(new_n822), .B1(new_n825), .B2(new_n827), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n391), .A2(new_n764), .ZN(new_n1006));
  NOR3_X1   g820(.A1(new_n815), .A2(new_n733), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(new_n834), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1008), .A2(new_n802), .A3(new_n805), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1005), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1011), .A2(G953), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n335), .A2(new_n345), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n498), .A2(new_n503), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1013), .B(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(G900), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1015), .B1(new_n1016), .B2(new_n465), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n1012), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT62), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n738), .A2(new_n1019), .A3(new_n1008), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(KEYINPUT126), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n799), .A2(new_n391), .ZN(new_n1022));
  AOI211_X1 g836(.A(new_n733), .B(new_n1022), .C1(new_n658), .C2(new_n861), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n738), .A2(new_n1008), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1023), .B1(new_n1024), .B2(KEYINPUT62), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1021), .A2(new_n1005), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1026), .A2(new_n465), .ZN(new_n1027));
  XOR2_X1   g841(.A(new_n1015), .B(KEYINPUT125), .Z(new_n1028));
  AOI21_X1  g842(.A(new_n1018), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g843(.A(G953), .B1(new_n438), .B2(new_n1016), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n1029), .B(new_n1030), .ZN(G72));
  NAND4_X1  g845(.A1(new_n1021), .A2(new_n1001), .A3(new_n1005), .A4(new_n1025), .ZN(new_n1032));
  NAND2_X1  g846(.A1(G472), .A2(G902), .ZN(new_n1033));
  XOR2_X1   g847(.A(new_n1033), .B(KEYINPUT63), .Z(new_n1034));
  NAND2_X1  g848(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1035), .A2(new_n719), .ZN(new_n1036));
  INV_X1    g850(.A(new_n375), .ZN(new_n1037));
  NAND4_X1  g851(.A1(new_n883), .A2(new_n1037), .A3(new_n718), .A4(new_n1034), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1001), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1034), .B1(new_n1011), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n954), .B1(new_n1040), .B2(new_n375), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n1036), .A2(new_n1038), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1042), .A2(KEYINPUT127), .ZN(new_n1043));
  INV_X1    g857(.A(KEYINPUT127), .ZN(new_n1044));
  NAND4_X1  g858(.A1(new_n1036), .A2(new_n1041), .A3(new_n1044), .A4(new_n1038), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1043), .A2(new_n1045), .ZN(G57));
endmodule


