

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784;

  XNOR2_X1 U376 ( .A(n386), .B(n364), .ZN(n609) );
  XNOR2_X1 U377 ( .A(n577), .B(G146), .ZN(n529) );
  XNOR2_X1 U378 ( .A(G134), .B(G107), .ZN(n492) );
  XNOR2_X1 U379 ( .A(n474), .B(KEYINPUT3), .ZN(n476) );
  NAND2_X1 U380 ( .A1(n646), .A2(n645), .ZN(n622) );
  AND2_X2 U381 ( .A1(n717), .A2(n621), .ZN(n646) );
  NAND2_X1 U382 ( .A1(n590), .A2(n683), .ZN(n633) );
  XNOR2_X2 U383 ( .A(n530), .B(G469), .ZN(n590) );
  NOR2_X2 U384 ( .A1(n456), .A2(n553), .ZN(n446) );
  AND2_X2 U385 ( .A1(n447), .A2(n445), .ZN(n444) );
  NAND2_X2 U386 ( .A1(n430), .A2(n432), .ZN(n621) );
  NAND2_X2 U387 ( .A1(n568), .A2(n567), .ZN(n570) );
  OR2_X2 U388 ( .A1(n753), .A2(G902), .ZN(n530) );
  XNOR2_X1 U389 ( .A(n541), .B(n480), .ZN(n574) );
  INV_X2 U390 ( .A(G146), .ZN(n479) );
  NOR2_X1 U391 ( .A1(G953), .A2(G237), .ZN(n481) );
  XNOR2_X1 U392 ( .A(n437), .B(n620), .ZN(n717) );
  AND2_X1 U393 ( .A1(n581), .A2(n580), .ZN(n763) );
  NOR2_X2 U394 ( .A1(n685), .A2(n686), .ZN(n683) );
  INV_X1 U395 ( .A(KEYINPUT69), .ZN(n463) );
  AND2_X1 U396 ( .A1(n616), .A2(n571), .ZN(n623) );
  AND2_X1 U397 ( .A1(n391), .A2(n367), .ZN(n357) );
  NAND2_X1 U398 ( .A1(n371), .A2(n369), .ZN(n625) );
  NOR2_X1 U399 ( .A1(n373), .A2(n372), .ZN(n371) );
  AND2_X1 U400 ( .A1(n381), .A2(n380), .ZN(n379) );
  XNOR2_X1 U401 ( .A(n427), .B(n424), .ZN(n546) );
  XNOR2_X1 U402 ( .A(n541), .B(n425), .ZN(n424) );
  XNOR2_X1 U403 ( .A(KEYINPUT75), .B(KEYINPUT16), .ZN(n537) );
  XNOR2_X1 U404 ( .A(G122), .B(KEYINPUT74), .ZN(n536) );
  XNOR2_X1 U405 ( .A(G113), .B(KEYINPUT71), .ZN(n475) );
  XNOR2_X1 U406 ( .A(n354), .B(n355), .ZN(n711) );
  NOR2_X1 U407 ( .A1(n629), .A2(n625), .ZN(n354) );
  XOR2_X1 U408 ( .A(n560), .B(KEYINPUT33), .Z(n355) );
  XNOR2_X1 U409 ( .A(n545), .B(n544), .ZN(n427) );
  INV_X2 U410 ( .A(n628), .ZN(n635) );
  NOR2_X2 U411 ( .A1(n678), .A2(n677), .ZN(n679) );
  OR2_X1 U412 ( .A1(n718), .A2(n452), .ZN(n451) );
  XNOR2_X2 U413 ( .A(n559), .B(n558), .ZN(n568) );
  OR2_X2 U414 ( .A1(n592), .A2(n557), .ZN(n559) );
  NOR2_X1 U415 ( .A1(n450), .A2(n601), .ZN(n449) );
  XNOR2_X1 U416 ( .A(n388), .B(n462), .ZN(n387) );
  INV_X1 U417 ( .A(KEYINPUT46), .ZN(n462) );
  OR2_X1 U418 ( .A1(n781), .A2(n782), .ZN(n388) );
  NAND2_X1 U419 ( .A1(n379), .A2(n375), .ZN(n572) );
  INV_X1 U420 ( .A(KEYINPUT15), .ZN(n500) );
  XNOR2_X1 U421 ( .A(G902), .B(KEYINPUT97), .ZN(n501) );
  XNOR2_X1 U422 ( .A(n545), .B(n409), .ZN(n577) );
  XNOR2_X1 U423 ( .A(n467), .B(KEYINPUT4), .ZN(n409) );
  NOR2_X1 U424 ( .A1(n633), .A2(n582), .ZN(n368) );
  NAND2_X1 U425 ( .A1(n444), .A2(n440), .ZN(n579) );
  NAND2_X1 U426 ( .A1(n443), .A2(n441), .ZN(n440) );
  NOR2_X1 U427 ( .A1(n379), .A2(n374), .ZN(n372) );
  XNOR2_X1 U428 ( .A(KEYINPUT67), .B(G137), .ZN(n525) );
  INV_X1 U429 ( .A(G140), .ZN(n526) );
  XNOR2_X1 U430 ( .A(n525), .B(KEYINPUT101), .ZN(n575) );
  XNOR2_X1 U431 ( .A(n600), .B(KEYINPUT39), .ZN(n396) );
  AND2_X1 U432 ( .A1(n357), .A2(n697), .ZN(n600) );
  NOR2_X1 U433 ( .A1(n436), .A2(n624), .ZN(n435) );
  NOR2_X1 U434 ( .A1(n632), .A2(n573), .ZN(n436) );
  INV_X2 U435 ( .A(G953), .ZN(n726) );
  XNOR2_X1 U436 ( .A(n461), .B(n460), .ZN(n459) );
  INV_X1 U437 ( .A(KEYINPUT85), .ZN(n460) );
  XNOR2_X1 U438 ( .A(n767), .B(n405), .ZN(n404) );
  INV_X1 U439 ( .A(KEYINPUT47), .ZN(n405) );
  AND2_X1 U440 ( .A1(n646), .A2(n644), .ZN(n412) );
  INV_X1 U441 ( .A(KEYINPUT73), .ZN(n410) );
  NAND2_X1 U442 ( .A1(G237), .A2(G234), .ZN(n506) );
  INV_X1 U443 ( .A(G237), .ZN(n531) );
  XNOR2_X1 U444 ( .A(G101), .B(G137), .ZN(n471) );
  INV_X1 U445 ( .A(KEYINPUT103), .ZN(n470) );
  XOR2_X1 U446 ( .A(KEYINPUT104), .B(KEYINPUT5), .Z(n469) );
  XNOR2_X1 U447 ( .A(n421), .B(n420), .ZN(n511) );
  INV_X1 U448 ( .A(KEYINPUT8), .ZN(n420) );
  NAND2_X1 U449 ( .A1(n726), .A2(G234), .ZN(n421) );
  XNOR2_X1 U450 ( .A(n457), .B(KEYINPUT11), .ZN(n486) );
  INV_X1 U451 ( .A(KEYINPUT105), .ZN(n457) );
  XNOR2_X1 U452 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n543) );
  XNOR2_X1 U453 ( .A(n426), .B(KEYINPUT4), .ZN(n425) );
  XNOR2_X1 U454 ( .A(KEYINPUT79), .B(KEYINPUT98), .ZN(n426) );
  NAND2_X1 U455 ( .A1(n550), .A2(n650), .ZN(n455) );
  NAND2_X1 U456 ( .A1(n454), .A2(n453), .ZN(n452) );
  INV_X1 U457 ( .A(n650), .ZN(n453) );
  INV_X1 U458 ( .A(n550), .ZN(n454) );
  OR2_X1 U459 ( .A1(n665), .A2(n376), .ZN(n375) );
  NAND2_X1 U460 ( .A1(n378), .A2(n377), .ZN(n376) );
  INV_X1 U461 ( .A(G472), .ZN(n378) );
  INV_X1 U462 ( .A(KEYINPUT6), .ZN(n374) );
  NAND2_X1 U463 ( .A1(G902), .A2(G472), .ZN(n380) );
  XNOR2_X1 U464 ( .A(G128), .B(G110), .ZN(n514) );
  XOR2_X1 U465 ( .A(G122), .B(G116), .Z(n493) );
  NOR2_X1 U466 ( .A1(n588), .A2(n423), .ZN(n578) );
  OR2_X1 U467 ( .A1(n625), .A2(n769), .ZN(n423) );
  XNOR2_X1 U468 ( .A(n393), .B(n392), .ZN(n391) );
  XNOR2_X1 U469 ( .A(n579), .B(KEYINPUT19), .ZN(n592) );
  XNOR2_X1 U470 ( .A(n466), .B(n465), .ZN(n581) );
  XNOR2_X1 U471 ( .A(n491), .B(n744), .ZN(n465) );
  XNOR2_X1 U472 ( .A(n464), .B(G478), .ZN(n580) );
  NOR2_X1 U473 ( .A1(n434), .A2(n433), .ZN(n747) );
  BUF_X1 U474 ( .A(n739), .Z(n751) );
  XNOR2_X1 U475 ( .A(n529), .B(n407), .ZN(n753) );
  XNOR2_X1 U476 ( .A(n408), .B(n575), .ZN(n407) );
  XNOR2_X1 U477 ( .A(n670), .B(n669), .ZN(n778) );
  INV_X1 U478 ( .A(n606), .ZN(n395) );
  XNOR2_X1 U479 ( .A(n366), .B(n365), .ZN(n782) );
  INV_X1 U480 ( .A(KEYINPUT40), .ZN(n365) );
  OR2_X1 U481 ( .A1(n396), .A2(n769), .ZN(n366) );
  XNOR2_X1 U482 ( .A(n382), .B(KEYINPUT113), .ZN(n419) );
  XNOR2_X1 U483 ( .A(n385), .B(n384), .ZN(n383) );
  INV_X1 U484 ( .A(KEYINPUT36), .ZN(n384) );
  NAND2_X1 U485 ( .A1(n429), .A2(n431), .ZN(n432) );
  NAND2_X1 U486 ( .A1(n435), .A2(n573), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n627), .B(KEYINPUT109), .ZN(n779) );
  INV_X1 U488 ( .A(KEYINPUT53), .ZN(n397) );
  INV_X1 U489 ( .A(G953), .ZN(n399) );
  AND2_X1 U490 ( .A1(n751), .A2(G478), .ZN(n356) );
  INV_X1 U491 ( .A(n572), .ZN(n632) );
  AND2_X1 U492 ( .A1(n609), .A2(n608), .ZN(n358) );
  INV_X1 U493 ( .A(G902), .ZN(n377) );
  AND2_X1 U494 ( .A1(n618), .A2(n617), .ZN(n359) );
  AND2_X1 U495 ( .A1(n632), .A2(n573), .ZN(n360) );
  AND2_X1 U496 ( .A1(n451), .A2(n455), .ZN(n361) );
  AND2_X1 U497 ( .A1(n435), .A2(n571), .ZN(n362) );
  AND2_X1 U498 ( .A1(n608), .A2(KEYINPUT2), .ZN(n363) );
  INV_X1 U499 ( .A(KEYINPUT66), .ZN(n573) );
  XNOR2_X1 U500 ( .A(n532), .B(KEYINPUT99), .ZN(n601) );
  INV_X1 U501 ( .A(n601), .ZN(n394) );
  XOR2_X1 U502 ( .A(n605), .B(KEYINPUT91), .Z(n364) );
  XNOR2_X1 U503 ( .A(n368), .B(KEYINPUT78), .ZN(n367) );
  NAND2_X1 U504 ( .A1(n370), .A2(n379), .ZN(n369) );
  AND2_X1 U505 ( .A1(n375), .A2(n374), .ZN(n370) );
  NOR2_X1 U506 ( .A1(n375), .A2(n374), .ZN(n373) );
  NAND2_X1 U507 ( .A1(n665), .A2(G472), .ZN(n381) );
  NAND2_X1 U508 ( .A1(n383), .A2(n682), .ZN(n382) );
  NAND2_X1 U509 ( .A1(n422), .A2(n579), .ZN(n385) );
  NAND2_X1 U510 ( .A1(n389), .A2(n387), .ZN(n386) );
  XNOR2_X1 U511 ( .A(n390), .B(n463), .ZN(n389) );
  NOR2_X2 U512 ( .A1(n599), .A2(n419), .ZN(n390) );
  INV_X1 U513 ( .A(KEYINPUT30), .ZN(n392) );
  NAND2_X1 U514 ( .A1(n572), .A2(n394), .ZN(n393) );
  OR2_X1 U515 ( .A1(n396), .A2(n395), .ZN(n775) );
  XNOR2_X1 U516 ( .A(n398), .B(n397), .ZN(G75) );
  NAND2_X1 U517 ( .A1(n400), .A2(n399), .ZN(n398) );
  XNOR2_X1 U518 ( .A(n402), .B(n401), .ZN(n400) );
  INV_X1 U519 ( .A(KEYINPUT120), .ZN(n401) );
  NAND2_X1 U520 ( .A1(n715), .A2(n714), .ZN(n402) );
  XNOR2_X1 U521 ( .A(n403), .B(n528), .ZN(n408) );
  XNOR2_X2 U522 ( .A(n403), .B(n538), .ZN(n540) );
  XNOR2_X2 U523 ( .A(n439), .B(n438), .ZN(n403) );
  XNOR2_X1 U524 ( .A(n411), .B(n410), .ZN(n647) );
  NAND2_X1 U525 ( .A1(n595), .A2(n404), .ZN(n596) );
  XNOR2_X1 U526 ( .A(n598), .B(KEYINPUT76), .ZN(n599) );
  NAND2_X1 U527 ( .A1(n623), .A2(n360), .ZN(n430) );
  NOR2_X1 U528 ( .A1(n406), .A2(n779), .ZN(n640) );
  XNOR2_X1 U529 ( .A(n639), .B(n638), .ZN(n406) );
  XNOR2_X2 U530 ( .A(n631), .B(n630), .ZN(n771) );
  XNOR2_X1 U531 ( .A(n517), .B(n518), .ZN(n740) );
  NOR2_X2 U532 ( .A1(n603), .A2(n593), .ZN(n767) );
  NAND2_X1 U533 ( .A1(n680), .A2(n681), .ZN(n715) );
  XNOR2_X2 U534 ( .A(n476), .B(n475), .ZN(n539) );
  XNOR2_X2 U535 ( .A(n733), .B(n546), .ZN(n718) );
  XNOR2_X2 U536 ( .A(n540), .B(n539), .ZN(n733) );
  XNOR2_X2 U537 ( .A(n428), .B(G128), .ZN(n545) );
  NAND2_X1 U538 ( .A1(n412), .A2(n645), .ZN(n411) );
  NAND2_X1 U539 ( .A1(n413), .A2(n561), .ZN(n417) );
  NAND2_X1 U540 ( .A1(n414), .A2(n635), .ZN(n413) );
  INV_X1 U541 ( .A(n711), .ZN(n414) );
  NAND2_X1 U542 ( .A1(n415), .A2(n635), .ZN(n416) );
  NOR2_X1 U543 ( .A1(n711), .A2(n561), .ZN(n415) );
  NAND2_X1 U544 ( .A1(n417), .A2(n416), .ZN(n418) );
  NAND2_X1 U545 ( .A1(n418), .A2(n583), .ZN(n564) );
  XNOR2_X1 U546 ( .A(n419), .B(KEYINPUT118), .ZN(n783) );
  NAND2_X1 U547 ( .A1(n511), .A2(G221), .ZN(n512) );
  NAND2_X1 U548 ( .A1(n609), .A2(n363), .ZN(n658) );
  XNOR2_X1 U549 ( .A(n578), .B(KEYINPUT112), .ZN(n422) );
  XNOR2_X2 U550 ( .A(n479), .B(G125), .ZN(n541) );
  XNOR2_X2 U551 ( .A(G143), .B(KEYINPUT64), .ZN(n428) );
  NAND2_X1 U552 ( .A1(n616), .A2(n362), .ZN(n429) );
  XNOR2_X2 U553 ( .A(G119), .B(G116), .ZN(n474) );
  AND2_X2 U554 ( .A1(n662), .A2(n681), .ZN(n739) );
  NAND2_X1 U555 ( .A1(n587), .A2(n459), .ZN(n458) );
  INV_X1 U556 ( .A(n662), .ZN(n433) );
  NAND2_X1 U557 ( .A1(n681), .A2(G475), .ZN(n434) );
  NAND2_X1 U558 ( .A1(n616), .A2(n359), .ZN(n437) );
  XNOR2_X2 U559 ( .A(G110), .B(G107), .ZN(n438) );
  XNOR2_X2 U560 ( .A(G104), .B(G101), .ZN(n439) );
  NOR2_X1 U561 ( .A1(n442), .A2(KEYINPUT93), .ZN(n441) );
  INV_X1 U562 ( .A(n456), .ZN(n442) );
  INV_X1 U563 ( .A(n448), .ZN(n443) );
  INV_X1 U564 ( .A(n446), .ZN(n445) );
  NAND2_X1 U565 ( .A1(n448), .A2(KEYINPUT93), .ZN(n447) );
  NAND2_X1 U566 ( .A1(n361), .A2(n456), .ZN(n552) );
  NAND2_X1 U567 ( .A1(n451), .A2(n449), .ZN(n448) );
  INV_X1 U568 ( .A(n455), .ZN(n450) );
  NAND2_X1 U569 ( .A1(n718), .A2(n550), .ZN(n456) );
  XNOR2_X1 U570 ( .A(n458), .B(KEYINPUT83), .ZN(n597) );
  NAND2_X1 U571 ( .A1(n700), .A2(KEYINPUT47), .ZN(n461) );
  INV_X1 U572 ( .A(n580), .ZN(n566) );
  NAND2_X1 U573 ( .A1(n776), .A2(n377), .ZN(n464) );
  NOR2_X1 U574 ( .A1(n745), .A2(G902), .ZN(n466) );
  XNOR2_X2 U575 ( .A(n522), .B(n521), .ZN(n685) );
  INV_X1 U576 ( .A(KEYINPUT87), .ZN(n586) );
  XNOR2_X1 U577 ( .A(n674), .B(n586), .ZN(n587) );
  INV_X1 U578 ( .A(KEYINPUT92), .ZN(n642) );
  XNOR2_X1 U579 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U580 ( .A(n473), .B(n472), .ZN(n477) );
  XNOR2_X1 U581 ( .A(n527), .B(n526), .ZN(n528) );
  INV_X1 U582 ( .A(KEYINPUT93), .ZN(n553) );
  BUF_X1 U583 ( .A(n592), .Z(n593) );
  XNOR2_X1 U584 ( .A(G131), .B(G134), .ZN(n467) );
  NAND2_X1 U585 ( .A1(G210), .A2(n481), .ZN(n468) );
  XNOR2_X1 U586 ( .A(n469), .B(n468), .ZN(n473) );
  XNOR2_X1 U587 ( .A(n477), .B(n539), .ZN(n478) );
  XNOR2_X1 U588 ( .A(n529), .B(n478), .ZN(n665) );
  XNOR2_X1 U589 ( .A(G140), .B(KEYINPUT10), .ZN(n480) );
  NAND2_X1 U590 ( .A1(n481), .A2(G214), .ZN(n482) );
  XNOR2_X1 U591 ( .A(n574), .B(n482), .ZN(n490) );
  XOR2_X1 U592 ( .A(G113), .B(G104), .Z(n484) );
  XNOR2_X1 U593 ( .A(G143), .B(G131), .ZN(n483) );
  XNOR2_X1 U594 ( .A(n484), .B(n483), .ZN(n488) );
  XNOR2_X1 U595 ( .A(G122), .B(KEYINPUT12), .ZN(n485) );
  XNOR2_X1 U596 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U597 ( .A(n488), .B(n487), .Z(n489) );
  XNOR2_X1 U598 ( .A(n490), .B(n489), .ZN(n745) );
  XNOR2_X1 U599 ( .A(KEYINPUT106), .B(KEYINPUT13), .ZN(n491) );
  INV_X1 U600 ( .A(G475), .ZN(n744) );
  XNOR2_X1 U601 ( .A(n493), .B(n492), .ZN(n495) );
  INV_X1 U602 ( .A(n545), .ZN(n494) );
  XNOR2_X1 U603 ( .A(n495), .B(n494), .ZN(n499) );
  XOR2_X1 U604 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n497) );
  NAND2_X1 U605 ( .A1(G217), .A2(n511), .ZN(n496) );
  XNOR2_X1 U606 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U607 ( .A(n499), .B(n498), .ZN(n776) );
  OR2_X1 U608 ( .A1(n581), .A2(n580), .ZN(n769) );
  XNOR2_X1 U609 ( .A(n501), .B(n500), .ZN(n654) );
  NAND2_X1 U610 ( .A1(n654), .A2(G234), .ZN(n503) );
  XNOR2_X1 U611 ( .A(KEYINPUT102), .B(KEYINPUT20), .ZN(n502) );
  XNOR2_X1 U612 ( .A(n503), .B(n502), .ZN(n519) );
  NAND2_X1 U613 ( .A1(n519), .A2(G221), .ZN(n504) );
  XNOR2_X1 U614 ( .A(n504), .B(KEYINPUT21), .ZN(n686) );
  INV_X1 U615 ( .A(KEYINPUT14), .ZN(n505) );
  XNOR2_X1 U616 ( .A(n506), .B(n505), .ZN(n509) );
  NAND2_X1 U617 ( .A1(G953), .A2(G902), .ZN(n507) );
  NOR2_X1 U618 ( .A1(n509), .A2(n507), .ZN(n554) );
  XOR2_X1 U619 ( .A(KEYINPUT110), .B(n554), .Z(n508) );
  NOR2_X1 U620 ( .A1(G900), .A2(n508), .ZN(n510) );
  INV_X1 U621 ( .A(G952), .ZN(n668) );
  OR2_X1 U622 ( .A1(n509), .A2(n668), .ZN(n708) );
  NOR2_X1 U623 ( .A1(n708), .A2(G953), .ZN(n555) );
  NOR2_X1 U624 ( .A1(n510), .A2(n555), .ZN(n582) );
  NOR2_X1 U625 ( .A1(n686), .A2(n582), .ZN(n523) );
  XNOR2_X1 U626 ( .A(n525), .B(KEYINPUT23), .ZN(n513) );
  XNOR2_X1 U627 ( .A(n513), .B(n512), .ZN(n518) );
  XOR2_X1 U628 ( .A(KEYINPUT24), .B(G119), .Z(n515) );
  XNOR2_X1 U629 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U630 ( .A(n574), .B(n516), .ZN(n517) );
  NAND2_X1 U631 ( .A1(n740), .A2(n377), .ZN(n522) );
  NAND2_X1 U632 ( .A1(G217), .A2(n519), .ZN(n520) );
  XNOR2_X1 U633 ( .A(KEYINPUT25), .B(n520), .ZN(n521) );
  NAND2_X1 U634 ( .A1(n523), .A2(n685), .ZN(n524) );
  XNOR2_X1 U635 ( .A(KEYINPUT70), .B(n524), .ZN(n588) );
  NAND2_X1 U636 ( .A1(n726), .A2(G227), .ZN(n527) );
  XNOR2_X2 U637 ( .A(n590), .B(KEYINPUT1), .ZN(n682) );
  NAND2_X1 U638 ( .A1(n377), .A2(n531), .ZN(n547) );
  NAND2_X1 U639 ( .A1(n547), .A2(G214), .ZN(n532) );
  NOR2_X1 U640 ( .A1(n682), .A2(n601), .ZN(n533) );
  NAND2_X1 U641 ( .A1(n578), .A2(n533), .ZN(n534) );
  XNOR2_X1 U642 ( .A(KEYINPUT111), .B(n534), .ZN(n535) );
  XOR2_X1 U643 ( .A(n535), .B(KEYINPUT43), .Z(n551) );
  XNOR2_X1 U644 ( .A(n537), .B(n536), .ZN(n538) );
  NAND2_X1 U645 ( .A1(n726), .A2(G224), .ZN(n542) );
  XNOR2_X1 U646 ( .A(n543), .B(n542), .ZN(n544) );
  INV_X1 U647 ( .A(n654), .ZN(n650) );
  NAND2_X1 U648 ( .A1(n547), .A2(G210), .ZN(n549) );
  INV_X1 U649 ( .A(KEYINPUT81), .ZN(n548) );
  XNOR2_X1 U650 ( .A(n549), .B(n548), .ZN(n550) );
  NAND2_X1 U651 ( .A1(n551), .A2(n552), .ZN(n607) );
  XNOR2_X1 U652 ( .A(n607), .B(G140), .ZN(G42) );
  XOR2_X1 U653 ( .A(G898), .B(KEYINPUT100), .Z(n734) );
  AND2_X1 U654 ( .A1(n734), .A2(n554), .ZN(n556) );
  NOR2_X1 U655 ( .A1(n556), .A2(n555), .ZN(n557) );
  INV_X1 U656 ( .A(KEYINPUT0), .ZN(n558) );
  INV_X1 U657 ( .A(n568), .ZN(n628) );
  NAND2_X1 U658 ( .A1(n682), .A2(n683), .ZN(n629) );
  INV_X1 U659 ( .A(KEYINPUT72), .ZN(n560) );
  INV_X1 U660 ( .A(KEYINPUT34), .ZN(n561) );
  INV_X1 U661 ( .A(n581), .ZN(n562) );
  AND2_X1 U662 ( .A1(n562), .A2(n580), .ZN(n583) );
  INV_X1 U663 ( .A(KEYINPUT35), .ZN(n563) );
  XNOR2_X2 U664 ( .A(n564), .B(n563), .ZN(n645) );
  XOR2_X1 U665 ( .A(G122), .B(KEYINPUT125), .Z(n565) );
  XNOR2_X1 U666 ( .A(n645), .B(n565), .ZN(G24) );
  NAND2_X1 U667 ( .A1(n581), .A2(n566), .ZN(n699) );
  NOR2_X1 U668 ( .A1(n699), .A2(n686), .ZN(n567) );
  INV_X1 U669 ( .A(KEYINPUT22), .ZN(n569) );
  XNOR2_X2 U670 ( .A(n570), .B(n569), .ZN(n616) );
  INV_X1 U671 ( .A(n682), .ZN(n571) );
  INV_X1 U672 ( .A(n685), .ZN(n624) );
  XNOR2_X1 U673 ( .A(n621), .B(G110), .ZN(G12) );
  XNOR2_X1 U674 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U675 ( .A(n577), .B(n576), .ZN(n611) );
  INV_X1 U676 ( .A(n769), .ZN(n766) );
  XOR2_X1 U677 ( .A(KEYINPUT107), .B(n763), .Z(n606) );
  NOR2_X1 U678 ( .A1(n766), .A2(n606), .ZN(n700) );
  INV_X1 U679 ( .A(n583), .ZN(n584) );
  NOR2_X1 U680 ( .A1(n584), .A2(n552), .ZN(n585) );
  NAND2_X1 U681 ( .A1(n357), .A2(n585), .ZN(n674) );
  NOR2_X1 U682 ( .A1(n588), .A2(n632), .ZN(n589) );
  XNOR2_X1 U683 ( .A(KEYINPUT28), .B(n589), .ZN(n591) );
  NAND2_X1 U684 ( .A1(n591), .A2(n590), .ZN(n603) );
  XOR2_X1 U685 ( .A(KEYINPUT86), .B(n700), .Z(n636) );
  INV_X1 U686 ( .A(n636), .ZN(n594) );
  NAND2_X1 U687 ( .A1(n767), .A2(n594), .ZN(n595) );
  NAND2_X1 U688 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U689 ( .A(n552), .B(KEYINPUT38), .ZN(n697) );
  NAND2_X1 U690 ( .A1(n697), .A2(n394), .ZN(n701) );
  NOR2_X1 U691 ( .A1(n701), .A2(n699), .ZN(n602) );
  XNOR2_X1 U692 ( .A(n602), .B(KEYINPUT41), .ZN(n710) );
  NOR2_X1 U693 ( .A1(n603), .A2(n710), .ZN(n604) );
  XNOR2_X1 U694 ( .A(n604), .B(KEYINPUT42), .ZN(n781) );
  XOR2_X1 U695 ( .A(KEYINPUT48), .B(KEYINPUT68), .Z(n605) );
  AND2_X1 U696 ( .A1(n607), .A2(n775), .ZN(n608) );
  XOR2_X1 U697 ( .A(n611), .B(n358), .Z(n610) );
  NAND2_X1 U698 ( .A1(n610), .A2(n726), .ZN(n615) );
  XNOR2_X1 U699 ( .A(G227), .B(n611), .ZN(n612) );
  NAND2_X1 U700 ( .A1(n612), .A2(G900), .ZN(n613) );
  NAND2_X1 U701 ( .A1(G953), .A2(n613), .ZN(n614) );
  NAND2_X1 U702 ( .A1(n615), .A2(n614), .ZN(G72) );
  XNOR2_X1 U703 ( .A(n625), .B(KEYINPUT80), .ZN(n618) );
  AND2_X1 U704 ( .A1(n682), .A2(n685), .ZN(n617) );
  INV_X1 U705 ( .A(KEYINPUT65), .ZN(n619) );
  XNOR2_X1 U706 ( .A(n619), .B(KEYINPUT32), .ZN(n620) );
  NAND2_X1 U707 ( .A1(n622), .A2(KEYINPUT44), .ZN(n641) );
  AND2_X1 U708 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U709 ( .A1(n623), .A2(n626), .ZN(n627) );
  NOR2_X1 U710 ( .A1(n629), .A2(n632), .ZN(n694) );
  NAND2_X1 U711 ( .A1(n635), .A2(n694), .ZN(n631) );
  INV_X1 U712 ( .A(KEYINPUT31), .ZN(n630) );
  INV_X1 U713 ( .A(n632), .ZN(n692) );
  NOR2_X1 U714 ( .A1(n692), .A2(n633), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n760) );
  NAND2_X1 U716 ( .A1(n771), .A2(n760), .ZN(n637) );
  NAND2_X1 U717 ( .A1(n637), .A2(n636), .ZN(n639) );
  INV_X1 U718 ( .A(KEYINPUT108), .ZN(n638) );
  NAND2_X1 U719 ( .A1(n641), .A2(n640), .ZN(n643) );
  XNOR2_X1 U720 ( .A(n643), .B(n642), .ZN(n648) );
  INV_X1 U721 ( .A(KEYINPUT44), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X2 U723 ( .A(n649), .B(KEYINPUT45), .ZN(n675) );
  NAND2_X1 U724 ( .A1(n675), .A2(n650), .ZN(n651) );
  XNOR2_X1 U725 ( .A(n651), .B(KEYINPUT89), .ZN(n652) );
  NAND2_X1 U726 ( .A1(n652), .A2(n358), .ZN(n656) );
  INV_X1 U727 ( .A(KEYINPUT2), .ZN(n653) );
  OR2_X1 U728 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U729 ( .A1(n656), .A2(n655), .ZN(n662) );
  INV_X1 U730 ( .A(KEYINPUT90), .ZN(n657) );
  XNOR2_X1 U731 ( .A(n658), .B(n657), .ZN(n659) );
  BUF_X2 U732 ( .A(n675), .Z(n727) );
  NAND2_X1 U733 ( .A1(n659), .A2(n727), .ZN(n661) );
  INV_X1 U734 ( .A(KEYINPUT77), .ZN(n660) );
  XNOR2_X2 U735 ( .A(n661), .B(n660), .ZN(n681) );
  NAND2_X1 U736 ( .A1(n739), .A2(G472), .ZN(n667) );
  XNOR2_X1 U737 ( .A(KEYINPUT94), .B(KEYINPUT114), .ZN(n663) );
  XNOR2_X1 U738 ( .A(n663), .B(KEYINPUT62), .ZN(n664) );
  XNOR2_X1 U739 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U740 ( .A(n667), .B(n666), .ZN(n671) );
  NAND2_X1 U741 ( .A1(n668), .A2(G953), .ZN(n670) );
  INV_X1 U742 ( .A(KEYINPUT96), .ZN(n669) );
  NOR2_X2 U743 ( .A1(n671), .A2(n778), .ZN(n673) );
  XNOR2_X1 U744 ( .A(KEYINPUT95), .B(KEYINPUT63), .ZN(n672) );
  XNOR2_X1 U745 ( .A(n673), .B(n672), .ZN(G57) );
  XNOR2_X1 U746 ( .A(n674), .B(G143), .ZN(G45) );
  NOR2_X1 U747 ( .A1(n675), .A2(KEYINPUT2), .ZN(n676) );
  XNOR2_X1 U748 ( .A(n676), .B(KEYINPUT88), .ZN(n678) );
  NOR2_X1 U749 ( .A1(n358), .A2(KEYINPUT2), .ZN(n677) );
  XNOR2_X1 U750 ( .A(n679), .B(KEYINPUT82), .ZN(n680) );
  NOR2_X1 U751 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U752 ( .A(KEYINPUT50), .B(n684), .Z(n690) );
  NAND2_X1 U753 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U754 ( .A(n687), .B(KEYINPUT119), .ZN(n688) );
  XNOR2_X1 U755 ( .A(KEYINPUT49), .B(n688), .ZN(n689) );
  NAND2_X1 U756 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U757 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U758 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U759 ( .A(KEYINPUT51), .B(n695), .Z(n696) );
  NOR2_X1 U760 ( .A1(n710), .A2(n696), .ZN(n706) );
  NOR2_X1 U761 ( .A1(n697), .A2(n394), .ZN(n698) );
  NOR2_X1 U762 ( .A1(n699), .A2(n698), .ZN(n703) );
  NOR2_X1 U763 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U764 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U765 ( .A1(n711), .A2(n704), .ZN(n705) );
  NOR2_X1 U766 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U767 ( .A(n707), .B(KEYINPUT52), .ZN(n709) );
  NOR2_X1 U768 ( .A1(n709), .A2(n708), .ZN(n713) );
  NOR2_X1 U769 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U770 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U771 ( .A(G119), .B(KEYINPUT126), .ZN(n716) );
  XNOR2_X1 U772 ( .A(n717), .B(n716), .ZN(G21) );
  NAND2_X1 U773 ( .A1(n739), .A2(G210), .ZN(n722) );
  XOR2_X1 U774 ( .A(KEYINPUT84), .B(KEYINPUT54), .Z(n719) );
  XNOR2_X1 U775 ( .A(n719), .B(KEYINPUT55), .ZN(n720) );
  XNOR2_X1 U776 ( .A(n718), .B(n720), .ZN(n721) );
  XNOR2_X1 U777 ( .A(n722), .B(n721), .ZN(n723) );
  NOR2_X2 U778 ( .A1(n723), .A2(n778), .ZN(n725) );
  XOR2_X1 U779 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n724) );
  XNOR2_X1 U780 ( .A(n725), .B(n724), .ZN(G51) );
  NAND2_X1 U781 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U782 ( .A(KEYINPUT124), .B(n728), .Z(n732) );
  NAND2_X1 U783 ( .A1(G953), .A2(G224), .ZN(n729) );
  XOR2_X1 U784 ( .A(KEYINPUT61), .B(n729), .Z(n730) );
  NOR2_X1 U785 ( .A1(n734), .A2(n730), .ZN(n731) );
  NOR2_X1 U786 ( .A1(n732), .A2(n731), .ZN(n738) );
  INV_X1 U787 ( .A(n733), .ZN(n736) );
  NAND2_X1 U788 ( .A1(n734), .A2(G953), .ZN(n735) );
  NAND2_X1 U789 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U790 ( .A(n738), .B(n737), .ZN(G69) );
  NAND2_X1 U791 ( .A1(n751), .A2(G217), .ZN(n742) );
  XNOR2_X1 U792 ( .A(n740), .B(KEYINPUT123), .ZN(n741) );
  XNOR2_X1 U793 ( .A(n742), .B(n741), .ZN(n743) );
  NOR2_X1 U794 ( .A1(n743), .A2(n778), .ZN(G66) );
  XNOR2_X1 U795 ( .A(n745), .B(KEYINPUT59), .ZN(n746) );
  XNOR2_X1 U796 ( .A(n747), .B(n746), .ZN(n748) );
  NOR2_X1 U797 ( .A1(n748), .A2(n778), .ZN(n750) );
  XNOR2_X1 U798 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n749) );
  XNOR2_X1 U799 ( .A(n750), .B(n749), .ZN(G60) );
  NAND2_X1 U800 ( .A1(n751), .A2(G469), .ZN(n755) );
  XOR2_X1 U801 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n752) );
  XNOR2_X1 U802 ( .A(n753), .B(n752), .ZN(n754) );
  XNOR2_X1 U803 ( .A(n755), .B(n754), .ZN(n756) );
  NOR2_X1 U804 ( .A1(n756), .A2(n778), .ZN(G54) );
  NOR2_X1 U805 ( .A1(n760), .A2(n769), .ZN(n757) );
  XOR2_X1 U806 ( .A(G104), .B(n757), .Z(G6) );
  XOR2_X1 U807 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n759) );
  XNOR2_X1 U808 ( .A(G107), .B(KEYINPUT116), .ZN(n758) );
  XNOR2_X1 U809 ( .A(n759), .B(n758), .ZN(n762) );
  INV_X1 U810 ( .A(n763), .ZN(n772) );
  NOR2_X1 U811 ( .A1(n760), .A2(n772), .ZN(n761) );
  XOR2_X1 U812 ( .A(n762), .B(n761), .Z(G9) );
  XOR2_X1 U813 ( .A(G128), .B(KEYINPUT29), .Z(n765) );
  NAND2_X1 U814 ( .A1(n767), .A2(n763), .ZN(n764) );
  XNOR2_X1 U815 ( .A(n765), .B(n764), .ZN(G30) );
  NAND2_X1 U816 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U817 ( .A(n768), .B(G146), .ZN(G48) );
  NOR2_X1 U818 ( .A1(n769), .A2(n771), .ZN(n770) );
  XOR2_X1 U819 ( .A(G113), .B(n770), .Z(G15) );
  NOR2_X1 U820 ( .A1(n772), .A2(n771), .ZN(n774) );
  XNOR2_X1 U821 ( .A(G116), .B(KEYINPUT117), .ZN(n773) );
  XNOR2_X1 U822 ( .A(n774), .B(n773), .ZN(G18) );
  XNOR2_X1 U823 ( .A(G134), .B(n775), .ZN(G36) );
  XNOR2_X1 U824 ( .A(n356), .B(n776), .ZN(n777) );
  NOR2_X1 U825 ( .A1(n778), .A2(n777), .ZN(G63) );
  XNOR2_X1 U826 ( .A(G101), .B(n779), .ZN(n780) );
  XNOR2_X1 U827 ( .A(n780), .B(KEYINPUT115), .ZN(G3) );
  XOR2_X1 U828 ( .A(G137), .B(n781), .Z(G39) );
  XOR2_X1 U829 ( .A(n782), .B(G131), .Z(G33) );
  XNOR2_X1 U830 ( .A(n783), .B(KEYINPUT37), .ZN(n784) );
  XNOR2_X1 U831 ( .A(G125), .B(n784), .ZN(G27) );
endmodule

