//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981;
  INV_X1    g000(.A(KEYINPUT18), .ZN(new_n202));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203));
  INV_X1    g002(.A(KEYINPUT15), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  INV_X1    g005(.A(G36gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT14), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT14), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n209), .B1(G29gat), .B2(G36gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n205), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT86), .B(G36gat), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n203), .A2(new_n204), .B1(new_n213), .B2(G29gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT85), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n208), .A2(new_n210), .A3(KEYINPUT85), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n213), .A2(G29gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(new_n205), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n215), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT17), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n212), .A2(new_n214), .B1(new_n220), .B2(new_n205), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT17), .ZN(new_n226));
  XNOR2_X1  g025(.A(G15gat), .B(G22gat), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n227), .A2(G1gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT87), .ZN(new_n229));
  AOI21_X1  g028(.A(G8gat), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT16), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n227), .B1(new_n231), .B2(G1gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n228), .B(new_n232), .C1(new_n229), .C2(G8gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n224), .A2(new_n226), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n222), .A2(new_n235), .A3(new_n234), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G229gat), .A2(G233gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n202), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n237), .A2(KEYINPUT18), .A3(new_n240), .A4(new_n238), .ZN(new_n243));
  XOR2_X1   g042(.A(new_n240), .B(KEYINPUT13), .Z(new_n244));
  INV_X1    g043(.A(new_n238), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n222), .B1(new_n235), .B2(new_n234), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n242), .A2(new_n243), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G113gat), .B(G141gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(G197gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT11), .B(G169gat), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n250), .B(new_n251), .Z(new_n252));
  XOR2_X1   g051(.A(new_n252), .B(KEYINPUT12), .Z(new_n253));
  NAND2_X1  g052(.A1(new_n248), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n253), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n242), .A2(new_n255), .A3(new_n243), .A4(new_n247), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(G225gat), .A2(G233gat), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G155gat), .A2(G162gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT2), .ZN(new_n262));
  OR2_X1    g061(.A1(G141gat), .A2(G148gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(G141gat), .A2(G148gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT75), .ZN(new_n266));
  AND2_X1   g065(.A1(G155gat), .A2(G162gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G155gat), .ZN(new_n270));
  INV_X1    g069(.A(G162gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(KEYINPUT75), .A3(new_n261), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n265), .A2(new_n269), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n262), .A2(KEYINPUT76), .ZN(new_n275));
  AND2_X1   g074(.A1(G141gat), .A2(G148gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(G141gat), .A2(G148gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G155gat), .B(G162gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT76), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n261), .A2(new_n280), .A3(KEYINPUT2), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n275), .A2(new_n278), .A3(new_n279), .A4(new_n281), .ZN(new_n282));
  AND2_X1   g081(.A1(new_n274), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n284));
  AND2_X1   g083(.A1(KEYINPUT71), .A2(G113gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(KEYINPUT71), .A2(G113gat), .ZN(new_n286));
  INV_X1    g085(.A(G120gat), .ZN(new_n287));
  NOR3_X1   g086(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(G113gat), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n284), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n292));
  INV_X1    g091(.A(G113gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(KEYINPUT71), .A2(G113gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(G120gat), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n296), .A2(KEYINPUT72), .A3(new_n289), .ZN(new_n297));
  INV_X1    g096(.A(G134gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G127gat), .ZN(new_n299));
  INV_X1    g098(.A(G127gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G134gat), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT1), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n299), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n291), .A2(new_n297), .A3(new_n304), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n299), .A2(new_n301), .A3(KEYINPUT70), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n293), .A2(G120gat), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT1), .B1(new_n289), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n299), .A2(KEYINPUT70), .ZN(new_n309));
  NOR3_X1   g108(.A1(new_n306), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n283), .A2(new_n305), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n274), .A2(new_n282), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT3), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT3), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n274), .A2(new_n282), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n296), .A2(new_n289), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n303), .B1(new_n318), .B2(new_n284), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n310), .B1(new_n319), .B2(new_n297), .ZN(new_n320));
  OAI211_X1 g119(.A(KEYINPUT4), .B(new_n312), .C1(new_n317), .C2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT4), .ZN(new_n322));
  AND4_X1   g121(.A1(new_n322), .A2(new_n283), .A3(new_n305), .A4(new_n311), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n260), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n283), .A2(new_n305), .A3(new_n311), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n283), .B1(new_n311), .B2(new_n305), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n260), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT5), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT77), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT5), .ZN(new_n331));
  AND3_X1   g130(.A1(new_n296), .A2(KEYINPUT72), .A3(new_n289), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT72), .B1(new_n296), .B2(new_n289), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n332), .A2(new_n333), .A3(new_n303), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n313), .B1(new_n334), .B2(new_n310), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(new_n312), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n331), .B1(new_n336), .B2(new_n260), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT77), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n322), .B1(new_n320), .B2(new_n283), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n305), .A2(new_n311), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n340), .A2(new_n316), .A3(new_n314), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n323), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n337), .B(new_n338), .C1(new_n342), .C2(new_n260), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n325), .A2(new_n331), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n330), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n346), .B(KEYINPUT79), .ZN(new_n347));
  XOR2_X1   g146(.A(G1gat), .B(G29gat), .Z(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G57gat), .B(G85gat), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n349), .B(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n345), .A2(KEYINPUT6), .A3(new_n353), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n345), .A2(new_n353), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n330), .A2(new_n343), .A3(new_n352), .A4(new_n344), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT6), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n354), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G8gat), .B(G36gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(G64gat), .B(G92gat), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n360), .B(new_n361), .Z(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G183gat), .A2(G190gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(G169gat), .A2(G176gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n365), .B(KEYINPUT26), .ZN(new_n366));
  NAND2_X1  g165(.A1(G169gat), .A2(G176gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT66), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT66), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(G169gat), .A3(G176gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT27), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(G183gat), .ZN(new_n374));
  INV_X1    g173(.A(G183gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT27), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT69), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n374), .A2(new_n376), .A3(KEYINPUT69), .ZN(new_n380));
  INV_X1    g179(.A(G190gat), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n381), .A2(KEYINPUT28), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n379), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT68), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n377), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(G190gat), .B1(new_n374), .B2(KEYINPUT68), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT28), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n364), .B(new_n372), .C1(new_n383), .C2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n364), .A2(KEYINPUT24), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT24), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(G183gat), .A3(G190gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n392), .B1(G183gat), .B2(G190gat), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT23), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n365), .A2(new_n395), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n394), .A2(new_n396), .B1(new_n368), .B2(new_n370), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n393), .A2(KEYINPUT25), .A3(new_n397), .ZN(new_n398));
  XOR2_X1   g197(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n399));
  OAI21_X1  g198(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n400));
  OR3_X1    g199(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n392), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n399), .B1(new_n402), .B2(new_n397), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT67), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n398), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI211_X1 g204(.A(KEYINPUT67), .B(new_n399), .C1(new_n402), .C2(new_n397), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n388), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(G226gat), .A2(G233gat), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT29), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G197gat), .B(G204gat), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT22), .ZN(new_n414));
  INV_X1    g213(.A(G211gat), .ZN(new_n415));
  INV_X1    g214(.A(G218gat), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  XOR2_X1   g217(.A(G211gat), .B(G218gat), .Z(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n388), .B(new_n409), .C1(new_n405), .C2(new_n406), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n412), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n420), .B1(new_n412), .B2(new_n421), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n363), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n412), .A2(new_n421), .ZN(new_n425));
  INV_X1    g224(.A(new_n420), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n412), .A2(new_n420), .A3(new_n421), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n428), .A3(new_n362), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n424), .A2(new_n429), .A3(KEYINPUT30), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT30), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n427), .A2(new_n431), .A3(new_n428), .A4(new_n362), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n359), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n420), .B1(new_n410), .B2(new_n316), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n410), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n315), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n435), .B1(new_n437), .B2(new_n313), .ZN(new_n438));
  XNOR2_X1  g237(.A(G78gat), .B(G106gat), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n438), .B(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT80), .ZN(new_n442));
  INV_X1    g241(.A(G228gat), .ZN(new_n443));
  INV_X1    g242(.A(G233gat), .ZN(new_n444));
  OAI22_X1  g243(.A1(new_n435), .A2(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(G22gat), .ZN(new_n446));
  INV_X1    g245(.A(G22gat), .ZN(new_n447));
  OAI221_X1 g246(.A(new_n447), .B1(new_n443), .B2(new_n444), .C1(new_n435), .C2(new_n442), .ZN(new_n448));
  XNOR2_X1  g247(.A(KEYINPUT31), .B(G50gat), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n446), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n450), .B1(new_n446), .B2(new_n448), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n441), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n446), .A2(new_n448), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n449), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n438), .B(new_n439), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n446), .A2(new_n448), .A3(new_n450), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT81), .B1(new_n453), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n453), .A2(new_n458), .A3(KEYINPUT81), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n434), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT36), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n407), .A2(new_n320), .ZN(new_n465));
  AND2_X1   g264(.A1(G227gat), .A2(G233gat), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n388), .B(new_n340), .C1(new_n405), .C2(new_n406), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  XOR2_X1   g267(.A(G71gat), .B(G99gat), .Z(new_n469));
  XNOR2_X1  g268(.A(G15gat), .B(G43gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT33), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n468), .A2(KEYINPUT32), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT73), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n468), .A2(KEYINPUT73), .A3(KEYINPUT32), .A4(new_n472), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n468), .A2(KEYINPUT32), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT33), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n468), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n480), .A3(new_n471), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n466), .B1(new_n465), .B2(new_n467), .ZN(new_n482));
  XOR2_X1   g281(.A(KEYINPUT74), .B(KEYINPUT34), .Z(new_n483));
  OR2_X1    g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT74), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n482), .A2(new_n485), .A3(KEYINPUT34), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n477), .A2(new_n481), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n487), .B1(new_n477), .B2(new_n481), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n464), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n477), .A2(new_n481), .ZN(new_n491));
  INV_X1    g290(.A(new_n487), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n481), .A3(new_n487), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(KEYINPUT36), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n427), .A2(new_n428), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n363), .B1(new_n497), .B2(KEYINPUT37), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT37), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n499), .B1(new_n427), .B2(new_n428), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT38), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n424), .B1(new_n499), .B2(new_n362), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT38), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n499), .B1(new_n422), .B2(KEYINPUT84), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT84), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n427), .A2(new_n505), .A3(new_n428), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n502), .A2(new_n503), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n501), .A2(new_n508), .A3(new_n429), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n352), .B1(new_n345), .B2(KEYINPUT83), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT83), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n330), .A2(new_n343), .A3(new_n511), .A4(new_n344), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n358), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n354), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n509), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n430), .A2(new_n432), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n345), .A2(KEYINPUT83), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(new_n353), .A3(new_n512), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n342), .A2(new_n260), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n519), .B(KEYINPUT39), .C1(new_n260), .C2(new_n336), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT39), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n321), .A2(new_n324), .A3(new_n521), .A4(new_n260), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT82), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n522), .A2(new_n523), .A3(new_n352), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n523), .B1(new_n522), .B2(new_n352), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n520), .B(KEYINPUT40), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n520), .B1(new_n524), .B2(new_n525), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT40), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n516), .A2(new_n518), .A3(new_n526), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n453), .A2(new_n458), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n463), .B(new_n496), .C1(new_n515), .C2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n358), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n354), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n453), .A2(new_n458), .ZN(new_n537));
  NOR3_X1   g336(.A1(new_n488), .A2(new_n489), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT35), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n536), .A2(new_n538), .A3(new_n539), .A4(new_n433), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n493), .A2(new_n531), .A3(new_n494), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT35), .B1(new_n434), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n258), .B1(new_n533), .B2(new_n543), .ZN(new_n544));
  AND2_X1   g343(.A1(G232gat), .A2(G233gat), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n545), .A2(KEYINPUT41), .ZN(new_n546));
  XNOR2_X1  g345(.A(G134gat), .B(G162gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(G85gat), .A2(G92gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT92), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n551), .A2(KEYINPUT7), .ZN(new_n552));
  NAND2_X1  g351(.A1(G85gat), .A2(G92gat), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(KEYINPUT7), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT7), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT92), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n555), .A2(new_n557), .A3(G85gat), .A4(G92gat), .ZN(new_n558));
  INV_X1    g357(.A(G99gat), .ZN(new_n559));
  INV_X1    g358(.A(G106gat), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT8), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n554), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(G99gat), .B(G106gat), .Z(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n563), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n565), .A2(new_n558), .A3(new_n561), .A4(new_n554), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n224), .A2(new_n226), .A3(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G190gat), .B(G218gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n569), .B(new_n570), .Z(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n567), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n222), .A2(new_n573), .B1(KEYINPUT41), .B2(new_n545), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n568), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n572), .B1(new_n568), .B2(new_n574), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n549), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n577), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n579), .A2(new_n548), .A3(new_n575), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G71gat), .B(G78gat), .Z(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n585));
  INV_X1    g384(.A(G57gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(G64gat), .ZN(new_n587));
  INV_X1    g386(.A(G64gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(G57gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT88), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n585), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n587), .A2(new_n589), .A3(KEYINPUT88), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n584), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT89), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n587), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n589), .B(KEYINPUT90), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n583), .A2(new_n585), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n594), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n600), .A2(KEYINPUT21), .ZN(new_n601));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n601), .B(new_n602), .Z(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(new_n300), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n598), .A2(new_n599), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n592), .A2(new_n593), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n605), .B1(new_n584), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT91), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT91), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n600), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n610), .A3(KEYINPUT21), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(new_n236), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n604), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n603), .B(G127gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(new_n612), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(new_n270), .ZN(new_n619));
  XNOR2_X1  g418(.A(G183gat), .B(G211gat), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n619), .B(new_n620), .Z(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n614), .A2(new_n616), .A3(new_n621), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n582), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT97), .ZN(new_n626));
  NAND2_X1  g425(.A1(G230gat), .A2(G233gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n567), .A2(KEYINPUT95), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT95), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n564), .A2(new_n629), .A3(new_n566), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n628), .A2(new_n607), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n600), .A2(KEYINPUT95), .A3(new_n567), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT10), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT10), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n567), .A2(new_n634), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n608), .A2(new_n610), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n627), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n627), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n631), .A2(new_n638), .A3(new_n632), .ZN(new_n639));
  XNOR2_X1  g438(.A(G120gat), .B(G148gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT96), .ZN(new_n641));
  XNOR2_X1  g440(.A(G176gat), .B(G204gat), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n641), .B(new_n642), .Z(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n637), .A2(new_n639), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n644), .B1(new_n637), .B2(new_n639), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n626), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n647), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n649), .A2(KEYINPUT97), .A3(new_n645), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n544), .A2(new_n625), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n359), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g454(.A1(new_n652), .A2(new_n516), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n656), .A2(G8gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT16), .B(G8gat), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(KEYINPUT42), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n660), .B1(KEYINPUT42), .B2(new_n659), .ZN(G1325gat));
  INV_X1    g460(.A(G15gat), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n493), .A2(new_n494), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n652), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n496), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n652), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n665), .B1(new_n667), .B2(new_n662), .ZN(G1326gat));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n462), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT43), .B(G22gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  NAND2_X1  g470(.A1(new_n623), .A2(new_n624), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n673), .A2(new_n582), .A3(new_n651), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT98), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n675), .A2(new_n544), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n676), .A2(new_n206), .A3(new_n653), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT45), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n533), .A2(new_n543), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT44), .B1(new_n679), .B2(new_n581), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n496), .B1(new_n515), .B2(new_n532), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n345), .A2(new_n353), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n682), .A2(new_n357), .A3(new_n356), .ZN(new_n683));
  AOI22_X1  g482(.A1(new_n683), .A2(new_n354), .B1(new_n432), .B2(new_n430), .ZN(new_n684));
  INV_X1    g483(.A(new_n461), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(new_n459), .ZN(new_n686));
  OAI21_X1  g485(.A(KEYINPUT99), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT99), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n434), .A2(new_n688), .A3(new_n462), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n543), .B1(new_n681), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT100), .B(KEYINPUT44), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(new_n582), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n680), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n651), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n672), .A2(new_n258), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(G29gat), .B1(new_n697), .B2(new_n359), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n678), .A2(new_n698), .ZN(G1328gat));
  INV_X1    g498(.A(new_n213), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n676), .A2(new_n516), .A3(new_n700), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n701), .B(KEYINPUT46), .Z(new_n702));
  OAI21_X1  g501(.A(new_n213), .B1(new_n697), .B2(new_n433), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(G1329gat));
  OAI21_X1  g503(.A(G43gat), .B1(new_n697), .B2(new_n496), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT101), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT47), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(G43gat), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n676), .A2(new_n708), .A3(new_n664), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n707), .B(new_n710), .ZN(G1330gat));
  INV_X1    g510(.A(G50gat), .ZN(new_n712));
  AND3_X1   g511(.A1(new_n676), .A2(new_n712), .A3(new_n462), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT102), .ZN(new_n714));
  OAI21_X1  g513(.A(G50gat), .B1(new_n697), .B2(new_n531), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n713), .B1(KEYINPUT102), .B2(KEYINPUT48), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n712), .A2(KEYINPUT48), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n718), .B1(new_n697), .B2(new_n686), .ZN(new_n719));
  AOI22_X1  g518(.A1(new_n716), .A2(KEYINPUT48), .B1(new_n717), .B2(new_n719), .ZN(G1331gat));
  AND3_X1   g519(.A1(new_n625), .A2(new_n258), .A3(new_n695), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n691), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n653), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(G57gat), .ZN(G1332gat));
  INV_X1    g523(.A(new_n722), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(new_n433), .ZN(new_n726));
  NOR2_X1   g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  AND2_X1   g526(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n729), .B1(new_n726), .B2(new_n727), .ZN(G1333gat));
  NAND3_X1  g529(.A1(new_n722), .A2(G71gat), .A3(new_n666), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT103), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n725), .A2(new_n663), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(G71gat), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g534(.A1(new_n722), .A2(new_n462), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g536(.A1(new_n672), .A2(new_n257), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n695), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n739), .B1(new_n680), .B2(new_n693), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n740), .A2(G85gat), .A3(new_n653), .ZN(new_n741));
  INV_X1    g540(.A(new_n738), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n531), .B(new_n530), .C1(new_n536), .C2(new_n509), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n743), .A2(new_n496), .A3(new_n687), .A4(new_n689), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n581), .B1(new_n744), .B2(new_n543), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n742), .B1(new_n745), .B2(KEYINPUT104), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n691), .A2(new_n582), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT104), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n746), .A2(KEYINPUT51), .A3(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n691), .A2(KEYINPUT104), .A3(new_n582), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n738), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT104), .B1(new_n691), .B2(new_n582), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n753), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n750), .B2(new_n751), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n653), .B(new_n695), .C1(new_n752), .C2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(G85gat), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n741), .B1(new_n759), .B2(new_n760), .ZN(G1336gat));
  NOR2_X1   g560(.A1(new_n651), .A2(new_n433), .ZN(new_n762));
  INV_X1    g561(.A(G92gat), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n752), .B2(new_n758), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n740), .A2(new_n516), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G92gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n755), .A2(new_n753), .A3(new_n756), .ZN(new_n771));
  AOI21_X1  g570(.A(KEYINPUT51), .B1(new_n746), .B2(new_n749), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n765), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n769), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT106), .B1(new_n774), .B2(KEYINPUT52), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n764), .B1(new_n757), .B2(new_n750), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n763), .B1(new_n740), .B2(new_n516), .ZN(new_n777));
  OAI211_X1 g576(.A(KEYINPUT106), .B(KEYINPUT52), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n770), .B1(new_n775), .B2(new_n779), .ZN(G1337gat));
  NAND2_X1  g579(.A1(new_n740), .A2(new_n666), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT107), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n559), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n783), .B1(new_n782), .B2(new_n781), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n663), .A2(new_n651), .A3(G99gat), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(new_n752), .B2(new_n758), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(G1338gat));
  INV_X1    g586(.A(new_n739), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n694), .A2(new_n462), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G106gat), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT108), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n789), .A2(KEYINPUT108), .A3(G106gat), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n651), .A2(G106gat), .A3(new_n531), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT109), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(new_n771), .B2(new_n772), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n792), .A2(new_n793), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT53), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n740), .A2(new_n537), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n560), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n740), .A2(KEYINPUT110), .A3(new_n537), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT53), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n794), .B1(new_n752), .B2(new_n758), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n798), .A2(new_n805), .ZN(G1339gat));
  INV_X1    g605(.A(KEYINPUT113), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n608), .A2(new_n610), .A3(new_n635), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n631), .A2(new_n632), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n638), .B(new_n809), .C1(new_n810), .C2(KEYINPUT10), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n811), .A2(new_n637), .A3(KEYINPUT54), .ZN(new_n812));
  XOR2_X1   g611(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n813));
  OAI211_X1 g612(.A(new_n627), .B(new_n813), .C1(new_n633), .C2(new_n636), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n643), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n808), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n811), .A2(new_n637), .A3(KEYINPUT54), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n817), .A2(KEYINPUT55), .A3(new_n643), .A4(new_n814), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n816), .A2(new_n645), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n239), .A2(new_n241), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT112), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n245), .A2(new_n246), .ZN(new_n822));
  INV_X1    g621(.A(new_n244), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n820), .A2(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n239), .A2(KEYINPUT112), .A3(new_n241), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n252), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n827), .A2(new_n582), .A3(new_n256), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n807), .B1(new_n819), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n818), .A2(new_n645), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n252), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n832), .B1(new_n824), .B2(new_n825), .ZN(new_n833));
  AND4_X1   g632(.A1(new_n255), .A2(new_n242), .A3(new_n243), .A4(new_n247), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n833), .A2(new_n834), .A3(new_n581), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n831), .A2(new_n835), .A3(KEYINPUT113), .A4(new_n816), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n829), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n648), .A2(new_n650), .A3(new_n256), .A4(new_n827), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n816), .A2(new_n257), .A3(new_n645), .A4(new_n818), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n582), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n673), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n625), .A2(new_n258), .A3(new_n651), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n359), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n843), .A2(new_n433), .A3(new_n538), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n844), .A2(new_n294), .A3(new_n295), .A4(new_n257), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n462), .B1(new_n841), .B2(new_n842), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n653), .A2(new_n433), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(new_n663), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(G113gat), .B1(new_n849), .B2(new_n258), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n845), .A2(new_n850), .ZN(G1340gat));
  NAND3_X1  g650(.A1(new_n846), .A2(new_n695), .A3(new_n848), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(G120gat), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(KEYINPUT114), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n844), .A2(new_n287), .A3(new_n695), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT115), .ZN(G1341gat));
  NAND3_X1  g656(.A1(new_n844), .A2(new_n300), .A3(new_n672), .ZN(new_n858));
  OAI21_X1  g657(.A(G127gat), .B1(new_n849), .B2(new_n673), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1342gat));
  NAND3_X1  g659(.A1(new_n844), .A2(new_n298), .A3(new_n582), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n862));
  OAI21_X1  g661(.A(G134gat), .B1(new_n849), .B2(new_n581), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(G1343gat));
  INV_X1    g664(.A(KEYINPUT120), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT58), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n841), .A2(new_n842), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n666), .A2(new_n531), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n653), .A3(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n258), .A2(new_n516), .A3(G141gat), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n843), .A2(KEYINPUT118), .A3(new_n869), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT119), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n666), .A2(new_n847), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n531), .B1(new_n841), .B2(new_n842), .ZN(new_n878));
  XOR2_X1   g677(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n462), .A2(KEYINPUT57), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n883));
  INV_X1    g682(.A(new_n815), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT55), .B1(new_n884), .B2(new_n817), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n883), .B1(new_n830), .B2(new_n885), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n816), .A2(KEYINPUT117), .A3(new_n645), .A4(new_n818), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n257), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n582), .B1(new_n888), .B2(new_n838), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n673), .B1(new_n889), .B2(new_n837), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n882), .B1(new_n890), .B2(new_n842), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n257), .B(new_n877), .C1(new_n881), .C2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(G141gat), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n872), .A2(new_n894), .A3(new_n873), .A4(new_n874), .ZN(new_n895));
  AND4_X1   g694(.A1(new_n867), .A2(new_n876), .A3(new_n893), .A4(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n843), .A2(new_n869), .A3(new_n873), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n867), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n866), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n898), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n876), .A2(new_n893), .A3(new_n867), .A4(new_n895), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n900), .A2(KEYINPUT120), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n899), .A2(new_n902), .ZN(G1344gat));
  INV_X1    g702(.A(new_n877), .ZN(new_n904));
  INV_X1    g703(.A(new_n881), .ZN(new_n905));
  INV_X1    g704(.A(new_n891), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n695), .ZN(new_n908));
  AOI21_X1  g707(.A(KEYINPUT59), .B1(new_n908), .B2(G148gat), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n872), .A2(new_n433), .A3(new_n874), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n651), .A2(G148gat), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n819), .A2(new_n828), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n673), .B1(new_n889), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n842), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n915), .A2(KEYINPUT121), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n686), .B1(new_n915), .B2(KEYINPUT121), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT57), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n878), .A2(new_n880), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n877), .A2(new_n695), .ZN(new_n921));
  OAI211_X1 g720(.A(KEYINPUT59), .B(G148gat), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n912), .A2(new_n922), .ZN(G1345gat));
  AOI21_X1  g722(.A(G155gat), .B1(new_n910), .B2(new_n672), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n672), .A2(G155gat), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT122), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n924), .B1(new_n907), .B2(new_n926), .ZN(G1346gat));
  NAND2_X1  g726(.A1(new_n907), .A2(new_n582), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT123), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n271), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n930), .B1(new_n929), .B2(new_n928), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n910), .A2(new_n271), .A3(new_n582), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1347gat));
  NAND2_X1  g732(.A1(new_n359), .A2(new_n516), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT124), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n935), .A2(new_n663), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n846), .A2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(G169gat), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n937), .A2(new_n938), .A3(new_n258), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n653), .B1(new_n841), .B2(new_n842), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(new_n538), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n941), .A2(new_n433), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(new_n257), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n939), .B1(new_n943), .B2(new_n938), .ZN(G1348gat));
  OAI21_X1  g743(.A(G176gat), .B1(new_n937), .B2(new_n651), .ZN(new_n945));
  INV_X1    g744(.A(G176gat), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n762), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n945), .B1(new_n941), .B2(new_n947), .ZN(G1349gat));
  NAND4_X1  g747(.A1(new_n942), .A2(new_n379), .A3(new_n380), .A4(new_n672), .ZN(new_n949));
  OAI21_X1  g748(.A(G183gat), .B1(new_n937), .B2(new_n673), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g750(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n951), .B(new_n952), .ZN(G1350gat));
  NAND3_X1  g752(.A1(new_n942), .A2(new_n381), .A3(new_n582), .ZN(new_n954));
  XNOR2_X1  g753(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n846), .A2(new_n582), .A3(new_n936), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n955), .B1(new_n956), .B2(G190gat), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n956), .A2(G190gat), .A3(new_n955), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n954), .B1(new_n957), .B2(new_n958), .ZN(G1351gat));
  AND3_X1   g758(.A1(new_n940), .A2(new_n516), .A3(new_n869), .ZN(new_n960));
  AOI21_X1  g759(.A(G197gat), .B1(new_n960), .B2(new_n257), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n920), .A2(new_n666), .A3(new_n935), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n257), .A2(G197gat), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(G1352gat));
  OR2_X1    g763(.A1(new_n918), .A2(new_n919), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n935), .A2(new_n666), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n965), .A2(new_n695), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(G204gat), .ZN(new_n968));
  INV_X1    g767(.A(G204gat), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n960), .A2(new_n969), .A3(new_n695), .ZN(new_n970));
  XOR2_X1   g769(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n971));
  XNOR2_X1  g770(.A(new_n970), .B(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n968), .A2(new_n972), .ZN(G1353gat));
  NAND3_X1  g772(.A1(new_n960), .A2(new_n415), .A3(new_n672), .ZN(new_n974));
  OAI211_X1 g773(.A(new_n672), .B(new_n966), .C1(new_n918), .C2(new_n919), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n975), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n976));
  AOI21_X1  g775(.A(KEYINPUT63), .B1(new_n975), .B2(G211gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(G1354gat));
  NAND3_X1  g777(.A1(new_n965), .A2(new_n582), .A3(new_n966), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(G218gat), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n960), .A2(new_n416), .A3(new_n582), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(G1355gat));
endmodule


