

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777;

  BUF_X1 U378 ( .A(n723), .Z(n356) );
  AND2_X1 U379 ( .A1(n589), .A2(n533), .ZN(n479) );
  OR2_X1 U380 ( .A1(n680), .A2(G902), .ZN(n466) );
  XNOR2_X1 U381 ( .A(n452), .B(n451), .ZN(n645) );
  XNOR2_X2 U382 ( .A(n593), .B(n426), .ZN(n580) );
  INV_X1 U383 ( .A(G953), .ZN(n760) );
  NOR2_X1 U384 ( .A1(G953), .A2(G237), .ZN(n496) );
  XOR2_X2 U385 ( .A(KEYINPUT90), .B(KEYINPUT0), .Z(n434) );
  XNOR2_X2 U386 ( .A(KEYINPUT74), .B(KEYINPUT22), .ZN(n516) );
  AND2_X2 U387 ( .A1(n479), .A2(n597), .ZN(n480) );
  XNOR2_X2 U388 ( .A(n416), .B(n766), .ZN(n436) );
  XNOR2_X2 U389 ( .A(n528), .B(n527), .ZN(n544) );
  INV_X1 U390 ( .A(KEYINPUT10), .ZN(n450) );
  INV_X1 U391 ( .A(G101), .ZN(n766) );
  OR2_X1 U392 ( .A1(n540), .A2(n542), .ZN(n382) );
  NOR2_X2 U393 ( .A1(n540), .A2(n364), .ZN(n528) );
  XNOR2_X2 U394 ( .A(n517), .B(n516), .ZN(n540) );
  AND2_X2 U395 ( .A1(n375), .A2(n376), .ZN(n374) );
  AND2_X2 U396 ( .A1(n361), .A2(n385), .ZN(n360) );
  NAND2_X2 U397 ( .A1(n360), .A2(n358), .ZN(n593) );
  NOR2_X1 U398 ( .A1(n379), .A2(n380), .ZN(n373) );
  INV_X1 U399 ( .A(n383), .ZN(n380) );
  XNOR2_X1 U400 ( .A(n532), .B(KEYINPUT31), .ZN(n705) );
  INV_X1 U401 ( .A(n530), .ZN(n357) );
  NAND2_X1 U402 ( .A1(n359), .A2(n365), .ZN(n358) );
  NOR2_X1 U403 ( .A1(n737), .A2(KEYINPUT89), .ZN(n365) );
  INV_X1 U404 ( .A(G237), .ZN(n421) );
  NAND2_X1 U405 ( .A1(G234), .A2(G237), .ZN(n427) );
  INV_X1 U406 ( .A(n554), .ZN(n359) );
  NAND2_X1 U407 ( .A1(n554), .A2(KEYINPUT89), .ZN(n361) );
  XNOR2_X2 U408 ( .A(n424), .B(n423), .ZN(n554) );
  NAND2_X1 U409 ( .A1(n644), .A2(n777), .ZN(n392) );
  XNOR2_X1 U410 ( .A(G110), .B(G107), .ZN(n417) );
  XNOR2_X1 U411 ( .A(KEYINPUT70), .B(G131), .ZN(n504) );
  NAND2_X1 U412 ( .A1(n362), .A2(n617), .ZN(n401) );
  NAND2_X1 U413 ( .A1(n362), .A2(KEYINPUT85), .ZN(n404) );
  XNOR2_X1 U414 ( .A(G137), .B(KEYINPUT71), .ZN(n475) );
  XNOR2_X1 U415 ( .A(n392), .B(n391), .ZN(n390) );
  XNOR2_X1 U416 ( .A(n418), .B(n767), .ZN(n474) );
  XNOR2_X1 U417 ( .A(n393), .B(KEYINPUT39), .ZN(n609) );
  NAND2_X1 U418 ( .A1(n382), .A2(n381), .ZN(n379) );
  INV_X1 U419 ( .A(KEYINPUT46), .ZN(n391) );
  NAND2_X1 U420 ( .A1(n737), .A2(KEYINPUT89), .ZN(n385) );
  XNOR2_X1 U421 ( .A(G113), .B(G122), .ZN(n499) );
  XNOR2_X1 U422 ( .A(G143), .B(G104), .ZN(n503) );
  INV_X1 U423 ( .A(G902), .ZN(n508) );
  XNOR2_X1 U424 ( .A(KEYINPUT95), .B(KEYINPUT5), .ZN(n441) );
  XNOR2_X1 U425 ( .A(n437), .B(n414), .ZN(n769) );
  XNOR2_X1 U426 ( .A(KEYINPUT16), .B(G122), .ZN(n414) );
  XNOR2_X1 U427 ( .A(G119), .B(KEYINPUT23), .ZN(n457) );
  XNOR2_X1 U428 ( .A(G128), .B(G110), .ZN(n458) );
  XNOR2_X1 U429 ( .A(KEYINPUT24), .B(KEYINPUT72), .ZN(n456) );
  XNOR2_X1 U430 ( .A(G116), .B(G107), .ZN(n482) );
  NAND2_X1 U431 ( .A1(n401), .A2(n400), .ZN(n399) );
  NAND2_X1 U432 ( .A1(KEYINPUT64), .A2(KEYINPUT85), .ZN(n400) );
  NAND2_X1 U433 ( .A1(n404), .A2(n403), .ZN(n402) );
  NAND2_X1 U434 ( .A1(n617), .A2(KEYINPUT64), .ZN(n403) );
  NOR2_X1 U435 ( .A1(n629), .A2(n628), .ZN(n712) );
  BUF_X1 U436 ( .A(n707), .Z(n746) );
  INV_X1 U437 ( .A(KEYINPUT32), .ZN(n527) );
  XNOR2_X1 U438 ( .A(n394), .B(KEYINPUT75), .ZN(n600) );
  NAND2_X1 U439 ( .A1(n395), .A2(n363), .ZN(n394) );
  OR2_X1 U440 ( .A1(n628), .A2(n396), .ZN(n764) );
  XOR2_X1 U441 ( .A(n630), .B(KEYINPUT59), .Z(n631) );
  XNOR2_X1 U442 ( .A(G146), .B(G140), .ZN(n473) );
  XNOR2_X1 U443 ( .A(n576), .B(KEYINPUT40), .ZN(n644) );
  BUF_X1 U444 ( .A(n544), .Z(n675) );
  NAND2_X1 U445 ( .A1(n357), .A2(n371), .ZN(n532) );
  INV_X1 U446 ( .A(n730), .ZN(n371) );
  BUF_X1 U447 ( .A(n545), .Z(n642) );
  INV_X1 U448 ( .A(n382), .ZN(n640) );
  INV_X1 U449 ( .A(n760), .ZN(n396) );
  NAND2_X1 U450 ( .A1(n620), .A2(KEYINPUT64), .ZN(n362) );
  AND2_X1 U451 ( .A1(n574), .A2(n573), .ZN(n363) );
  XNOR2_X1 U452 ( .A(KEYINPUT78), .B(n526), .ZN(n364) );
  AND2_X1 U453 ( .A1(n714), .A2(n402), .ZN(n366) );
  XOR2_X1 U454 ( .A(KEYINPUT65), .B(KEYINPUT1), .Z(n367) );
  XNOR2_X1 U455 ( .A(KEYINPUT106), .B(KEYINPUT33), .ZN(n368) );
  NOR2_X1 U456 ( .A1(n620), .A2(KEYINPUT64), .ZN(n369) );
  AND2_X1 U457 ( .A1(KEYINPUT44), .A2(KEYINPUT88), .ZN(n370) );
  NOR2_X1 U458 ( .A1(n712), .A2(n369), .ZN(n397) );
  AND2_X2 U459 ( .A1(n398), .A2(n397), .ZN(n678) );
  INV_X2 U460 ( .A(n518), .ZN(n570) );
  XNOR2_X1 U461 ( .A(n435), .B(n434), .ZN(n530) );
  NAND2_X1 U462 ( .A1(n374), .A2(n372), .ZN(n550) );
  NAND2_X1 U463 ( .A1(n373), .A2(n378), .ZN(n372) );
  NAND2_X1 U464 ( .A1(n384), .A2(n370), .ZN(n375) );
  NAND2_X1 U465 ( .A1(n377), .A2(KEYINPUT88), .ZN(n376) );
  NAND2_X1 U466 ( .A1(n382), .A2(n383), .ZN(n377) );
  OR2_X2 U467 ( .A1(n539), .A2(n577), .ZN(n383) );
  NAND2_X1 U468 ( .A1(n384), .A2(KEYINPUT44), .ZN(n378) );
  INV_X1 U469 ( .A(KEYINPUT88), .ZN(n381) );
  NAND2_X1 U470 ( .A1(n529), .A2(n544), .ZN(n384) );
  NAND2_X1 U471 ( .A1(n387), .A2(n386), .ZN(n398) );
  NAND2_X1 U472 ( .A1(n389), .A2(n366), .ZN(n386) );
  NAND2_X1 U473 ( .A1(n388), .A2(n399), .ZN(n387) );
  NAND2_X1 U474 ( .A1(n389), .A2(n714), .ZN(n388) );
  XNOR2_X1 U475 ( .A(n553), .B(KEYINPUT86), .ZN(n389) );
  NAND2_X1 U476 ( .A1(n390), .A2(n606), .ZN(n607) );
  NAND2_X1 U477 ( .A1(n600), .A2(n736), .ZN(n393) );
  INV_X1 U478 ( .A(n575), .ZN(n395) );
  BUF_X1 U479 ( .A(n678), .Z(n682) );
  XNOR2_X2 U480 ( .A(G143), .B(G128), .ZN(n445) );
  XOR2_X1 U481 ( .A(n473), .B(n472), .Z(n405) );
  INV_X1 U482 ( .A(n589), .ZN(n523) );
  INV_X1 U483 ( .A(KEYINPUT85), .ZN(n617) );
  XNOR2_X1 U484 ( .A(n474), .B(n405), .ZN(n477) );
  BUF_X1 U485 ( .A(n518), .Z(n726) );
  BUF_X1 U486 ( .A(n676), .Z(n677) );
  INV_X1 U487 ( .A(G953), .ZN(n406) );
  NAND2_X1 U488 ( .A1(n406), .A2(G224), .ZN(n407) );
  XNOR2_X1 U489 ( .A(n407), .B(KEYINPUT92), .ZN(n408) );
  XNOR2_X1 U490 ( .A(n408), .B(n445), .ZN(n411) );
  XNOR2_X2 U491 ( .A(G146), .B(G125), .ZN(n452) );
  XNOR2_X1 U492 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n409) );
  XNOR2_X1 U493 ( .A(n452), .B(n409), .ZN(n410) );
  XNOR2_X1 U494 ( .A(n411), .B(n410), .ZN(n415) );
  XNOR2_X2 U495 ( .A(G116), .B(G113), .ZN(n413) );
  XNOR2_X2 U496 ( .A(KEYINPUT3), .B(G119), .ZN(n412) );
  XNOR2_X2 U497 ( .A(n413), .B(n412), .ZN(n437) );
  XNOR2_X1 U498 ( .A(n415), .B(n769), .ZN(n419) );
  XNOR2_X2 U499 ( .A(KEYINPUT66), .B(KEYINPUT4), .ZN(n416) );
  XNOR2_X1 U500 ( .A(n436), .B(KEYINPUT73), .ZN(n418) );
  XNOR2_X1 U501 ( .A(n417), .B(G104), .ZN(n767) );
  XNOR2_X1 U502 ( .A(n419), .B(n474), .ZN(n665) );
  INV_X1 U503 ( .A(KEYINPUT15), .ZN(n420) );
  XNOR2_X1 U504 ( .A(n420), .B(G902), .ZN(n618) );
  OR2_X2 U505 ( .A1(n665), .A2(n618), .ZN(n424) );
  NAND2_X1 U506 ( .A1(n508), .A2(n421), .ZN(n425) );
  NAND2_X1 U507 ( .A1(n425), .A2(G210), .ZN(n422) );
  XNOR2_X1 U508 ( .A(n422), .B(KEYINPUT80), .ZN(n423) );
  AND2_X1 U509 ( .A1(n425), .A2(G214), .ZN(n737) );
  XNOR2_X1 U510 ( .A(KEYINPUT76), .B(KEYINPUT19), .ZN(n426) );
  XNOR2_X1 U511 ( .A(n427), .B(KEYINPUT14), .ZN(n430) );
  NAND2_X1 U512 ( .A1(G952), .A2(n430), .ZN(n753) );
  NOR2_X1 U513 ( .A1(n753), .A2(n396), .ZN(n429) );
  INV_X1 U514 ( .A(KEYINPUT93), .ZN(n428) );
  XNOR2_X1 U515 ( .A(n429), .B(n428), .ZN(n561) );
  NAND2_X1 U516 ( .A1(G902), .A2(n430), .ZN(n558) );
  INV_X1 U517 ( .A(G898), .ZN(n431) );
  NAND2_X1 U518 ( .A1(n431), .A2(n396), .ZN(n770) );
  NOR2_X1 U519 ( .A1(n558), .A2(n770), .ZN(n432) );
  NOR2_X1 U520 ( .A1(n561), .A2(n432), .ZN(n433) );
  NOR2_X1 U521 ( .A1(n580), .A2(n433), .ZN(n435) );
  INV_X1 U522 ( .A(n436), .ZN(n438) );
  XNOR2_X1 U523 ( .A(n438), .B(n437), .ZN(n444) );
  NAND2_X1 U524 ( .A1(n496), .A2(G210), .ZN(n440) );
  XNOR2_X1 U525 ( .A(G146), .B(G137), .ZN(n439) );
  XNOR2_X1 U526 ( .A(n440), .B(n439), .ZN(n442) );
  XNOR2_X1 U527 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U528 ( .A(n444), .B(n443), .ZN(n447) );
  XNOR2_X1 U529 ( .A(n445), .B(G134), .ZN(n490) );
  INV_X1 U530 ( .A(n490), .ZN(n446) );
  XNOR2_X1 U531 ( .A(n446), .B(n504), .ZN(n476) );
  XNOR2_X1 U532 ( .A(n447), .B(n476), .ZN(n660) );
  OR2_X2 U533 ( .A1(n660), .A2(G902), .ZN(n449) );
  XNOR2_X1 U534 ( .A(KEYINPUT96), .B(G472), .ZN(n448) );
  XNOR2_X2 U535 ( .A(n449), .B(n448), .ZN(n518) );
  XNOR2_X2 U536 ( .A(n570), .B(KEYINPUT6), .ZN(n589) );
  XNOR2_X1 U537 ( .A(n450), .B(G140), .ZN(n451) );
  XNOR2_X1 U538 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n454) );
  NAND2_X1 U539 ( .A1(n760), .A2(G234), .ZN(n453) );
  XNOR2_X1 U540 ( .A(n454), .B(n453), .ZN(n488) );
  NAND2_X1 U541 ( .A1(n488), .A2(G221), .ZN(n455) );
  XNOR2_X1 U542 ( .A(n645), .B(n455), .ZN(n462) );
  XNOR2_X1 U543 ( .A(n475), .B(n456), .ZN(n460) );
  XNOR2_X1 U544 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U545 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U546 ( .A(n462), .B(n461), .ZN(n680) );
  INV_X1 U547 ( .A(n618), .ZN(n552) );
  NAND2_X1 U548 ( .A1(n552), .A2(G234), .ZN(n463) );
  XNOR2_X1 U549 ( .A(n463), .B(KEYINPUT20), .ZN(n467) );
  NAND2_X1 U550 ( .A1(n467), .A2(G217), .ZN(n464) );
  XNOR2_X1 U551 ( .A(n464), .B(KEYINPUT25), .ZN(n465) );
  XNOR2_X2 U552 ( .A(n466), .B(n465), .ZN(n723) );
  INV_X1 U553 ( .A(n467), .ZN(n469) );
  INV_X1 U554 ( .A(G221), .ZN(n468) );
  OR2_X1 U555 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U556 ( .A(n470), .B(KEYINPUT21), .ZN(n722) );
  NOR2_X2 U557 ( .A1(n723), .A2(n722), .ZN(n471) );
  XNOR2_X2 U558 ( .A(n471), .B(KEYINPUT68), .ZN(n533) );
  INV_X1 U559 ( .A(n533), .ZN(n719) );
  NAND2_X1 U560 ( .A1(n760), .A2(G227), .ZN(n472) );
  XNOR2_X1 U561 ( .A(n476), .B(n475), .ZN(n647) );
  XNOR2_X1 U562 ( .A(n477), .B(n647), .ZN(n683) );
  OR2_X2 U563 ( .A1(n683), .A2(G902), .ZN(n478) );
  XNOR2_X2 U564 ( .A(n478), .B(G469), .ZN(n567) );
  XNOR2_X2 U565 ( .A(n567), .B(n367), .ZN(n597) );
  XNOR2_X1 U566 ( .A(n480), .B(n368), .ZN(n707) );
  NOR2_X1 U567 ( .A1(n530), .A2(n707), .ZN(n481) );
  XNOR2_X1 U568 ( .A(n481), .B(KEYINPUT34), .ZN(n511) );
  XOR2_X1 U569 ( .A(KEYINPUT101), .B(G122), .Z(n483) );
  XNOR2_X1 U570 ( .A(n483), .B(n482), .ZN(n487) );
  XOR2_X1 U571 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n485) );
  XNOR2_X1 U572 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n484) );
  XNOR2_X1 U573 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U574 ( .A(n487), .B(n486), .Z(n492) );
  NAND2_X1 U575 ( .A1(n488), .A2(G217), .ZN(n489) );
  XNOR2_X1 U576 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U577 ( .A(n492), .B(n491), .ZN(n657) );
  NAND2_X1 U578 ( .A1(n657), .A2(n508), .ZN(n495) );
  XNOR2_X1 U579 ( .A(G478), .B(KEYINPUT102), .ZN(n493) );
  XNOR2_X1 U580 ( .A(n493), .B(KEYINPUT103), .ZN(n494) );
  XNOR2_X1 U581 ( .A(n495), .B(n494), .ZN(n537) );
  XOR2_X1 U582 ( .A(KEYINPUT97), .B(KEYINPUT12), .Z(n498) );
  NAND2_X1 U583 ( .A1(G214), .A2(n496), .ZN(n497) );
  XNOR2_X1 U584 ( .A(n498), .B(n497), .ZN(n502) );
  XOR2_X1 U585 ( .A(KEYINPUT11), .B(KEYINPUT98), .Z(n500) );
  XNOR2_X1 U586 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U587 ( .A(n502), .B(n501), .ZN(n507) );
  XNOR2_X1 U588 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U589 ( .A(n645), .B(n505), .ZN(n506) );
  XNOR2_X1 U590 ( .A(n507), .B(n506), .ZN(n630) );
  NAND2_X1 U591 ( .A1(n630), .A2(n508), .ZN(n510) );
  XNOR2_X1 U592 ( .A(KEYINPUT13), .B(G475), .ZN(n509) );
  XNOR2_X1 U593 ( .A(n510), .B(n509), .ZN(n536) );
  NOR2_X1 U594 ( .A1(n537), .A2(n536), .ZN(n601) );
  NAND2_X1 U595 ( .A1(n511), .A2(n601), .ZN(n513) );
  XOR2_X1 U596 ( .A(KEYINPUT77), .B(KEYINPUT35), .Z(n512) );
  XNOR2_X2 U597 ( .A(n513), .B(n512), .ZN(n676) );
  AND2_X1 U598 ( .A1(n537), .A2(n536), .ZN(n739) );
  INV_X1 U599 ( .A(n739), .ZN(n514) );
  NOR2_X1 U600 ( .A1(n514), .A2(n722), .ZN(n515) );
  NAND2_X1 U601 ( .A1(n357), .A2(n515), .ZN(n517) );
  INV_X1 U602 ( .A(n597), .ZN(n720) );
  INV_X1 U603 ( .A(n356), .ZN(n519) );
  NOR2_X1 U604 ( .A1(n726), .A2(n519), .ZN(n520) );
  NAND2_X1 U605 ( .A1(n720), .A2(n520), .ZN(n521) );
  NOR2_X1 U606 ( .A1(n540), .A2(n521), .ZN(n545) );
  NOR2_X2 U607 ( .A1(n676), .A2(n545), .ZN(n529) );
  NAND2_X1 U608 ( .A1(n597), .A2(n356), .ZN(n522) );
  XNOR2_X1 U609 ( .A(n522), .B(KEYINPUT105), .ZN(n525) );
  XOR2_X1 U610 ( .A(KEYINPUT79), .B(n523), .Z(n524) );
  NAND2_X1 U611 ( .A1(n525), .A2(n524), .ZN(n526) );
  NAND2_X1 U612 ( .A1(n533), .A2(n726), .ZN(n531) );
  OR2_X1 U613 ( .A1(n720), .A2(n531), .ZN(n730) );
  NAND2_X1 U614 ( .A1(n567), .A2(n533), .ZN(n534) );
  XNOR2_X1 U615 ( .A(n534), .B(KEYINPUT94), .ZN(n575) );
  NOR2_X1 U616 ( .A1(n575), .A2(n726), .ZN(n535) );
  AND2_X1 U617 ( .A1(n357), .A2(n535), .ZN(n692) );
  NOR2_X1 U618 ( .A1(n705), .A2(n692), .ZN(n539) );
  INV_X1 U619 ( .A(n536), .ZN(n538) );
  NOR2_X1 U620 ( .A1(n538), .A2(n537), .ZN(n704) );
  XNOR2_X1 U621 ( .A(n704), .B(KEYINPUT104), .ZN(n608) );
  AND2_X1 U622 ( .A1(n538), .A2(n537), .ZN(n701) );
  NOR2_X1 U623 ( .A1(n608), .A2(n701), .ZN(n741) );
  XOR2_X1 U624 ( .A(KEYINPUT83), .B(n741), .Z(n577) );
  NOR2_X1 U625 ( .A1(n589), .A2(n356), .ZN(n541) );
  NAND2_X1 U626 ( .A1(n720), .A2(n541), .ZN(n542) );
  NOR2_X1 U627 ( .A1(n676), .A2(KEYINPUT44), .ZN(n543) );
  XNOR2_X1 U628 ( .A(n543), .B(KEYINPUT67), .ZN(n548) );
  INV_X1 U629 ( .A(n642), .ZN(n546) );
  NAND2_X1 U630 ( .A1(n675), .A2(n546), .ZN(n547) );
  NOR2_X1 U631 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U632 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U633 ( .A(n551), .B(KEYINPUT45), .ZN(n627) );
  NOR2_X1 U634 ( .A1(n627), .A2(n552), .ZN(n553) );
  BUF_X1 U635 ( .A(n554), .Z(n555) );
  XNOR2_X1 U636 ( .A(n555), .B(KEYINPUT38), .ZN(n736) );
  INV_X1 U637 ( .A(n737), .ZN(n610) );
  NAND2_X1 U638 ( .A1(n736), .A2(n610), .ZN(n556) );
  XOR2_X1 U639 ( .A(KEYINPUT112), .B(n556), .Z(n743) );
  NAND2_X1 U640 ( .A1(n739), .A2(n743), .ZN(n557) );
  XNOR2_X1 U641 ( .A(KEYINPUT41), .B(n557), .ZN(n735) );
  NOR2_X1 U642 ( .A1(G900), .A2(n558), .ZN(n559) );
  NAND2_X1 U643 ( .A1(n396), .A2(n559), .ZN(n560) );
  XNOR2_X1 U644 ( .A(n560), .B(KEYINPUT107), .ZN(n562) );
  OR2_X1 U645 ( .A1(n562), .A2(n561), .ZN(n573) );
  INV_X1 U646 ( .A(n573), .ZN(n563) );
  NOR2_X1 U647 ( .A1(n563), .A2(n722), .ZN(n564) );
  AND2_X1 U648 ( .A1(n356), .A2(n564), .ZN(n588) );
  NAND2_X1 U649 ( .A1(n726), .A2(n588), .ZN(n566) );
  XNOR2_X1 U650 ( .A(KEYINPUT28), .B(KEYINPUT111), .ZN(n565) );
  XNOR2_X1 U651 ( .A(n566), .B(n565), .ZN(n568) );
  AND2_X1 U652 ( .A1(n568), .A2(n567), .ZN(n578) );
  NAND2_X1 U653 ( .A1(n735), .A2(n578), .ZN(n569) );
  XNOR2_X1 U654 ( .A(n569), .B(KEYINPUT42), .ZN(n777) );
  NOR2_X1 U655 ( .A1(n570), .A2(n737), .ZN(n572) );
  XNOR2_X1 U656 ( .A(KEYINPUT110), .B(KEYINPUT30), .ZN(n571) );
  XNOR2_X1 U657 ( .A(n572), .B(n571), .ZN(n574) );
  NAND2_X1 U658 ( .A1(n609), .A2(n701), .ZN(n576) );
  NOR2_X1 U659 ( .A1(n577), .A2(KEYINPUT47), .ZN(n581) );
  INV_X1 U660 ( .A(n578), .ZN(n579) );
  OR2_X1 U661 ( .A1(n580), .A2(n579), .ZN(n582) );
  NOR2_X1 U662 ( .A1(n581), .A2(n582), .ZN(n584) );
  INV_X1 U663 ( .A(n582), .ZN(n699) );
  NOR2_X1 U664 ( .A1(n699), .A2(KEYINPUT47), .ZN(n583) );
  NOR2_X1 U665 ( .A1(n584), .A2(n583), .ZN(n587) );
  NAND2_X1 U666 ( .A1(n741), .A2(KEYINPUT47), .ZN(n585) );
  XOR2_X1 U667 ( .A(n585), .B(KEYINPUT82), .Z(n586) );
  NOR2_X1 U668 ( .A1(n587), .A2(n586), .ZN(n599) );
  NAND2_X1 U669 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U670 ( .A(n590), .B(KEYINPUT108), .ZN(n592) );
  INV_X1 U671 ( .A(n701), .ZN(n591) );
  OR2_X1 U672 ( .A1(n592), .A2(n591), .ZN(n612) );
  BUF_X1 U673 ( .A(n593), .Z(n594) );
  INV_X1 U674 ( .A(n594), .ZN(n595) );
  NOR2_X1 U675 ( .A1(n612), .A2(n595), .ZN(n596) );
  XNOR2_X1 U676 ( .A(n596), .B(KEYINPUT36), .ZN(n598) );
  NAND2_X1 U677 ( .A1(n598), .A2(n597), .ZN(n638) );
  NAND2_X1 U678 ( .A1(n599), .A2(n638), .ZN(n605) );
  INV_X1 U679 ( .A(n600), .ZN(n604) );
  INV_X1 U680 ( .A(n555), .ZN(n602) );
  NAND2_X1 U681 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U682 ( .A1(n604), .A2(n603), .ZN(n639) );
  NOR2_X1 U683 ( .A1(n605), .A2(n639), .ZN(n606) );
  XNOR2_X1 U684 ( .A(n607), .B(KEYINPUT48), .ZN(n621) );
  NAND2_X1 U685 ( .A1(n609), .A2(n608), .ZN(n641) );
  NAND2_X1 U686 ( .A1(n720), .A2(n610), .ZN(n611) );
  NOR2_X1 U687 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U688 ( .A(KEYINPUT43), .B(n613), .Z(n614) );
  NAND2_X1 U689 ( .A1(n614), .A2(n555), .ZN(n615) );
  XOR2_X1 U690 ( .A(KEYINPUT109), .B(n615), .Z(n776) );
  NAND2_X1 U691 ( .A1(n641), .A2(n776), .ZN(n616) );
  NOR2_X2 U692 ( .A1(n621), .A2(n616), .ZN(n714) );
  XOR2_X1 U693 ( .A(KEYINPUT87), .B(n618), .Z(n619) );
  NAND2_X1 U694 ( .A1(n619), .A2(KEYINPUT2), .ZN(n620) );
  INV_X1 U695 ( .A(n621), .ZN(n626) );
  NAND2_X1 U696 ( .A1(n641), .A2(KEYINPUT2), .ZN(n622) );
  XOR2_X1 U697 ( .A(KEYINPUT81), .B(n622), .Z(n624) );
  INV_X1 U698 ( .A(n776), .ZN(n623) );
  NOR2_X1 U699 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U700 ( .A1(n626), .A2(n625), .ZN(n629) );
  BUF_X1 U701 ( .A(n627), .Z(n628) );
  NAND2_X1 U702 ( .A1(n678), .A2(G475), .ZN(n632) );
  XNOR2_X1 U703 ( .A(n632), .B(n631), .ZN(n634) );
  INV_X1 U704 ( .A(G952), .ZN(n633) );
  NAND2_X1 U705 ( .A1(n633), .A2(n396), .ZN(n670) );
  NAND2_X1 U706 ( .A1(n634), .A2(n670), .ZN(n636) );
  INV_X1 U707 ( .A(KEYINPUT60), .ZN(n635) );
  XNOR2_X1 U708 ( .A(n636), .B(n635), .ZN(G60) );
  XOR2_X1 U709 ( .A(G125), .B(KEYINPUT37), .Z(n637) );
  XNOR2_X1 U710 ( .A(n638), .B(n637), .ZN(G27) );
  XOR2_X1 U711 ( .A(G143), .B(n639), .Z(G45) );
  XNOR2_X1 U712 ( .A(n640), .B(n766), .ZN(G3) );
  XNOR2_X1 U713 ( .A(n641), .B(G134), .ZN(G36) );
  XOR2_X1 U714 ( .A(G110), .B(KEYINPUT115), .Z(n643) );
  XOR2_X1 U715 ( .A(n643), .B(n642), .Z(G12) );
  XNOR2_X1 U716 ( .A(n644), .B(G131), .ZN(G33) );
  XOR2_X1 U717 ( .A(KEYINPUT4), .B(n645), .Z(n646) );
  XNOR2_X1 U718 ( .A(n647), .B(n646), .ZN(n649) );
  XNOR2_X1 U719 ( .A(n714), .B(n649), .ZN(n648) );
  NAND2_X1 U720 ( .A1(n648), .A2(n760), .ZN(n655) );
  XNOR2_X1 U721 ( .A(n649), .B(KEYINPUT125), .ZN(n650) );
  XNOR2_X1 U722 ( .A(G227), .B(n650), .ZN(n651) );
  NAND2_X1 U723 ( .A1(G900), .A2(n651), .ZN(n652) );
  NAND2_X1 U724 ( .A1(n396), .A2(n652), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n653), .B(KEYINPUT126), .ZN(n654) );
  NAND2_X1 U726 ( .A1(n655), .A2(n654), .ZN(G72) );
  NAND2_X1 U727 ( .A1(n678), .A2(G478), .ZN(n656) );
  XOR2_X1 U728 ( .A(n657), .B(n656), .Z(n658) );
  INV_X1 U729 ( .A(n670), .ZN(n688) );
  NOR2_X1 U730 ( .A1(n658), .A2(n688), .ZN(G63) );
  NAND2_X1 U731 ( .A1(n678), .A2(G472), .ZN(n662) );
  XNOR2_X1 U732 ( .A(KEYINPUT91), .B(KEYINPUT62), .ZN(n659) );
  XNOR2_X1 U733 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U734 ( .A(n662), .B(n661), .ZN(n663) );
  NAND2_X1 U735 ( .A1(n663), .A2(n670), .ZN(n664) );
  XNOR2_X1 U736 ( .A(n664), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U737 ( .A1(n678), .A2(G210), .ZN(n669) );
  BUF_X1 U738 ( .A(n665), .Z(n666) );
  XNOR2_X1 U739 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n667) );
  XNOR2_X1 U740 ( .A(n666), .B(n667), .ZN(n668) );
  XNOR2_X1 U741 ( .A(n669), .B(n668), .ZN(n671) );
  NAND2_X1 U742 ( .A1(n671), .A2(n670), .ZN(n673) );
  XNOR2_X1 U743 ( .A(KEYINPUT121), .B(KEYINPUT56), .ZN(n672) );
  XNOR2_X1 U744 ( .A(n673), .B(n672), .ZN(G51) );
  XOR2_X1 U745 ( .A(G119), .B(KEYINPUT127), .Z(n674) );
  XNOR2_X1 U746 ( .A(n675), .B(n674), .ZN(G21) );
  XOR2_X1 U747 ( .A(n677), .B(G122), .Z(G24) );
  NAND2_X1 U748 ( .A1(n682), .A2(G217), .ZN(n679) );
  XNOR2_X1 U749 ( .A(n680), .B(n679), .ZN(n681) );
  NOR2_X1 U750 ( .A1(n681), .A2(n688), .ZN(G66) );
  NAND2_X1 U751 ( .A1(n682), .A2(G469), .ZN(n687) );
  XOR2_X1 U752 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n684) );
  XNOR2_X1 U753 ( .A(n684), .B(KEYINPUT58), .ZN(n685) );
  XNOR2_X1 U754 ( .A(n683), .B(n685), .ZN(n686) );
  XNOR2_X1 U755 ( .A(n687), .B(n686), .ZN(n689) );
  NOR2_X1 U756 ( .A1(n689), .A2(n688), .ZN(G54) );
  XOR2_X1 U757 ( .A(G104), .B(KEYINPUT113), .Z(n691) );
  NAND2_X1 U758 ( .A1(n692), .A2(n701), .ZN(n690) );
  XNOR2_X1 U759 ( .A(n691), .B(n690), .ZN(G6) );
  XNOR2_X1 U760 ( .A(G107), .B(KEYINPUT114), .ZN(n696) );
  XOR2_X1 U761 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n694) );
  NAND2_X1 U762 ( .A1(n692), .A2(n704), .ZN(n693) );
  XNOR2_X1 U763 ( .A(n694), .B(n693), .ZN(n695) );
  XNOR2_X1 U764 ( .A(n696), .B(n695), .ZN(G9) );
  XOR2_X1 U765 ( .A(G128), .B(KEYINPUT29), .Z(n698) );
  NAND2_X1 U766 ( .A1(n699), .A2(n704), .ZN(n697) );
  XNOR2_X1 U767 ( .A(n698), .B(n697), .ZN(G30) );
  NAND2_X1 U768 ( .A1(n699), .A2(n701), .ZN(n700) );
  XNOR2_X1 U769 ( .A(n700), .B(G146), .ZN(G48) );
  NAND2_X1 U770 ( .A1(n705), .A2(n701), .ZN(n702) );
  XNOR2_X1 U771 ( .A(n702), .B(KEYINPUT116), .ZN(n703) );
  XNOR2_X1 U772 ( .A(G113), .B(n703), .ZN(G15) );
  NAND2_X1 U773 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U774 ( .A(n706), .B(G116), .ZN(G18) );
  INV_X1 U775 ( .A(n735), .ZN(n708) );
  NOR2_X1 U776 ( .A1(n708), .A2(n746), .ZN(n709) );
  NOR2_X1 U777 ( .A1(n709), .A2(n396), .ZN(n758) );
  INV_X1 U778 ( .A(KEYINPUT2), .ZN(n715) );
  AND2_X1 U779 ( .A1(n628), .A2(n715), .ZN(n710) );
  NOR2_X1 U780 ( .A1(n710), .A2(KEYINPUT84), .ZN(n711) );
  NOR2_X1 U781 ( .A1(n712), .A2(n711), .ZN(n718) );
  NAND2_X1 U782 ( .A1(n628), .A2(KEYINPUT84), .ZN(n713) );
  NAND2_X1 U783 ( .A1(n714), .A2(n713), .ZN(n716) );
  NAND2_X1 U784 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U785 ( .A1(n718), .A2(n717), .ZN(n756) );
  NAND2_X1 U786 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U787 ( .A(n721), .B(KEYINPUT50), .ZN(n729) );
  XOR2_X1 U788 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n725) );
  NAND2_X1 U789 ( .A1(n356), .A2(n722), .ZN(n724) );
  XOR2_X1 U790 ( .A(n725), .B(n724), .Z(n727) );
  NOR2_X1 U791 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U792 ( .A1(n729), .A2(n728), .ZN(n731) );
  AND2_X1 U793 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U794 ( .A(n732), .B(KEYINPUT119), .Z(n733) );
  XNOR2_X1 U795 ( .A(KEYINPUT51), .B(n733), .ZN(n734) );
  NAND2_X1 U796 ( .A1(n735), .A2(n734), .ZN(n750) );
  INV_X1 U797 ( .A(n736), .ZN(n738) );
  NAND2_X1 U798 ( .A1(n738), .A2(n737), .ZN(n740) );
  NAND2_X1 U799 ( .A1(n740), .A2(n739), .ZN(n745) );
  INV_X1 U800 ( .A(n741), .ZN(n742) );
  NAND2_X1 U801 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U802 ( .A1(n745), .A2(n744), .ZN(n748) );
  INV_X1 U803 ( .A(n746), .ZN(n747) );
  NAND2_X1 U804 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U805 ( .A1(n750), .A2(n749), .ZN(n752) );
  XOR2_X1 U806 ( .A(KEYINPUT52), .B(KEYINPUT120), .Z(n751) );
  XNOR2_X1 U807 ( .A(n752), .B(n751), .ZN(n754) );
  NOR2_X1 U808 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U809 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U810 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U811 ( .A(KEYINPUT53), .B(n759), .Z(G75) );
  NAND2_X1 U812 ( .A1(n396), .A2(G224), .ZN(n761) );
  XNOR2_X1 U813 ( .A(KEYINPUT61), .B(n761), .ZN(n762) );
  NAND2_X1 U814 ( .A1(n762), .A2(G898), .ZN(n763) );
  NAND2_X1 U815 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U816 ( .A(n765), .B(KEYINPUT123), .ZN(n773) );
  XNOR2_X1 U817 ( .A(n767), .B(n766), .ZN(n768) );
  XNOR2_X1 U818 ( .A(n769), .B(n768), .ZN(n771) );
  AND2_X1 U819 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U820 ( .A(n773), .B(n772), .Z(n774) );
  XNOR2_X1 U821 ( .A(KEYINPUT124), .B(n774), .ZN(G69) );
  XOR2_X1 U822 ( .A(G140), .B(KEYINPUT117), .Z(n775) );
  XNOR2_X1 U823 ( .A(n776), .B(n775), .ZN(G42) );
  XNOR2_X1 U824 ( .A(G137), .B(n777), .ZN(G39) );
endmodule

