//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 0 0 0 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n530, new_n531, new_n532, new_n533, new_n534, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n546,
    new_n547, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  AND2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI211_X1 g037(.A(G137), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT65), .B1(new_n465), .B2(G101), .ZN(new_n466));
  AND4_X1   g041(.A1(KEYINPUT65), .A2(new_n460), .A3(G101), .A4(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n460), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(G160));
  OR2_X1    g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n460), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n460), .A2(G112), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G136), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n473), .A2(new_n474), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n460), .ZN(new_n481));
  OAI221_X1 g056(.A(new_n476), .B1(new_n477), .B2(new_n478), .C1(new_n479), .C2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n482), .B(new_n483), .ZN(G162));
  OAI211_X1 g059(.A(G138), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n460), .A2(G138), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n480), .A2(KEYINPUT67), .A3(new_n488), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n487), .A2(new_n489), .A3(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n485), .A2(new_n486), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n492), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n490), .A2(new_n497), .ZN(G164));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(KEYINPUT69), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(KEYINPUT5), .A3(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  OR3_X1    g082(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT68), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n499), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT68), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(new_n516), .A3(G50), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n501), .A2(new_n503), .B1(new_n513), .B2(new_n514), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n512), .A2(new_n517), .B1(G88), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n506), .B1(new_n505), .B2(new_n507), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n508), .A2(new_n519), .A3(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  NAND2_X1  g097(.A1(new_n518), .A2(G89), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n515), .A2(G51), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n523), .A2(new_n524), .A3(new_n526), .A4(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  AND2_X1   g104(.A1(G77), .A2(G543), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n530), .B1(new_n504), .B2(G64), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(new_n507), .ZN(new_n532));
  XOR2_X1   g107(.A(KEYINPUT71), .B(G90), .Z(new_n533));
  AOI22_X1  g108(.A1(new_n518), .A2(new_n533), .B1(new_n515), .B2(G52), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(G301));
  INV_X1    g110(.A(G301), .ZN(G171));
  AOI22_X1  g111(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n507), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n515), .A2(G43), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n504), .A2(new_n509), .ZN(new_n540));
  INV_X1    g115(.A(G81), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(G188));
  NAND3_X1  g123(.A1(new_n509), .A2(G53), .A3(G543), .ZN(new_n549));
  XOR2_X1   g124(.A(KEYINPUT72), .B(KEYINPUT9), .Z(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n518), .A2(G91), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n515), .A2(KEYINPUT72), .A3(KEYINPUT9), .A4(G53), .ZN(new_n553));
  AND3_X1   g128(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  AND2_X1   g129(.A1(new_n504), .A2(G65), .ZN(new_n555));
  AND2_X1   g130(.A1(G78), .A2(G543), .ZN(new_n556));
  OAI211_X1 g131(.A(KEYINPUT73), .B(G651), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT73), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n556), .B1(new_n504), .B2(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n559), .B2(new_n507), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n554), .A2(new_n557), .A3(new_n560), .ZN(G299));
  NAND3_X1  g136(.A1(new_n504), .A2(G87), .A3(new_n509), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT74), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n518), .A2(new_n564), .A3(G87), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n515), .A2(KEYINPUT75), .A3(G49), .ZN(new_n567));
  INV_X1    g142(.A(new_n514), .ZN(new_n568));
  NOR2_X1   g143(.A1(KEYINPUT6), .A2(G651), .ZN(new_n569));
  OAI211_X1 g144(.A(G49), .B(G543), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(G74), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n501), .A2(new_n573), .A3(new_n503), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n567), .A2(new_n572), .B1(G651), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n566), .A2(new_n575), .ZN(G288));
  NAND3_X1  g151(.A1(new_n515), .A2(KEYINPUT77), .A3(G48), .ZN(new_n577));
  OAI211_X1 g152(.A(G48), .B(G543), .C1(new_n568), .C2(new_n569), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n518), .A2(G86), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(new_n501), .B2(new_n503), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT76), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI211_X1 g165(.A(KEYINPUT76), .B(G651), .C1(new_n585), .C2(new_n587), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n583), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G305));
  AOI22_X1  g168(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(new_n507), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n515), .A2(G47), .ZN(new_n596));
  INV_X1    g171(.A(G85), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n540), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n515), .A2(G54), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n504), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(new_n507), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n605));
  INV_X1    g180(.A(G92), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n540), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n518), .A2(KEYINPUT10), .A3(G92), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n604), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n601), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n601), .B1(new_n609), .B2(G868), .ZN(G321));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(G299), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(new_n612), .B2(G168), .ZN(G297));
  OAI21_X1  g189(.A(new_n613), .B1(new_n612), .B2(G168), .ZN(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n609), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n609), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G868), .B2(new_n543), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g196(.A1(new_n480), .A2(new_n465), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT78), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n625), .A2(G2100), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(G2100), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n461), .A2(new_n462), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n628), .A2(G2105), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G135), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n475), .A2(G123), .ZN(new_n631));
  OR2_X1    g206(.A1(G99), .A2(G2105), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n632), .B(G2104), .C1(G111), .C2(new_n460), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(G2096), .Z(new_n635));
  NAND3_X1  g210(.A1(new_n626), .A2(new_n627), .A3(new_n635), .ZN(G156));
  XOR2_X1   g211(.A(G2451), .B(G2454), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT79), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2443), .B(G2446), .Z(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n647), .ZN(new_n651));
  NAND4_X1  g226(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n651), .A4(new_n645), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n648), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n650), .B1(new_n648), .B2(new_n652), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n640), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n657), .A2(new_n639), .A3(new_n653), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n656), .A2(new_n658), .A3(G14), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(G401));
  XNOR2_X1  g235(.A(G2072), .B(G2078), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT17), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2084), .B(G2090), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT80), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT81), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n663), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT82), .ZN(new_n670));
  INV_X1    g245(.A(new_n661), .ZN(new_n671));
  AND2_X1   g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n663), .A2(new_n668), .ZN(new_n673));
  OR3_X1    g248(.A1(new_n672), .A2(new_n673), .A3(new_n665), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n665), .A2(new_n661), .A3(new_n666), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT18), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n670), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2096), .B(G2100), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g256(.A1(new_n670), .A2(new_n674), .A3(new_n677), .A4(new_n679), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(G227));
  XOR2_X1   g258(.A(G1991), .B(G1996), .Z(new_n684));
  XNOR2_X1  g259(.A(G1956), .B(G2474), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1961), .B(G1966), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1971), .B(G1976), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT19), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT20), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n685), .B(new_n686), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(new_n691), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n691), .A2(new_n685), .A3(new_n686), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NOR3_X1   g275(.A1(new_n694), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n698), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n692), .B(KEYINPUT20), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n699), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n684), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1981), .B(G1986), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n700), .B1(new_n694), .B2(new_n698), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n702), .A2(new_n703), .A3(new_n699), .ZN(new_n708));
  INV_X1    g283(.A(new_n684), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AND3_X1   g285(.A1(new_n705), .A2(new_n706), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n706), .B1(new_n705), .B2(new_n710), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(G229));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G22), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G166), .B2(new_n714), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G1971), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n592), .A2(new_n714), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G6), .B2(new_n714), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT32), .B(G1981), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n717), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(G16), .A2(G23), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT87), .ZN(new_n725));
  AND3_X1   g300(.A1(new_n566), .A2(new_n575), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n725), .B1(new_n566), .B2(new_n575), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n724), .B1(new_n728), .B2(G16), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT33), .B(G1976), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n723), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(KEYINPUT34), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT89), .B(KEYINPUT36), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT34), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n723), .A2(new_n736), .A3(new_n731), .A4(new_n732), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n475), .A2(G119), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT83), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n741));
  INV_X1    g316(.A(G107), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(G2105), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT84), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n745), .A2(new_n746), .B1(G131), .B2(new_n629), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n740), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(KEYINPUT85), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT85), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n740), .A2(new_n747), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT86), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n749), .A2(KEYINPUT86), .A3(new_n751), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n754), .A2(G29), .A3(new_n755), .ZN(new_n756));
  OR2_X1    g331(.A1(G25), .A2(G29), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT35), .B(G1991), .Z(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  AND3_X1   g334(.A1(new_n756), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n759), .B1(new_n756), .B2(new_n757), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n714), .A2(G24), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n599), .B2(new_n714), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1986), .ZN(new_n764));
  NOR3_X1   g339(.A1(new_n760), .A2(new_n761), .A3(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT88), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n737), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n766), .B1(new_n737), .B2(new_n765), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n734), .B(new_n735), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(G29), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(G35), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G162), .B2(new_n771), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G2090), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n609), .A2(new_n714), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G4), .B2(new_n714), .ZN(new_n778));
  INV_X1    g353(.A(G1348), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT24), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G34), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n771), .B1(new_n781), .B2(G34), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT92), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n784), .B2(new_n783), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G160), .B2(G29), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G2084), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n771), .A2(G32), .ZN(new_n789));
  NAND3_X1  g364(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT26), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n475), .A2(G129), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n465), .A2(G105), .ZN(new_n794));
  INV_X1    g369(.A(G141), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n481), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n789), .B1(new_n797), .B2(new_n771), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT27), .B(G1996), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NOR3_X1   g375(.A1(new_n780), .A2(new_n788), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT25), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G139), .B2(new_n629), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n480), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(new_n460), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n804), .A2(new_n806), .A3(G29), .ZN(new_n807));
  NOR2_X1   g382(.A1(G29), .A2(G33), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT91), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(G2072), .Z(new_n811));
  NAND2_X1  g386(.A1(new_n714), .A2(G5), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G171), .B2(new_n714), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n714), .A2(G21), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G168), .B2(new_n714), .ZN(new_n815));
  OAI22_X1  g390(.A1(new_n813), .A2(G1961), .B1(G1966), .B2(new_n815), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n634), .A2(KEYINPUT94), .A3(new_n771), .ZN(new_n817));
  OAI21_X1  g392(.A(KEYINPUT94), .B1(new_n634), .B2(new_n771), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT31), .B(G11), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT95), .B(G28), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n820), .A2(KEYINPUT30), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(KEYINPUT30), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(new_n771), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n818), .B(new_n819), .C1(new_n821), .C2(new_n823), .ZN(new_n824));
  NOR4_X1   g399(.A1(new_n811), .A2(new_n816), .A3(new_n817), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n815), .A2(G1966), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT93), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n813), .A2(G1961), .ZN(new_n828));
  INV_X1    g403(.A(G2078), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n487), .A2(new_n489), .A3(KEYINPUT4), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n496), .A2(new_n495), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n830), .A2(new_n492), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(G29), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n771), .A2(G27), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n828), .B1(new_n829), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(new_n829), .B2(new_n836), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n801), .A2(new_n825), .A3(new_n827), .A4(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n771), .A2(G26), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT28), .Z(new_n841));
  OAI21_X1  g416(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n842));
  INV_X1    g417(.A(G116), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n842), .B1(new_n843), .B2(G2105), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(G128), .B2(new_n475), .ZN(new_n845));
  AOI21_X1  g420(.A(KEYINPUT90), .B1(new_n629), .B2(G140), .ZN(new_n846));
  AND4_X1   g421(.A1(KEYINPUT90), .A2(new_n480), .A3(G140), .A4(new_n460), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n841), .B1(new_n848), .B2(G29), .ZN(new_n849));
  INV_X1    g424(.A(G2067), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(new_n779), .B2(new_n778), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n714), .A2(G20), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT23), .Z(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(G299), .B2(G16), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(G1956), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n714), .A2(G19), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n543), .B2(new_n714), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(G1341), .Z(new_n859));
  NAND3_X1  g434(.A1(new_n852), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  NOR3_X1   g435(.A1(new_n776), .A2(new_n839), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n770), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT36), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT89), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n737), .A2(new_n765), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT88), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(new_n767), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n864), .B1(new_n867), .B2(new_n734), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n862), .A2(new_n868), .ZN(G311));
  AOI22_X1  g444(.A1(new_n866), .A2(new_n767), .B1(KEYINPUT34), .B2(new_n733), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n770), .B(new_n861), .C1(new_n870), .C2(new_n864), .ZN(G150));
  NAND2_X1  g446(.A1(new_n609), .A2(G559), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT38), .ZN(new_n873));
  XNOR2_X1  g448(.A(KEYINPUT98), .B(G55), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n515), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(G93), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n875), .B1(new_n540), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(KEYINPUT99), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT99), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n875), .B(new_n879), .C1(new_n540), .C2(new_n876), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(G67), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n882), .B1(new_n501), .B2(new_n503), .ZN(new_n883));
  AND2_X1   g458(.A1(G80), .A2(G543), .ZN(new_n884));
  OAI21_X1  g459(.A(G651), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(KEYINPUT97), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT97), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n887), .B(G651), .C1(new_n883), .C2(new_n884), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n881), .A2(new_n543), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n543), .B1(new_n881), .B2(new_n889), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n873), .B(new_n892), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n893), .A2(KEYINPUT39), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(KEYINPUT39), .ZN(new_n895));
  XOR2_X1   g470(.A(KEYINPUT100), .B(G860), .Z(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n896), .B1(new_n881), .B2(new_n889), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT37), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(G145));
  XNOR2_X1  g475(.A(G164), .B(new_n848), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n624), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n629), .A2(G142), .ZN(new_n903));
  OR3_X1    g478(.A1(new_n460), .A2(KEYINPUT102), .A3(G118), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT102), .B1(new_n460), .B2(G118), .ZN(new_n905));
  OR2_X1    g480(.A1(G106), .A2(G2105), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n904), .A2(G2104), .A3(new_n905), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n475), .A2(G130), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n903), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n752), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT101), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n804), .A2(new_n806), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(new_n797), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n749), .A2(new_n751), .A3(new_n909), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n911), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n914), .B1(new_n911), .B2(new_n915), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n902), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(G162), .A2(new_n634), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(G162), .A2(new_n634), .ZN(new_n921));
  OAI22_X1  g496(.A1(new_n920), .A2(new_n921), .B1(new_n471), .B2(new_n468), .ZN(new_n922));
  INV_X1    g497(.A(new_n921), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n923), .A2(new_n919), .A3(G160), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n624), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n901), .B(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n914), .ZN(new_n928));
  INV_X1    g503(.A(new_n915), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n909), .B1(new_n749), .B2(new_n751), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n911), .A2(new_n914), .A3(new_n915), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n927), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n918), .A2(new_n925), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(G37), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n925), .B1(new_n918), .B2(new_n933), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n938), .B(KEYINPUT40), .Z(G395));
  XOR2_X1   g514(.A(new_n892), .B(new_n618), .Z(new_n940));
  OAI21_X1  g515(.A(KEYINPUT103), .B1(G299), .B2(new_n609), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n942));
  OAI21_X1  g517(.A(G651), .B1(new_n555), .B2(new_n556), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n942), .B1(new_n943), .B2(new_n558), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n607), .A2(new_n608), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n603), .A2(new_n507), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(new_n946), .A3(new_n602), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT103), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n944), .A2(new_n947), .A3(new_n948), .A4(new_n557), .ZN(new_n949));
  NAND2_X1  g524(.A1(G299), .A2(new_n609), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n941), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n940), .A2(new_n951), .ZN(new_n952));
  XOR2_X1   g527(.A(new_n952), .B(KEYINPUT104), .Z(new_n953));
  AND2_X1   g528(.A1(new_n949), .A2(new_n950), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n954), .A2(new_n955), .A3(KEYINPUT41), .A4(new_n941), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT41), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT105), .B1(new_n951), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n951), .A2(new_n957), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n956), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  OR2_X1    g536(.A1(new_n961), .A2(new_n940), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n592), .B(G303), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n728), .A2(G290), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n726), .A2(new_n727), .A3(new_n599), .ZN(new_n965));
  OR3_X1    g540(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT42), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n953), .A2(new_n962), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n969), .B1(new_n953), .B2(new_n962), .ZN(new_n971));
  OAI21_X1  g546(.A(G868), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n881), .A2(new_n889), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n612), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(G295));
  NAND2_X1  g550(.A1(new_n972), .A2(new_n974), .ZN(G331));
  XNOR2_X1  g551(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n891), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n524), .A2(new_n527), .A3(new_n526), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n532), .A2(new_n980), .A3(new_n523), .A4(new_n534), .ZN(new_n981));
  INV_X1    g556(.A(new_n534), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n531), .A2(new_n507), .ZN(new_n983));
  OAI21_X1  g558(.A(G286), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n881), .A2(new_n543), .A3(new_n889), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n979), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n985), .B1(new_n890), .B2(new_n891), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT107), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n988), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n892), .A2(KEYINPUT107), .A3(new_n986), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n960), .A2(new_n990), .B1(new_n994), .B2(new_n951), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n935), .B1(new_n995), .B2(new_n968), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n960), .A2(new_n990), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n994), .A2(new_n951), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n997), .A2(new_n968), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n978), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n995), .A2(new_n968), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n951), .B(KEYINPUT41), .ZN(new_n1002));
  INV_X1    g577(.A(new_n951), .ZN(new_n1003));
  OAI22_X1  g578(.A1(new_n1002), .A2(new_n994), .B1(new_n1003), .B2(new_n990), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1004), .A2(new_n966), .A3(new_n967), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1001), .A2(new_n1005), .A3(new_n935), .A4(new_n977), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1000), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1007), .A2(KEYINPUT44), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n1009));
  OR3_X1    g584(.A1(new_n996), .A2(new_n999), .A3(new_n978), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1001), .A2(new_n1005), .A3(new_n935), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT43), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1009), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1008), .A2(new_n1013), .ZN(G397));
  XOR2_X1   g589(.A(KEYINPUT108), .B(G1384), .Z(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT45), .B1(new_n833), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G40), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n468), .A2(new_n471), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n848), .B(new_n850), .ZN(new_n1020));
  INV_X1    g595(.A(new_n797), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(G1996), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1019), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  OR3_X1    g598(.A1(new_n1019), .A2(KEYINPUT109), .A3(G1996), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT109), .B1(new_n1019), .B2(G1996), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1023), .B1(new_n1026), .B2(new_n797), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1019), .B1(new_n752), .B2(new_n758), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(new_n752), .B2(new_n758), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1019), .ZN(new_n1032));
  INV_X1    g607(.A(G1986), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n599), .B(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1031), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n577), .A2(new_n580), .B1(G86), .B2(new_n518), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n588), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n1037), .A2(G1981), .ZN(new_n1038));
  XOR2_X1   g613(.A(KEYINPUT115), .B(G1981), .Z(new_n1039));
  AND3_X1   g614(.A1(new_n502), .A2(KEYINPUT5), .A3(G543), .ZN(new_n1040));
  AOI21_X1  g615(.A(G543), .B1(new_n502), .B2(KEYINPUT5), .ZN(new_n1041));
  OAI21_X1  g616(.A(G61), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n586), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT76), .B1(new_n1043), .B2(G651), .ZN(new_n1044));
  INV_X1    g619(.A(new_n591), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1036), .B(new_n1039), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n590), .A2(new_n591), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1049), .A2(KEYINPUT116), .A3(new_n1036), .A4(new_n1039), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1038), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G1384), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n833), .A2(new_n1052), .A3(new_n1018), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(G8), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1054), .B1(new_n1053), .B2(G8), .ZN(new_n1057));
  OAI22_X1  g632(.A1(new_n1051), .A2(KEYINPUT49), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT49), .ZN(new_n1059));
  AOI211_X1 g634(.A(new_n1059), .B(new_n1038), .C1(new_n1048), .C2(new_n1050), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n727), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n566), .A2(new_n575), .A3(new_n725), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1062), .A2(G1976), .A3(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT114), .B(G1976), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT52), .B1(G288), .B2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1064), .B(new_n1066), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1053), .A2(G8), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT113), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1069), .A2(new_n1055), .B1(G1976), .B2(new_n728), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1067), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1061), .A2(new_n1072), .ZN(new_n1073));
  OAI211_X1 g648(.A(KEYINPUT45), .B(new_n1015), .C1(new_n490), .C2(new_n497), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT67), .B1(new_n480), .B2(new_n488), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n831), .B1(new_n491), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(G1384), .B1(new_n1076), .B2(new_n830), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1074), .B(new_n1018), .C1(new_n1077), .C2(KEYINPUT45), .ZN(new_n1078));
  INV_X1    g653(.A(G1971), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT110), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n833), .A2(new_n1052), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT50), .ZN(new_n1083));
  INV_X1    g658(.A(G2090), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT50), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n833), .A2(new_n1085), .A3(new_n1052), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1083), .A2(new_n1084), .A3(new_n1018), .A4(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT111), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT110), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1078), .A2(new_n1089), .A3(new_n1079), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1018), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n1082), .B2(KEYINPUT50), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT111), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1092), .A2(new_n1093), .A3(new_n1084), .A4(new_n1086), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1081), .A2(new_n1088), .A3(new_n1090), .A4(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT112), .ZN(new_n1096));
  NAND2_X1  g671(.A1(G303), .A2(G8), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT55), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1100));
  NAND4_X1  g675(.A1(G303), .A2(KEYINPUT112), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1095), .A2(G8), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(G8), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1104), .B1(new_n1080), .B2(new_n1087), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n1105), .A2(new_n1102), .ZN(new_n1106));
  INV_X1    g681(.A(G1966), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1018), .B1(new_n1077), .B2(KEYINPUT45), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT45), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1082), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1107), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  XOR2_X1   g686(.A(KEYINPUT120), .B(G2084), .Z(new_n1112));
  NAND3_X1  g687(.A1(new_n1092), .A2(new_n1086), .A3(new_n1112), .ZN(new_n1113));
  AOI211_X1 g688(.A(new_n1104), .B(G286), .C1(new_n1111), .C2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1073), .A2(new_n1103), .A3(new_n1106), .A4(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT121), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT63), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT117), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(new_n1061), .B2(new_n1072), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1038), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n1059), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1051), .A2(KEYINPUT49), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1069), .A2(new_n1055), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1064), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT52), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1127), .A2(KEYINPUT117), .A3(new_n1129), .A4(new_n1067), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1120), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1095), .A2(G8), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1102), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1114), .A2(KEYINPUT63), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1134), .A2(new_n1103), .A3(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1131), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1116), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1118), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n833), .A2(new_n1018), .A3(new_n1052), .A4(new_n850), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(KEYINPUT122), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1077), .A2(new_n1142), .A3(new_n850), .A4(new_n1018), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1018), .B1(new_n1077), .B2(new_n1085), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1086), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n779), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n609), .B(KEYINPUT124), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1145), .A2(new_n1148), .A3(new_n1149), .A4(KEYINPUT60), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT60), .ZN(new_n1151));
  AOI21_X1  g726(.A(G1348), .B1(new_n1092), .B2(new_n1086), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1151), .B1(new_n1152), .B2(new_n1144), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1152), .A2(new_n1144), .A3(new_n1151), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n947), .A2(KEYINPUT124), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1150), .B(new_n1153), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  XOR2_X1   g731(.A(KEYINPUT58), .B(G1341), .Z(new_n1157));
  NAND2_X1  g732(.A1(new_n1053), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1158), .B1(new_n1078), .B2(G1996), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(new_n543), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(KEYINPUT59), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT59), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1159), .A2(new_n1162), .A3(new_n543), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(G1956), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1165), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT57), .ZN(new_n1167));
  XNOR2_X1  g742(.A(G299), .B(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1091), .B1(new_n1082), .B2(new_n1109), .ZN(new_n1169));
  XNOR2_X1  g744(.A(KEYINPUT56), .B(G2072), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1169), .A2(new_n1074), .A3(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1166), .A2(new_n1168), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1168), .B1(new_n1166), .B2(new_n1171), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1172), .B1(new_n1173), .B2(KEYINPUT61), .ZN(new_n1174));
  OR2_X1    g749(.A1(new_n1172), .A2(KEYINPUT61), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1156), .A2(new_n1164), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1166), .A2(new_n1171), .ZN(new_n1177));
  OR2_X1    g752(.A1(new_n1177), .A2(KEYINPUT123), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1168), .B1(new_n1177), .B2(KEYINPUT123), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n947), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1180));
  AOI22_X1  g755(.A1(new_n1178), .A2(new_n1179), .B1(new_n1180), .B2(new_n1172), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1176), .A2(new_n1181), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1073), .A2(new_n1103), .A3(new_n1106), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT53), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1184), .B1(new_n1078), .B2(G2078), .ZN(new_n1185));
  INV_X1    g760(.A(G1961), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1186), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1169), .B1(new_n1109), .B2(new_n1082), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n829), .A2(KEYINPUT53), .ZN(new_n1189));
  OAI211_X1 g764(.A(new_n1185), .B(new_n1187), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g765(.A(G301), .B(KEYINPUT54), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1016), .A2(new_n1091), .A3(new_n1189), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1191), .B1(new_n1193), .B2(new_n1074), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1194), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1192), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1111), .A2(new_n1113), .A3(G168), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT51), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1104), .B1(KEYINPUT125), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(KEYINPUT51), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1197), .A2(new_n1199), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1203), .A2(G8), .A3(G286), .ZN(new_n1204));
  AND2_X1   g779(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1201), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1206));
  INV_X1    g781(.A(new_n1206), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1196), .B1(new_n1205), .B2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1182), .A2(new_n1183), .A3(new_n1208), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n1126), .B(KEYINPUT118), .ZN(new_n1210));
  NOR2_X1   g785(.A1(G288), .A2(G1976), .ZN(new_n1211));
  XOR2_X1   g786(.A(new_n1211), .B(KEYINPUT119), .Z(new_n1212));
  NAND2_X1  g787(.A1(new_n1127), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1210), .B1(new_n1213), .B2(new_n1121), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1120), .A2(new_n1130), .ZN(new_n1215));
  INV_X1    g790(.A(new_n1103), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1214), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1218));
  OAI21_X1  g793(.A(KEYINPUT62), .B1(new_n1218), .B2(new_n1206), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1219), .A2(KEYINPUT126), .ZN(new_n1220));
  INV_X1    g795(.A(KEYINPUT126), .ZN(new_n1221));
  OAI211_X1 g796(.A(new_n1221), .B(KEYINPUT62), .C1(new_n1218), .C2(new_n1206), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1223));
  AND2_X1   g798(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1224));
  INV_X1    g799(.A(KEYINPUT62), .ZN(new_n1225));
  NAND4_X1  g800(.A1(new_n1207), .A2(new_n1225), .A3(new_n1204), .A4(new_n1202), .ZN(new_n1226));
  AND2_X1   g801(.A1(new_n1190), .A2(G171), .ZN(new_n1227));
  NAND4_X1  g802(.A1(new_n1224), .A2(new_n1226), .A3(new_n1073), .A4(new_n1227), .ZN(new_n1228));
  OAI211_X1 g803(.A(new_n1209), .B(new_n1217), .C1(new_n1223), .C2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g804(.A(new_n1035), .B1(new_n1139), .B2(new_n1229), .ZN(new_n1230));
  AND4_X1   g805(.A1(new_n755), .A2(new_n1027), .A3(new_n754), .A4(new_n758), .ZN(new_n1231));
  NOR2_X1   g806(.A1(new_n848), .A2(G2067), .ZN(new_n1232));
  OAI21_X1  g807(.A(new_n1032), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  NOR3_X1   g808(.A1(new_n1019), .A2(G1986), .A3(G290), .ZN(new_n1234));
  XNOR2_X1  g809(.A(new_n1234), .B(KEYINPUT48), .ZN(new_n1235));
  XOR2_X1   g810(.A(new_n1026), .B(KEYINPUT46), .Z(new_n1236));
  INV_X1    g811(.A(KEYINPUT47), .ZN(new_n1237));
  INV_X1    g812(.A(new_n1020), .ZN(new_n1238));
  OAI21_X1  g813(.A(new_n1032), .B1(new_n1238), .B2(new_n1021), .ZN(new_n1239));
  NAND3_X1  g814(.A1(new_n1236), .A2(new_n1237), .A3(new_n1239), .ZN(new_n1240));
  INV_X1    g815(.A(new_n1240), .ZN(new_n1241));
  AOI21_X1  g816(.A(new_n1237), .B1(new_n1236), .B2(new_n1239), .ZN(new_n1242));
  OAI221_X1 g817(.A(new_n1233), .B1(new_n1031), .B2(new_n1235), .C1(new_n1241), .C2(new_n1242), .ZN(new_n1243));
  INV_X1    g818(.A(new_n1243), .ZN(new_n1244));
  NAND2_X1  g819(.A1(new_n1230), .A2(new_n1244), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g820(.A(KEYINPUT127), .ZN(new_n1247));
  AND3_X1   g821(.A1(new_n681), .A2(G319), .A3(new_n682), .ZN(new_n1248));
  NAND2_X1  g822(.A1(new_n659), .A2(new_n1248), .ZN(new_n1249));
  NOR2_X1   g823(.A1(G229), .A2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g824(.A(new_n1250), .B1(new_n936), .B2(new_n937), .ZN(new_n1251));
  INV_X1    g825(.A(new_n1251), .ZN(new_n1252));
  AOI21_X1  g826(.A(new_n1247), .B1(new_n1007), .B2(new_n1252), .ZN(new_n1253));
  AOI211_X1 g827(.A(KEYINPUT127), .B(new_n1251), .C1(new_n1000), .C2(new_n1006), .ZN(new_n1254));
  NOR2_X1   g828(.A1(new_n1253), .A2(new_n1254), .ZN(G308));
  NAND2_X1  g829(.A1(new_n1007), .A2(new_n1252), .ZN(G225));
endmodule


