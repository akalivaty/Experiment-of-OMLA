

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U552 ( .A1(n537), .A2(n762), .ZN(n766) );
  AND2_X1 U553 ( .A1(G2104), .A2(G2105), .ZN(n926) );
  NAND2_X1 U554 ( .A1(n596), .A2(n593), .ZN(n539) );
  INV_X1 U555 ( .A(G2105), .ZN(n621) );
  AND2_X1 U556 ( .A1(n575), .A2(n561), .ZN(n557) );
  AND2_X1 U557 ( .A1(n577), .A2(n578), .ZN(n574) );
  NOR2_X1 U558 ( .A1(n585), .A2(n589), .ZN(n538) );
  NOR2_X1 U559 ( .A1(n720), .A2(n719), .ZN(n734) );
  XNOR2_X1 U560 ( .A(n718), .B(KEYINPUT27), .ZN(n720) );
  AND2_X1 U561 ( .A1(n598), .A2(n597), .ZN(n596) );
  NAND2_X1 U562 ( .A1(n595), .A2(n594), .ZN(n593) );
  AND2_X1 U563 ( .A1(n544), .A2(n600), .ZN(n545) );
  AND2_X1 U564 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X2 U565 ( .A1(n554), .A2(n553), .ZN(n933) );
  NOR2_X1 U566 ( .A1(G2104), .A2(n621), .ZN(n620) );
  AND2_X2 U567 ( .A1(n621), .A2(G2104), .ZN(n930) );
  NOR2_X1 U568 ( .A1(G2104), .A2(KEYINPUT17), .ZN(n568) );
  BUF_X2 U569 ( .A(n629), .Z(n520) );
  XNOR2_X1 U570 ( .A(n620), .B(KEYINPUT68), .ZN(n629) );
  NAND2_X1 U571 ( .A1(n706), .A2(n705), .ZN(n729) );
  XNOR2_X1 U572 ( .A(n704), .B(KEYINPUT94), .ZN(n705) );
  OR2_X1 U573 ( .A1(G286), .A2(KEYINPUT96), .ZN(n572) );
  AND2_X1 U574 ( .A1(n593), .A2(n543), .ZN(n541) );
  AND2_X1 U575 ( .A1(G286), .A2(KEYINPUT96), .ZN(n573) );
  INV_X1 U576 ( .A(n573), .ZN(n551) );
  NAND2_X1 U577 ( .A1(n522), .A2(G8), .ZN(n549) );
  NAND2_X1 U578 ( .A1(n743), .A2(n742), .ZN(n751) );
  NOR2_X1 U579 ( .A1(n525), .A2(n684), .ZN(n685) );
  INV_X1 U580 ( .A(KEYINPUT64), .ZN(n604) );
  AND2_X1 U581 ( .A1(n761), .A2(n591), .ZN(n588) );
  INV_X1 U582 ( .A(n774), .ZN(n590) );
  XNOR2_X1 U583 ( .A(n759), .B(KEYINPUT98), .ZN(n592) );
  NOR2_X1 U584 ( .A1(n633), .A2(n603), .ZN(n602) );
  INV_X1 U585 ( .A(G40), .ZN(n603) );
  NAND2_X1 U586 ( .A1(G2104), .A2(KEYINPUT17), .ZN(n570) );
  NAND2_X1 U587 ( .A1(n765), .A2(n582), .ZN(n580) );
  NAND2_X1 U588 ( .A1(n583), .A2(n582), .ZN(n581) );
  NAND2_X1 U589 ( .A1(n565), .A2(n562), .ZN(n561) );
  NAND2_X1 U590 ( .A1(n822), .A2(n563), .ZN(n562) );
  NAND2_X1 U591 ( .A1(n567), .A2(n566), .ZN(n565) );
  NAND2_X1 U592 ( .A1(n564), .A2(n566), .ZN(n563) );
  NOR2_X1 U593 ( .A1(G651), .A2(n653), .ZN(n858) );
  NAND2_X1 U594 ( .A1(n933), .A2(G138), .ZN(n619) );
  XNOR2_X1 U595 ( .A(n571), .B(n625), .ZN(n628) );
  NAND2_X1 U596 ( .A1(n933), .A2(G137), .ZN(n571) );
  NOR2_X1 U597 ( .A1(n653), .A2(n610), .ZN(n863) );
  INV_X1 U598 ( .A(G168), .ZN(n680) );
  INV_X1 U599 ( .A(G1384), .ZN(n599) );
  NAND2_X1 U600 ( .A1(KEYINPUT66), .A2(G1384), .ZN(n600) );
  NOR2_X1 U601 ( .A1(n703), .A2(G2084), .ZN(n675) );
  NAND2_X1 U602 ( .A1(n751), .A2(n529), .ZN(n552) );
  NOR2_X1 U603 ( .A1(n789), .A2(n604), .ZN(n594) );
  INV_X1 U604 ( .A(KEYINPUT102), .ZN(n582) );
  NAND2_X1 U605 ( .A1(n1014), .A2(KEYINPUT100), .ZN(n586) );
  INV_X1 U606 ( .A(n605), .ZN(n564) );
  INV_X1 U607 ( .A(n822), .ZN(n567) );
  INV_X1 U608 ( .A(KEYINPUT40), .ZN(n566) );
  AND2_X1 U609 ( .A1(n569), .A2(n570), .ZN(n553) );
  NAND2_X1 U610 ( .A1(G2105), .A2(KEYINPUT17), .ZN(n569) );
  NAND2_X1 U611 ( .A1(n581), .A2(n579), .ZN(n578) );
  NAND2_X1 U612 ( .A1(n524), .A2(n580), .ZN(n579) );
  NAND2_X1 U613 ( .A1(n561), .A2(n534), .ZN(n555) );
  NOR2_X1 U614 ( .A1(n726), .A2(n725), .ZN(n1010) );
  NAND2_X1 U615 ( .A1(n526), .A2(n624), .ZN(n546) );
  NOR2_X1 U616 ( .A1(n628), .A2(n627), .ZN(n631) );
  XOR2_X1 U617 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  AND2_X1 U618 ( .A1(n748), .A2(n572), .ZN(n521) );
  NAND2_X1 U619 ( .A1(n521), .A2(KEYINPUT96), .ZN(n522) );
  AND2_X1 U620 ( .A1(n584), .A2(KEYINPUT102), .ZN(n523) );
  AND2_X1 U621 ( .A1(n777), .A2(n776), .ZN(n524) );
  AND2_X1 U622 ( .A1(n681), .A2(n680), .ZN(n525) );
  AND2_X1 U623 ( .A1(n619), .A2(n618), .ZN(n526) );
  AND2_X1 U624 ( .A1(n596), .A2(n593), .ZN(n703) );
  XOR2_X1 U625 ( .A(KEYINPUT28), .B(n735), .Z(n527) );
  AND2_X1 U626 ( .A1(n673), .A2(n599), .ZN(n528) );
  AND2_X1 U627 ( .A1(n521), .A2(n551), .ZN(n529) );
  AND2_X1 U628 ( .A1(n526), .A2(KEYINPUT66), .ZN(n530) );
  AND2_X1 U629 ( .A1(n573), .A2(G8), .ZN(n531) );
  AND2_X1 U630 ( .A1(n524), .A2(n582), .ZN(n532) );
  OR2_X1 U631 ( .A1(n764), .A2(n774), .ZN(n533) );
  NAND2_X1 U632 ( .A1(n545), .A2(n547), .ZN(n788) );
  NAND2_X1 U633 ( .A1(n605), .A2(KEYINPUT40), .ZN(n534) );
  INV_X1 U634 ( .A(n765), .ZN(n584) );
  NAND2_X1 U635 ( .A1(n533), .A2(n1005), .ZN(n765) );
  AND2_X1 U636 ( .A1(n822), .A2(n566), .ZN(n535) );
  AND2_X1 U637 ( .A1(n590), .A2(n586), .ZN(n536) );
  INV_X1 U638 ( .A(KEYINPUT100), .ZN(n591) );
  XNOR2_X1 U639 ( .A(n538), .B(KEYINPUT65), .ZN(n537) );
  NAND2_X1 U640 ( .A1(n539), .A2(KEYINPUT92), .ZN(n542) );
  NAND2_X1 U641 ( .A1(n542), .A2(n540), .ZN(n717) );
  NAND2_X1 U642 ( .A1(n541), .A2(n596), .ZN(n540) );
  INV_X1 U643 ( .A(KEYINPUT92), .ZN(n543) );
  NAND2_X1 U644 ( .A1(n546), .A2(n528), .ZN(n544) );
  INV_X1 U645 ( .A(n546), .ZN(G164) );
  NAND2_X1 U646 ( .A1(n530), .A2(n624), .ZN(n547) );
  NAND2_X1 U647 ( .A1(n552), .A2(n548), .ZN(n749) );
  NAND2_X1 U648 ( .A1(n550), .A2(n549), .ZN(n548) );
  NAND2_X1 U649 ( .A1(n751), .A2(n531), .ZN(n550) );
  NAND2_X1 U650 ( .A1(n568), .A2(n621), .ZN(n554) );
  NAND2_X1 U651 ( .A1(n556), .A2(n555), .ZN(n560) );
  NAND2_X1 U652 ( .A1(n557), .A2(n574), .ZN(n556) );
  NAND2_X1 U653 ( .A1(n558), .A2(n574), .ZN(n559) );
  AND2_X1 U654 ( .A1(n575), .A2(n535), .ZN(n558) );
  NAND2_X1 U655 ( .A1(n560), .A2(n559), .ZN(G329) );
  NOR2_X1 U656 ( .A1(n753), .A2(n678), .ZN(n679) );
  NAND2_X1 U657 ( .A1(n587), .A2(n536), .ZN(n585) );
  NAND2_X1 U658 ( .A1(n766), .A2(n532), .ZN(n577) );
  NAND2_X1 U659 ( .A1(n576), .A2(n523), .ZN(n575) );
  INV_X1 U660 ( .A(n766), .ZN(n576) );
  INV_X1 U661 ( .A(n524), .ZN(n583) );
  NAND2_X1 U662 ( .A1(n592), .A2(n588), .ZN(n587) );
  NOR2_X1 U663 ( .A1(n592), .A2(n591), .ZN(n589) );
  INV_X1 U664 ( .A(n788), .ZN(n595) );
  NAND2_X1 U665 ( .A1(n789), .A2(n604), .ZN(n597) );
  NAND2_X1 U666 ( .A1(n788), .A2(n604), .ZN(n598) );
  NAND2_X1 U667 ( .A1(n601), .A2(n602), .ZN(n789) );
  INV_X1 U668 ( .A(n634), .ZN(n601) );
  NOR2_X1 U669 ( .A1(n634), .A2(n633), .ZN(G160) );
  AND2_X1 U670 ( .A1(n816), .A2(n807), .ZN(n605) );
  INV_X1 U671 ( .A(KEYINPUT93), .ZN(n688) );
  XNOR2_X1 U672 ( .A(n689), .B(n688), .ZN(n690) );
  NOR2_X1 U673 ( .A1(n732), .A2(n731), .ZN(n733) );
  INV_X1 U674 ( .A(KEYINPUT29), .ZN(n737) );
  INV_X1 U675 ( .A(n1014), .ZN(n761) );
  INV_X1 U676 ( .A(KEYINPUT66), .ZN(n673) );
  INV_X1 U677 ( .A(KEYINPUT70), .ZN(n625) );
  NOR2_X1 U678 ( .A1(G543), .A2(G651), .ZN(n862) );
  NAND2_X1 U679 ( .A1(n862), .A2(G89), .ZN(n606) );
  XNOR2_X1 U680 ( .A(n606), .B(KEYINPUT4), .ZN(n608) );
  XOR2_X1 U681 ( .A(G543), .B(KEYINPUT0), .Z(n653) );
  INV_X1 U682 ( .A(G651), .ZN(n610) );
  NAND2_X1 U683 ( .A1(G76), .A2(n863), .ZN(n607) );
  NAND2_X1 U684 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U685 ( .A(n609), .B(KEYINPUT5), .ZN(n616) );
  NAND2_X1 U686 ( .A1(G51), .A2(n858), .ZN(n613) );
  NOR2_X1 U687 ( .A1(G543), .A2(n610), .ZN(n611) );
  XOR2_X2 U688 ( .A(KEYINPUT1), .B(n611), .Z(n859) );
  NAND2_X1 U689 ( .A1(G63), .A2(n859), .ZN(n612) );
  NAND2_X1 U690 ( .A1(n613), .A2(n612), .ZN(n614) );
  XOR2_X1 U691 ( .A(KEYINPUT6), .B(n614), .Z(n615) );
  NAND2_X1 U692 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U693 ( .A(n617), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U694 ( .A1(G102), .A2(n930), .ZN(n618) );
  NAND2_X1 U695 ( .A1(G126), .A2(n629), .ZN(n623) );
  NAND2_X1 U696 ( .A1(G114), .A2(n926), .ZN(n622) );
  NAND2_X1 U697 ( .A1(G101), .A2(n930), .ZN(n626) );
  XNOR2_X1 U698 ( .A(n626), .B(KEYINPUT23), .ZN(n627) );
  NAND2_X1 U699 ( .A1(G125), .A2(n520), .ZN(n630) );
  NAND2_X1 U700 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U701 ( .A1(G113), .A2(n926), .ZN(n632) );
  XNOR2_X1 U702 ( .A(KEYINPUT69), .B(n632), .ZN(n633) );
  NAND2_X1 U703 ( .A1(G52), .A2(n858), .ZN(n636) );
  NAND2_X1 U704 ( .A1(G64), .A2(n859), .ZN(n635) );
  NAND2_X1 U705 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U706 ( .A(KEYINPUT72), .B(n637), .ZN(n642) );
  NAND2_X1 U707 ( .A1(G90), .A2(n862), .ZN(n639) );
  NAND2_X1 U708 ( .A1(G77), .A2(n863), .ZN(n638) );
  NAND2_X1 U709 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U710 ( .A(KEYINPUT9), .B(n640), .Z(n641) );
  NOR2_X1 U711 ( .A1(n642), .A2(n641), .ZN(G171) );
  NAND2_X1 U712 ( .A1(G88), .A2(n862), .ZN(n644) );
  NAND2_X1 U713 ( .A1(G75), .A2(n863), .ZN(n643) );
  NAND2_X1 U714 ( .A1(n644), .A2(n643), .ZN(n649) );
  NAND2_X1 U715 ( .A1(n858), .A2(G50), .ZN(n645) );
  XNOR2_X1 U716 ( .A(n645), .B(KEYINPUT80), .ZN(n647) );
  NAND2_X1 U717 ( .A1(G62), .A2(n859), .ZN(n646) );
  NAND2_X1 U718 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U719 ( .A1(n649), .A2(n648), .ZN(G166) );
  XNOR2_X1 U720 ( .A(KEYINPUT87), .B(G166), .ZN(G303) );
  NAND2_X1 U721 ( .A1(G49), .A2(n858), .ZN(n651) );
  NAND2_X1 U722 ( .A1(G74), .A2(G651), .ZN(n650) );
  NAND2_X1 U723 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U724 ( .A1(n859), .A2(n652), .ZN(n656) );
  NAND2_X1 U725 ( .A1(G87), .A2(n653), .ZN(n654) );
  XOR2_X1 U726 ( .A(KEYINPUT77), .B(n654), .Z(n655) );
  NAND2_X1 U727 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U728 ( .A(KEYINPUT78), .B(n657), .ZN(G288) );
  NAND2_X1 U729 ( .A1(G73), .A2(n863), .ZN(n658) );
  XNOR2_X1 U730 ( .A(n658), .B(KEYINPUT2), .ZN(n665) );
  NAND2_X1 U731 ( .A1(G86), .A2(n862), .ZN(n660) );
  NAND2_X1 U732 ( .A1(G48), .A2(n858), .ZN(n659) );
  NAND2_X1 U733 ( .A1(n660), .A2(n659), .ZN(n663) );
  NAND2_X1 U734 ( .A1(G61), .A2(n859), .ZN(n661) );
  XNOR2_X1 U735 ( .A(KEYINPUT79), .B(n661), .ZN(n662) );
  NOR2_X1 U736 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U737 ( .A1(n665), .A2(n664), .ZN(G305) );
  NAND2_X1 U738 ( .A1(G47), .A2(n858), .ZN(n667) );
  NAND2_X1 U739 ( .A1(G60), .A2(n859), .ZN(n666) );
  NAND2_X1 U740 ( .A1(n667), .A2(n666), .ZN(n670) );
  NAND2_X1 U741 ( .A1(G85), .A2(n862), .ZN(n668) );
  XNOR2_X1 U742 ( .A(KEYINPUT71), .B(n668), .ZN(n669) );
  NOR2_X1 U743 ( .A1(n670), .A2(n669), .ZN(n672) );
  NAND2_X1 U744 ( .A1(n863), .A2(G72), .ZN(n671) );
  NAND2_X1 U745 ( .A1(n672), .A2(n671), .ZN(G290) );
  NAND2_X1 U746 ( .A1(n703), .A2(G8), .ZN(n774) );
  NOR2_X1 U747 ( .A1(G1966), .A2(n774), .ZN(n753) );
  INV_X1 U748 ( .A(KEYINPUT91), .ZN(n676) );
  XNOR2_X1 U749 ( .A(n676), .B(n675), .ZN(n750) );
  INV_X1 U750 ( .A(n750), .ZN(n677) );
  NAND2_X1 U751 ( .A1(G8), .A2(n677), .ZN(n678) );
  XNOR2_X1 U752 ( .A(n679), .B(KEYINPUT30), .ZN(n681) );
  INV_X1 U753 ( .A(G1961), .ZN(n954) );
  NAND2_X1 U754 ( .A1(n703), .A2(n954), .ZN(n683) );
  XNOR2_X1 U755 ( .A(KEYINPUT25), .B(G2078), .ZN(n1033) );
  NAND2_X1 U756 ( .A1(n717), .A2(n1033), .ZN(n682) );
  NAND2_X1 U757 ( .A1(n683), .A2(n682), .ZN(n739) );
  NOR2_X1 U758 ( .A1(G171), .A2(n739), .ZN(n684) );
  XOR2_X1 U759 ( .A(KEYINPUT31), .B(n685), .Z(n743) );
  NAND2_X1 U760 ( .A1(G1996), .A2(n539), .ZN(n687) );
  XOR2_X1 U761 ( .A(KEYINPUT67), .B(KEYINPUT26), .Z(n686) );
  XNOR2_X1 U762 ( .A(n687), .B(n686), .ZN(n691) );
  NAND2_X1 U763 ( .A1(G1341), .A2(n703), .ZN(n689) );
  NAND2_X1 U764 ( .A1(n691), .A2(n690), .ZN(n702) );
  NAND2_X1 U765 ( .A1(n862), .A2(G81), .ZN(n692) );
  XNOR2_X1 U766 ( .A(n692), .B(KEYINPUT12), .ZN(n694) );
  NAND2_X1 U767 ( .A1(G68), .A2(n863), .ZN(n693) );
  NAND2_X1 U768 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U769 ( .A(n695), .B(KEYINPUT13), .ZN(n697) );
  NAND2_X1 U770 ( .A1(G43), .A2(n858), .ZN(n696) );
  NAND2_X1 U771 ( .A1(n697), .A2(n696), .ZN(n700) );
  NAND2_X1 U772 ( .A1(n859), .A2(G56), .ZN(n698) );
  XOR2_X1 U773 ( .A(KEYINPUT14), .B(n698), .Z(n699) );
  NOR2_X1 U774 ( .A1(n700), .A2(n699), .ZN(n946) );
  INV_X1 U775 ( .A(n946), .ZN(n701) );
  NOR2_X1 U776 ( .A1(n702), .A2(n701), .ZN(n716) );
  NAND2_X1 U777 ( .A1(n717), .A2(G2067), .ZN(n706) );
  NAND2_X1 U778 ( .A1(n703), .A2(G1348), .ZN(n704) );
  NAND2_X1 U779 ( .A1(n858), .A2(G54), .ZN(n713) );
  NAND2_X1 U780 ( .A1(G92), .A2(n862), .ZN(n708) );
  NAND2_X1 U781 ( .A1(G79), .A2(n863), .ZN(n707) );
  NAND2_X1 U782 ( .A1(n708), .A2(n707), .ZN(n711) );
  NAND2_X1 U783 ( .A1(n859), .A2(G66), .ZN(n709) );
  XOR2_X1 U784 ( .A(KEYINPUT74), .B(n709), .Z(n710) );
  NOR2_X1 U785 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U786 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X2 U787 ( .A(KEYINPUT15), .B(n714), .ZN(n1025) );
  INV_X1 U788 ( .A(n1025), .ZN(n730) );
  NAND2_X1 U789 ( .A1(n729), .A2(n730), .ZN(n715) );
  NAND2_X1 U790 ( .A1(n716), .A2(n715), .ZN(n728) );
  NAND2_X1 U791 ( .A1(n717), .A2(G2072), .ZN(n718) );
  INV_X1 U792 ( .A(G1956), .ZN(n1068) );
  NOR2_X1 U793 ( .A1(n1068), .A2(n717), .ZN(n719) );
  NAND2_X1 U794 ( .A1(G53), .A2(n858), .ZN(n722) );
  NAND2_X1 U795 ( .A1(G65), .A2(n859), .ZN(n721) );
  NAND2_X1 U796 ( .A1(n722), .A2(n721), .ZN(n726) );
  NAND2_X1 U797 ( .A1(G91), .A2(n862), .ZN(n724) );
  NAND2_X1 U798 ( .A1(G78), .A2(n863), .ZN(n723) );
  NAND2_X1 U799 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U800 ( .A1(n734), .A2(n1010), .ZN(n727) );
  NAND2_X1 U801 ( .A1(n728), .A2(n727), .ZN(n732) );
  NOR2_X1 U802 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U803 ( .A(n733), .B(KEYINPUT95), .ZN(n736) );
  NOR2_X1 U804 ( .A1(n1010), .A2(n734), .ZN(n735) );
  NAND2_X1 U805 ( .A1(n736), .A2(n527), .ZN(n738) );
  XNOR2_X1 U806 ( .A(n738), .B(n737), .ZN(n741) );
  NAND2_X1 U807 ( .A1(G171), .A2(n739), .ZN(n740) );
  NAND2_X1 U808 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U809 ( .A1(n703), .A2(G2090), .ZN(n746) );
  NOR2_X1 U810 ( .A1(G1971), .A2(n774), .ZN(n744) );
  XOR2_X1 U811 ( .A(KEYINPUT97), .B(n744), .Z(n745) );
  NOR2_X1 U812 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U813 ( .A1(n747), .A2(G303), .ZN(n748) );
  XNOR2_X1 U814 ( .A(n749), .B(KEYINPUT32), .ZN(n757) );
  NAND2_X1 U815 ( .A1(G8), .A2(n750), .ZN(n755) );
  INV_X1 U816 ( .A(n751), .ZN(n752) );
  NOR2_X1 U817 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U818 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U819 ( .A1(n757), .A2(n756), .ZN(n769) );
  NOR2_X1 U820 ( .A1(G1976), .A2(G288), .ZN(n763) );
  NOR2_X1 U821 ( .A1(G1971), .A2(G303), .ZN(n758) );
  NOR2_X1 U822 ( .A1(n763), .A2(n758), .ZN(n1012) );
  NAND2_X1 U823 ( .A1(n769), .A2(n1012), .ZN(n759) );
  NAND2_X1 U824 ( .A1(G288), .A2(G1976), .ZN(n760) );
  XNOR2_X1 U825 ( .A(n760), .B(KEYINPUT99), .ZN(n1014) );
  INV_X1 U826 ( .A(KEYINPUT33), .ZN(n762) );
  NAND2_X1 U827 ( .A1(n763), .A2(KEYINPUT33), .ZN(n764) );
  XOR2_X1 U828 ( .A(G1981), .B(G305), .Z(n1005) );
  NOR2_X1 U829 ( .A1(G2090), .A2(G303), .ZN(n767) );
  XOR2_X1 U830 ( .A(KEYINPUT101), .B(n767), .Z(n768) );
  NAND2_X1 U831 ( .A1(G8), .A2(n768), .ZN(n770) );
  NAND2_X1 U832 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U833 ( .A1(n771), .A2(n774), .ZN(n777) );
  NOR2_X1 U834 ( .A1(G1981), .A2(G305), .ZN(n772) );
  XOR2_X1 U835 ( .A(n772), .B(KEYINPUT24), .Z(n773) );
  NOR2_X1 U836 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U837 ( .A(n775), .B(KEYINPUT90), .Z(n776) );
  NAND2_X1 U838 ( .A1(G104), .A2(n930), .ZN(n779) );
  NAND2_X1 U839 ( .A1(G140), .A2(n933), .ZN(n778) );
  NAND2_X1 U840 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U841 ( .A(KEYINPUT34), .B(n780), .ZN(n786) );
  NAND2_X1 U842 ( .A1(n926), .A2(G116), .ZN(n781) );
  XNOR2_X1 U843 ( .A(n781), .B(KEYINPUT88), .ZN(n783) );
  NAND2_X1 U844 ( .A1(G128), .A2(n520), .ZN(n782) );
  NAND2_X1 U845 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U846 ( .A(KEYINPUT35), .B(n784), .Z(n785) );
  NOR2_X1 U847 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U848 ( .A(KEYINPUT36), .B(n787), .ZN(n937) );
  XNOR2_X1 U849 ( .A(G2067), .B(KEYINPUT37), .ZN(n818) );
  NOR2_X1 U850 ( .A1(n937), .A2(n818), .ZN(n991) );
  NOR2_X1 U851 ( .A1(n595), .A2(n789), .ZN(n820) );
  NAND2_X1 U852 ( .A1(n991), .A2(n820), .ZN(n816) );
  XOR2_X1 U853 ( .A(G1986), .B(G290), .Z(n1018) );
  NAND2_X1 U854 ( .A1(G105), .A2(n930), .ZN(n790) );
  XNOR2_X1 U855 ( .A(n790), .B(KEYINPUT38), .ZN(n792) );
  NAND2_X1 U856 ( .A1(n926), .A2(G117), .ZN(n791) );
  NAND2_X1 U857 ( .A1(n792), .A2(n791), .ZN(n796) );
  NAND2_X1 U858 ( .A1(n933), .A2(G141), .ZN(n794) );
  NAND2_X1 U859 ( .A1(G129), .A2(n520), .ZN(n793) );
  NAND2_X1 U860 ( .A1(n794), .A2(n793), .ZN(n795) );
  OR2_X1 U861 ( .A1(n796), .A2(n795), .ZN(n912) );
  AND2_X1 U862 ( .A1(n912), .A2(G1996), .ZN(n805) );
  NAND2_X1 U863 ( .A1(G95), .A2(n930), .ZN(n798) );
  NAND2_X1 U864 ( .A1(G131), .A2(n933), .ZN(n797) );
  NAND2_X1 U865 ( .A1(n798), .A2(n797), .ZN(n803) );
  NAND2_X1 U866 ( .A1(G107), .A2(n926), .ZN(n800) );
  NAND2_X1 U867 ( .A1(G119), .A2(n520), .ZN(n799) );
  NAND2_X1 U868 ( .A1(n800), .A2(n799), .ZN(n801) );
  XOR2_X1 U869 ( .A(KEYINPUT89), .B(n801), .Z(n802) );
  OR2_X1 U870 ( .A1(n803), .A2(n802), .ZN(n913) );
  AND2_X1 U871 ( .A1(n913), .A2(G1991), .ZN(n804) );
  NOR2_X1 U872 ( .A1(n805), .A2(n804), .ZN(n979) );
  NAND2_X1 U873 ( .A1(n1018), .A2(n979), .ZN(n806) );
  NAND2_X1 U874 ( .A1(n806), .A2(n820), .ZN(n807) );
  XOR2_X1 U875 ( .A(KEYINPUT39), .B(KEYINPUT105), .Z(n815) );
  NOR2_X1 U876 ( .A1(G1996), .A2(n912), .ZN(n994) );
  NOR2_X1 U877 ( .A1(G1991), .A2(n913), .ZN(n988) );
  NOR2_X1 U878 ( .A1(G1986), .A2(G290), .ZN(n808) );
  XOR2_X1 U879 ( .A(n808), .B(KEYINPUT103), .Z(n809) );
  NOR2_X1 U880 ( .A1(n988), .A2(n809), .ZN(n811) );
  INV_X1 U881 ( .A(n979), .ZN(n810) );
  NOR2_X1 U882 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U883 ( .A(n812), .B(KEYINPUT104), .ZN(n813) );
  NOR2_X1 U884 ( .A1(n994), .A2(n813), .ZN(n814) );
  XNOR2_X1 U885 ( .A(n815), .B(n814), .ZN(n817) );
  NAND2_X1 U886 ( .A1(n817), .A2(n816), .ZN(n819) );
  NAND2_X1 U887 ( .A1(n937), .A2(n818), .ZN(n978) );
  NAND2_X1 U888 ( .A1(n819), .A2(n978), .ZN(n821) );
  NAND2_X1 U889 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U890 ( .A(G2451), .B(G2427), .ZN(n832) );
  XOR2_X1 U891 ( .A(G2430), .B(G2443), .Z(n824) );
  XNOR2_X1 U892 ( .A(G2435), .B(G2438), .ZN(n823) );
  XNOR2_X1 U893 ( .A(n824), .B(n823), .ZN(n828) );
  XOR2_X1 U894 ( .A(G2454), .B(KEYINPUT107), .Z(n826) );
  XNOR2_X1 U895 ( .A(G1341), .B(G1348), .ZN(n825) );
  XNOR2_X1 U896 ( .A(n826), .B(n825), .ZN(n827) );
  XOR2_X1 U897 ( .A(n828), .B(n827), .Z(n830) );
  XNOR2_X1 U898 ( .A(G2446), .B(KEYINPUT106), .ZN(n829) );
  XNOR2_X1 U899 ( .A(n830), .B(n829), .ZN(n831) );
  XNOR2_X1 U900 ( .A(n832), .B(n831), .ZN(n833) );
  AND2_X1 U901 ( .A1(n833), .A2(G14), .ZN(G401) );
  AND2_X1 U902 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U903 ( .A(G57), .ZN(G237) );
  NAND2_X1 U904 ( .A1(G7), .A2(G661), .ZN(n834) );
  XOR2_X1 U905 ( .A(n834), .B(KEYINPUT10), .Z(n977) );
  NAND2_X1 U906 ( .A1(n977), .A2(G567), .ZN(n835) );
  XOR2_X1 U907 ( .A(KEYINPUT11), .B(n835), .Z(G234) );
  NAND2_X1 U908 ( .A1(n946), .A2(G860), .ZN(G153) );
  INV_X1 U909 ( .A(G171), .ZN(G301) );
  NOR2_X1 U910 ( .A1(n1025), .A2(G868), .ZN(n836) );
  XNOR2_X1 U911 ( .A(n836), .B(KEYINPUT75), .ZN(n838) );
  NAND2_X1 U912 ( .A1(G868), .A2(G301), .ZN(n837) );
  NAND2_X1 U913 ( .A1(n838), .A2(n837), .ZN(G284) );
  XNOR2_X1 U914 ( .A(n1010), .B(KEYINPUT73), .ZN(G299) );
  NAND2_X1 U915 ( .A1(G286), .A2(G868), .ZN(n841) );
  INV_X1 U916 ( .A(G868), .ZN(n839) );
  NAND2_X1 U917 ( .A1(G299), .A2(n839), .ZN(n840) );
  NAND2_X1 U918 ( .A1(n841), .A2(n840), .ZN(G297) );
  INV_X1 U919 ( .A(G860), .ZN(n842) );
  NAND2_X1 U920 ( .A1(n842), .A2(G559), .ZN(n843) );
  NAND2_X1 U921 ( .A1(n843), .A2(n1025), .ZN(n844) );
  XNOR2_X1 U922 ( .A(n844), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U923 ( .A1(n1025), .A2(G868), .ZN(n845) );
  NOR2_X1 U924 ( .A1(G559), .A2(n845), .ZN(n847) );
  NOR2_X1 U925 ( .A1(G868), .A2(n701), .ZN(n846) );
  NOR2_X1 U926 ( .A1(n847), .A2(n846), .ZN(G282) );
  XOR2_X1 U927 ( .A(G2100), .B(KEYINPUT76), .Z(n856) );
  NAND2_X1 U928 ( .A1(G111), .A2(n926), .ZN(n849) );
  NAND2_X1 U929 ( .A1(G99), .A2(n930), .ZN(n848) );
  NAND2_X1 U930 ( .A1(n849), .A2(n848), .ZN(n852) );
  NAND2_X1 U931 ( .A1(n520), .A2(G123), .ZN(n850) );
  XOR2_X1 U932 ( .A(KEYINPUT18), .B(n850), .Z(n851) );
  NOR2_X1 U933 ( .A1(n852), .A2(n851), .ZN(n854) );
  NAND2_X1 U934 ( .A1(n933), .A2(G135), .ZN(n853) );
  NAND2_X1 U935 ( .A1(n854), .A2(n853), .ZN(n985) );
  XOR2_X1 U936 ( .A(G2096), .B(n985), .Z(n855) );
  NAND2_X1 U937 ( .A1(n856), .A2(n855), .ZN(G156) );
  NAND2_X1 U938 ( .A1(G559), .A2(n1025), .ZN(n857) );
  XOR2_X1 U939 ( .A(n857), .B(n946), .Z(n876) );
  NOR2_X1 U940 ( .A1(n876), .A2(G860), .ZN(n868) );
  NAND2_X1 U941 ( .A1(G55), .A2(n858), .ZN(n861) );
  NAND2_X1 U942 ( .A1(G67), .A2(n859), .ZN(n860) );
  NAND2_X1 U943 ( .A1(n861), .A2(n860), .ZN(n867) );
  NAND2_X1 U944 ( .A1(G93), .A2(n862), .ZN(n865) );
  NAND2_X1 U945 ( .A1(G80), .A2(n863), .ZN(n864) );
  NAND2_X1 U946 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U947 ( .A1(n867), .A2(n866), .ZN(n870) );
  XNOR2_X1 U948 ( .A(n868), .B(n870), .ZN(G145) );
  NOR2_X1 U949 ( .A1(G868), .A2(n870), .ZN(n869) );
  XNOR2_X1 U950 ( .A(n869), .B(KEYINPUT81), .ZN(n879) );
  XNOR2_X1 U951 ( .A(G166), .B(n870), .ZN(n873) );
  XNOR2_X1 U952 ( .A(G288), .B(G305), .ZN(n871) );
  XNOR2_X1 U953 ( .A(n871), .B(G299), .ZN(n872) );
  XNOR2_X1 U954 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U955 ( .A(KEYINPUT19), .B(n874), .ZN(n875) );
  XNOR2_X1 U956 ( .A(n875), .B(G290), .ZN(n949) );
  XOR2_X1 U957 ( .A(n876), .B(n949), .Z(n877) );
  NAND2_X1 U958 ( .A1(G868), .A2(n877), .ZN(n878) );
  NAND2_X1 U959 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U960 ( .A(KEYINPUT82), .B(n880), .ZN(G295) );
  NAND2_X1 U961 ( .A1(G2078), .A2(G2084), .ZN(n881) );
  XNOR2_X1 U962 ( .A(n881), .B(KEYINPUT20), .ZN(n882) );
  XNOR2_X1 U963 ( .A(n882), .B(KEYINPUT83), .ZN(n883) );
  NAND2_X1 U964 ( .A1(n883), .A2(G2090), .ZN(n886) );
  XOR2_X1 U965 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n884) );
  XNOR2_X1 U966 ( .A(KEYINPUT21), .B(n884), .ZN(n885) );
  XNOR2_X1 U967 ( .A(n886), .B(n885), .ZN(n887) );
  NAND2_X1 U968 ( .A1(n887), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U969 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U970 ( .A1(G132), .A2(G82), .ZN(n888) );
  XNOR2_X1 U971 ( .A(n888), .B(KEYINPUT86), .ZN(n889) );
  XNOR2_X1 U972 ( .A(n889), .B(KEYINPUT22), .ZN(n890) );
  NOR2_X1 U973 ( .A1(G218), .A2(n890), .ZN(n891) );
  NAND2_X1 U974 ( .A1(G96), .A2(n891), .ZN(n900) );
  NAND2_X1 U975 ( .A1(n900), .A2(G2106), .ZN(n895) );
  NAND2_X1 U976 ( .A1(G69), .A2(G120), .ZN(n892) );
  NOR2_X1 U977 ( .A1(G237), .A2(n892), .ZN(n893) );
  NAND2_X1 U978 ( .A1(G108), .A2(n893), .ZN(n901) );
  NAND2_X1 U979 ( .A1(n901), .A2(G567), .ZN(n894) );
  NAND2_X1 U980 ( .A1(n895), .A2(n894), .ZN(n902) );
  NAND2_X1 U981 ( .A1(G661), .A2(G483), .ZN(n896) );
  NOR2_X1 U982 ( .A1(n902), .A2(n896), .ZN(n899) );
  NAND2_X1 U983 ( .A1(n899), .A2(G36), .ZN(G176) );
  NAND2_X1 U984 ( .A1(G2106), .A2(n977), .ZN(G217) );
  AND2_X1 U985 ( .A1(G15), .A2(G2), .ZN(n897) );
  NAND2_X1 U986 ( .A1(G661), .A2(n897), .ZN(G259) );
  NAND2_X1 U987 ( .A1(G3), .A2(G1), .ZN(n898) );
  NAND2_X1 U988 ( .A1(n899), .A2(n898), .ZN(G188) );
  INV_X1 U990 ( .A(G132), .ZN(G219) );
  INV_X1 U991 ( .A(G120), .ZN(G236) );
  INV_X1 U992 ( .A(G82), .ZN(G220) );
  INV_X1 U993 ( .A(G69), .ZN(G235) );
  NOR2_X1 U994 ( .A1(n901), .A2(n900), .ZN(G325) );
  INV_X1 U995 ( .A(G325), .ZN(G261) );
  INV_X1 U996 ( .A(n902), .ZN(G319) );
  NAND2_X1 U997 ( .A1(G112), .A2(n926), .ZN(n904) );
  NAND2_X1 U998 ( .A1(G100), .A2(n930), .ZN(n903) );
  NAND2_X1 U999 ( .A1(n904), .A2(n903), .ZN(n910) );
  NAND2_X1 U1000 ( .A1(n520), .A2(G124), .ZN(n905) );
  XOR2_X1 U1001 ( .A(KEYINPUT44), .B(n905), .Z(n906) );
  XNOR2_X1 U1002 ( .A(n906), .B(KEYINPUT109), .ZN(n908) );
  NAND2_X1 U1003 ( .A1(G136), .A2(n933), .ZN(n907) );
  NAND2_X1 U1004 ( .A1(n908), .A2(n907), .ZN(n909) );
  NOR2_X1 U1005 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U1006 ( .A(KEYINPUT110), .B(n911), .ZN(G162) );
  XOR2_X1 U1007 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n915) );
  XNOR2_X1 U1008 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1009 ( .A(n915), .B(n914), .ZN(n944) );
  NAND2_X1 U1010 ( .A1(G130), .A2(n520), .ZN(n924) );
  NAND2_X1 U1011 ( .A1(n926), .A2(G118), .ZN(n916) );
  XNOR2_X1 U1012 ( .A(KEYINPUT111), .B(n916), .ZN(n922) );
  NAND2_X1 U1013 ( .A1(G106), .A2(n930), .ZN(n918) );
  NAND2_X1 U1014 ( .A1(G142), .A2(n933), .ZN(n917) );
  NAND2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1016 ( .A(KEYINPUT112), .B(n919), .Z(n920) );
  XNOR2_X1 U1017 ( .A(KEYINPUT45), .B(n920), .ZN(n921) );
  NOR2_X1 U1018 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1019 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1020 ( .A(n925), .B(n985), .ZN(n940) );
  NAND2_X1 U1021 ( .A1(G115), .A2(n926), .ZN(n928) );
  NAND2_X1 U1022 ( .A1(G127), .A2(n520), .ZN(n927) );
  NAND2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1024 ( .A(n929), .B(KEYINPUT47), .ZN(n932) );
  NAND2_X1 U1025 ( .A1(G103), .A2(n930), .ZN(n931) );
  NAND2_X1 U1026 ( .A1(n932), .A2(n931), .ZN(n936) );
  NAND2_X1 U1027 ( .A1(G139), .A2(n933), .ZN(n934) );
  XNOR2_X1 U1028 ( .A(KEYINPUT113), .B(n934), .ZN(n935) );
  NOR2_X1 U1029 ( .A1(n936), .A2(n935), .ZN(n981) );
  XNOR2_X1 U1030 ( .A(n981), .B(n937), .ZN(n938) );
  XNOR2_X1 U1031 ( .A(n938), .B(G162), .ZN(n939) );
  XNOR2_X1 U1032 ( .A(n940), .B(n939), .ZN(n942) );
  XNOR2_X1 U1033 ( .A(G164), .B(G160), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(n942), .B(n941), .ZN(n943) );
  XOR2_X1 U1035 ( .A(n944), .B(n943), .Z(n945) );
  NOR2_X1 U1036 ( .A1(G37), .A2(n945), .ZN(G395) );
  XOR2_X1 U1037 ( .A(n1025), .B(G286), .Z(n948) );
  XOR2_X1 U1038 ( .A(G301), .B(n946), .Z(n947) );
  XNOR2_X1 U1039 ( .A(n948), .B(n947), .ZN(n950) );
  XNOR2_X1 U1040 ( .A(n950), .B(n949), .ZN(n951) );
  NOR2_X1 U1041 ( .A1(G37), .A2(n951), .ZN(G397) );
  XNOR2_X1 U1042 ( .A(G1991), .B(KEYINPUT41), .ZN(n962) );
  XNOR2_X1 U1043 ( .A(n1068), .B(G1976), .ZN(n953) );
  XNOR2_X1 U1044 ( .A(G1986), .B(G1996), .ZN(n952) );
  XNOR2_X1 U1045 ( .A(n953), .B(n952), .ZN(n958) );
  XNOR2_X1 U1046 ( .A(n954), .B(G1966), .ZN(n956) );
  XNOR2_X1 U1047 ( .A(G1981), .B(G1971), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(n956), .B(n955), .ZN(n957) );
  XOR2_X1 U1049 ( .A(n958), .B(n957), .Z(n960) );
  XNOR2_X1 U1050 ( .A(KEYINPUT108), .B(G2474), .ZN(n959) );
  XNOR2_X1 U1051 ( .A(n960), .B(n959), .ZN(n961) );
  XNOR2_X1 U1052 ( .A(n962), .B(n961), .ZN(G229) );
  XOR2_X1 U1053 ( .A(G2096), .B(G2100), .Z(n964) );
  XNOR2_X1 U1054 ( .A(KEYINPUT42), .B(G2678), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(n964), .B(n963), .ZN(n968) );
  XOR2_X1 U1056 ( .A(KEYINPUT43), .B(G2090), .Z(n966) );
  XNOR2_X1 U1057 ( .A(G2067), .B(G2072), .ZN(n965) );
  XNOR2_X1 U1058 ( .A(n966), .B(n965), .ZN(n967) );
  XOR2_X1 U1059 ( .A(n968), .B(n967), .Z(n970) );
  XNOR2_X1 U1060 ( .A(G2078), .B(G2084), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(n970), .B(n969), .ZN(G227) );
  NOR2_X1 U1062 ( .A1(G395), .A2(G397), .ZN(n971) );
  XNOR2_X1 U1063 ( .A(n971), .B(KEYINPUT114), .ZN(n972) );
  NAND2_X1 U1064 ( .A1(G319), .A2(n972), .ZN(n973) );
  NOR2_X1 U1065 ( .A1(G401), .A2(n973), .ZN(n976) );
  NOR2_X1 U1066 ( .A1(G229), .A2(G227), .ZN(n974) );
  XOR2_X1 U1067 ( .A(KEYINPUT49), .B(n974), .Z(n975) );
  NAND2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(G225) );
  INV_X1 U1069 ( .A(G225), .ZN(G308) );
  INV_X1 U1070 ( .A(G96), .ZN(G221) );
  INV_X1 U1071 ( .A(G108), .ZN(G238) );
  INV_X1 U1072 ( .A(n977), .ZN(G223) );
  INV_X1 U1073 ( .A(KEYINPUT55), .ZN(n1049) );
  NAND2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n1001) );
  XNOR2_X1 U1075 ( .A(G164), .B(G2078), .ZN(n980) );
  XNOR2_X1 U1076 ( .A(n980), .B(KEYINPUT117), .ZN(n983) );
  XOR2_X1 U1077 ( .A(G2072), .B(n981), .Z(n982) );
  NOR2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1079 ( .A(KEYINPUT50), .B(n984), .ZN(n999) );
  XNOR2_X1 U1080 ( .A(G160), .B(G2084), .ZN(n986) );
  NAND2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1083 ( .A(n989), .B(KEYINPUT115), .ZN(n990) );
  NOR2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  XOR2_X1 U1085 ( .A(KEYINPUT116), .B(n992), .Z(n997) );
  XOR2_X1 U1086 ( .A(G2090), .B(G162), .Z(n993) );
  NOR2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1088 ( .A(KEYINPUT51), .B(n995), .ZN(n996) );
  NOR2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(KEYINPUT52), .B(n1002), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1049), .A2(n1003), .ZN(n1004) );
  NAND2_X1 U1094 ( .A1(n1004), .A2(G29), .ZN(n1056) );
  XNOR2_X1 U1095 ( .A(G1966), .B(G168), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(n1007), .B(KEYINPUT57), .ZN(n1024) );
  XOR2_X1 U1098 ( .A(n701), .B(G1341), .Z(n1009) );
  XOR2_X1 U1099 ( .A(G301), .B(G1961), .Z(n1008) );
  NAND2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1022) );
  XNOR2_X1 U1101 ( .A(n1010), .B(n1068), .ZN(n1017) );
  NAND2_X1 U1102 ( .A1(G1971), .A2(G303), .ZN(n1011) );
  NAND2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(KEYINPUT121), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1108 ( .A(KEYINPUT122), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1027) );
  XOR2_X1 U1111 ( .A(G1348), .B(n1025), .Z(n1026) );
  NOR2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1029) );
  XOR2_X1 U1113 ( .A(KEYINPUT56), .B(G16), .Z(n1028) );
  NOR2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1054) );
  XNOR2_X1 U1115 ( .A(G2067), .B(G26), .ZN(n1031) );
  XNOR2_X1 U1116 ( .A(G32), .B(G1996), .ZN(n1030) );
  NOR2_X1 U1117 ( .A1(n1031), .A2(n1030), .ZN(n1038) );
  XOR2_X1 U1118 ( .A(G2072), .B(G33), .Z(n1032) );
  NAND2_X1 U1119 ( .A1(n1032), .A2(G28), .ZN(n1036) );
  XNOR2_X1 U1120 ( .A(G27), .B(n1033), .ZN(n1034) );
  XNOR2_X1 U1121 ( .A(KEYINPUT119), .B(n1034), .ZN(n1035) );
  NOR2_X1 U1122 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NAND2_X1 U1123 ( .A1(n1038), .A2(n1037), .ZN(n1040) );
  XNOR2_X1 U1124 ( .A(G25), .B(G1991), .ZN(n1039) );
  NOR2_X1 U1125 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XOR2_X1 U1126 ( .A(KEYINPUT53), .B(n1041), .Z(n1044) );
  XOR2_X1 U1127 ( .A(G35), .B(KEYINPUT118), .Z(n1042) );
  XNOR2_X1 U1128 ( .A(G2090), .B(n1042), .ZN(n1043) );
  NAND2_X1 U1129 ( .A1(n1044), .A2(n1043), .ZN(n1047) );
  XNOR2_X1 U1130 ( .A(G34), .B(G2084), .ZN(n1045) );
  XNOR2_X1 U1131 ( .A(KEYINPUT54), .B(n1045), .ZN(n1046) );
  NOR2_X1 U1132 ( .A1(n1047), .A2(n1046), .ZN(n1048) );
  XNOR2_X1 U1133 ( .A(n1049), .B(n1048), .ZN(n1050) );
  NOR2_X1 U1134 ( .A1(G29), .A2(n1050), .ZN(n1051) );
  XOR2_X1 U1135 ( .A(KEYINPUT120), .B(n1051), .Z(n1052) );
  NAND2_X1 U1136 ( .A1(G11), .A2(n1052), .ZN(n1053) );
  NOR2_X1 U1137 ( .A1(n1054), .A2(n1053), .ZN(n1055) );
  NAND2_X1 U1138 ( .A1(n1056), .A2(n1055), .ZN(n1085) );
  XOR2_X1 U1139 ( .A(G16), .B(KEYINPUT123), .Z(n1083) );
  XNOR2_X1 U1140 ( .A(G1986), .B(G24), .ZN(n1061) );
  XNOR2_X1 U1141 ( .A(G1976), .B(G23), .ZN(n1058) );
  XNOR2_X1 U1142 ( .A(G1971), .B(G22), .ZN(n1057) );
  NOR2_X1 U1143 ( .A1(n1058), .A2(n1057), .ZN(n1059) );
  XNOR2_X1 U1144 ( .A(KEYINPUT127), .B(n1059), .ZN(n1060) );
  NOR2_X1 U1145 ( .A1(n1061), .A2(n1060), .ZN(n1062) );
  XNOR2_X1 U1146 ( .A(KEYINPUT58), .B(n1062), .ZN(n1080) );
  XOR2_X1 U1147 ( .A(G1966), .B(G21), .Z(n1074) );
  XNOR2_X1 U1148 ( .A(G1348), .B(KEYINPUT59), .ZN(n1063) );
  XNOR2_X1 U1149 ( .A(n1063), .B(G4), .ZN(n1067) );
  XNOR2_X1 U1150 ( .A(G1981), .B(G6), .ZN(n1065) );
  XNOR2_X1 U1151 ( .A(G1341), .B(G19), .ZN(n1064) );
  NOR2_X1 U1152 ( .A1(n1065), .A2(n1064), .ZN(n1066) );
  NAND2_X1 U1153 ( .A1(n1067), .A2(n1066), .ZN(n1071) );
  XNOR2_X1 U1154 ( .A(G20), .B(n1068), .ZN(n1069) );
  XNOR2_X1 U1155 ( .A(KEYINPUT125), .B(n1069), .ZN(n1070) );
  NOR2_X1 U1156 ( .A1(n1071), .A2(n1070), .ZN(n1072) );
  XNOR2_X1 U1157 ( .A(KEYINPUT60), .B(n1072), .ZN(n1073) );
  NAND2_X1 U1158 ( .A1(n1074), .A2(n1073), .ZN(n1077) );
  XNOR2_X1 U1159 ( .A(KEYINPUT124), .B(G1961), .ZN(n1075) );
  XNOR2_X1 U1160 ( .A(G5), .B(n1075), .ZN(n1076) );
  NOR2_X1 U1161 ( .A1(n1077), .A2(n1076), .ZN(n1078) );
  XNOR2_X1 U1162 ( .A(KEYINPUT126), .B(n1078), .ZN(n1079) );
  NAND2_X1 U1163 ( .A1(n1080), .A2(n1079), .ZN(n1081) );
  XNOR2_X1 U1164 ( .A(n1081), .B(KEYINPUT61), .ZN(n1082) );
  NOR2_X1 U1165 ( .A1(n1083), .A2(n1082), .ZN(n1084) );
  NOR2_X1 U1166 ( .A1(n1085), .A2(n1084), .ZN(n1086) );
  XOR2_X1 U1167 ( .A(n1086), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1168 ( .A(G150), .ZN(G311) );
endmodule

