//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n449, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n555, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n574, new_n575,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT65), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT66), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT67), .Z(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  INV_X1    g034(.A(new_n455), .ZN(new_n460));
  AOI22_X1  g035(.A1(new_n459), .A2(G2106), .B1(G567), .B2(new_n460), .ZN(G319));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n469), .A2(KEYINPUT68), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n462), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(KEYINPUT3), .B1(KEYINPUT69), .B2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(KEYINPUT69), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n468), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G101), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT70), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n479), .A2(KEYINPUT70), .A3(G101), .ZN(new_n483));
  AOI22_X1  g058(.A1(new_n478), .A2(G137), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n474), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G160));
  AND2_X1   g061(.A1(new_n478), .A2(G136), .ZN(new_n487));
  INV_X1    g062(.A(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(new_n488), .B2(G112), .ZN(new_n489));
  INV_X1    g064(.A(G100), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n489), .B1(new_n490), .B2(new_n488), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n476), .A2(new_n477), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT71), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n492), .A2(new_n495), .A3(G2105), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  AOI211_X1 g072(.A(new_n487), .B(new_n491), .C1(new_n497), .C2(G124), .ZN(G162));
  NAND2_X1  g073(.A1(new_n466), .A2(new_n471), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n488), .A2(G138), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g076(.A(KEYINPUT4), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  AND3_X1   g077(.A1(KEYINPUT69), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n503));
  OAI211_X1 g078(.A(KEYINPUT4), .B(G138), .C1(new_n503), .C2(new_n475), .ZN(new_n504));
  NAND2_X1  g079(.A1(G102), .A2(G2104), .ZN(new_n505));
  AOI21_X1  g080(.A(G2105), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g081(.A(G126), .B1(new_n503), .B2(new_n475), .ZN(new_n507));
  NAND2_X1  g082(.A1(G114), .A2(G2104), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n488), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR3_X1   g084(.A1(new_n502), .A2(new_n506), .A3(new_n509), .ZN(G164));
  XNOR2_X1  g085(.A(KEYINPUT5), .B(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n512));
  AND3_X1   g087(.A1(new_n512), .A2(KEYINPUT6), .A3(G651), .ZN(new_n513));
  AOI21_X1  g088(.A(KEYINPUT6), .B1(new_n512), .B2(G651), .ZN(new_n514));
  OAI211_X1 g089(.A(new_n511), .B(G88), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  OAI211_X1 g090(.A(G50), .B(G543), .C1(new_n513), .C2(new_n514), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT5), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G543), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n519), .A2(new_n521), .A3(G62), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n511), .A2(KEYINPUT73), .A3(G62), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n517), .B1(G651), .B2(new_n527), .ZN(G166));
  NOR2_X1   g103(.A1(new_n513), .A2(new_n514), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n519), .A2(new_n521), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G89), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n518), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G51), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n532), .A2(new_n534), .A3(new_n535), .A4(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G64), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n530), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n533), .A2(G52), .B1(new_n542), .B2(G651), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n531), .A2(G90), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(G171));
  OR2_X1    g120(.A1(new_n513), .A2(new_n514), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n546), .A2(G81), .A3(new_n511), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n546), .A2(G43), .A3(G543), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G56), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n530), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G651), .ZN(new_n552));
  AND3_X1   g127(.A1(new_n547), .A2(new_n548), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(G188));
  AND2_X1   g134(.A1(new_n511), .A2(G65), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  XOR2_X1   g136(.A(new_n561), .B(KEYINPUT75), .Z(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n531), .A2(G91), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n546), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n566));
  OAI211_X1 g141(.A(G53), .B(G543), .C1(new_n513), .C2(new_n514), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AND3_X1   g144(.A1(new_n566), .A2(KEYINPUT74), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g145(.A(KEYINPUT74), .B1(new_n566), .B2(new_n569), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n565), .B1(new_n570), .B2(new_n571), .ZN(G299));
  NAND2_X1  g147(.A1(new_n543), .A2(new_n544), .ZN(G301));
  NAND2_X1  g148(.A1(new_n527), .A2(G651), .ZN(new_n574));
  INV_X1    g149(.A(new_n517), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(G303));
  NAND2_X1  g151(.A1(new_n533), .A2(G49), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n531), .A2(G87), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G288));
  NAND3_X1  g155(.A1(new_n546), .A2(G48), .A3(G543), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n546), .A2(G86), .A3(new_n511), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT76), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n511), .A2(G61), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  AND2_X1   g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(G651), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n585), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n589), .B1(new_n586), .B2(new_n587), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(KEYINPUT76), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n584), .A2(new_n590), .A3(new_n592), .ZN(G305));
  AOI22_X1  g168(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(new_n589), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n531), .A2(G85), .ZN(new_n596));
  XNOR2_X1  g171(.A(KEYINPUT77), .B(G47), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n533), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(KEYINPUT78), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT78), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n595), .A2(new_n596), .A3(new_n598), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n600), .A2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n531), .A2(G92), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n530), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n533), .A2(G54), .B1(new_n609), .B2(G651), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n531), .A2(new_n611), .A3(G92), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n606), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT79), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n604), .B1(new_n615), .B2(G868), .ZN(G284));
  OAI21_X1  g191(.A(new_n604), .B1(new_n615), .B2(G868), .ZN(G321));
  NAND2_X1  g192(.A1(G286), .A2(G868), .ZN(new_n618));
  INV_X1    g193(.A(G299), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G868), .ZN(G280));
  XOR2_X1   g195(.A(G280), .B(KEYINPUT80), .Z(G297));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n615), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND3_X1  g198(.A1(new_n547), .A2(new_n548), .A3(new_n552), .ZN(new_n624));
  INV_X1    g199(.A(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g201(.A1(new_n615), .A2(new_n622), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(new_n625), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g204(.A1(new_n499), .A2(new_n479), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XOR2_X1   g206(.A(KEYINPUT81), .B(KEYINPUT13), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(KEYINPUT82), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n633), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n497), .A2(G123), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n478), .A2(G135), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT83), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n641), .B(new_n642), .C1(G111), .C2(new_n488), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n637), .A2(new_n638), .A3(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n644), .A2(G2096), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n634), .A2(KEYINPUT82), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(G2096), .ZN(new_n647));
  NAND4_X1  g222(.A1(new_n636), .A2(new_n645), .A3(new_n646), .A4(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT84), .B(KEYINPUT14), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2435), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT85), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2438), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2427), .B(G2430), .Z(new_n656));
  OAI21_X1  g231(.A(new_n651), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT86), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n655), .A2(new_n656), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n658), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1341), .B(G1348), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n661), .B1(new_n658), .B2(new_n662), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n664), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n658), .A2(new_n662), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(new_n660), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n665), .B1(new_n670), .B2(new_n663), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n650), .B1(new_n668), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n666), .B1(new_n664), .B2(new_n667), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n670), .A2(new_n665), .A3(new_n663), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n673), .A2(new_n649), .A3(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n672), .A2(G14), .A3(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G401));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G2067), .B(G2678), .Z(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G2072), .B(G2078), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n679), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT87), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n682), .B(KEYINPUT88), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT17), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n684), .B1(new_n686), .B2(new_n680), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n686), .A2(new_n680), .A3(new_n678), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n681), .A2(new_n678), .A3(new_n682), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT18), .Z(new_n690));
  NAND3_X1  g265(.A1(new_n687), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G2096), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G2100), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(G227));
  XOR2_X1   g269(.A(G1956), .B(G2474), .Z(new_n695));
  XOR2_X1   g270(.A(G1961), .B(G1966), .Z(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1971), .B(G1976), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT19), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n695), .A2(new_n696), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT20), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n701), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n698), .A2(new_n700), .A3(new_n702), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n705), .B(new_n706), .C1(new_n704), .C2(new_n703), .ZN(new_n707));
  XOR2_X1   g282(.A(G1991), .B(G1996), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT89), .B(G1986), .ZN(new_n712));
  INV_X1    g287(.A(G1981), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n711), .B(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(G229));
  NAND2_X1  g291(.A1(new_n615), .A2(G16), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G4), .B2(G16), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n718), .A2(KEYINPUT91), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(KEYINPUT91), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G1348), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(G27), .A2(G29), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G164), .B2(G29), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G2078), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT95), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n644), .A2(new_n728), .ZN(new_n729));
  OR2_X1    g304(.A1(G16), .A2(G21), .ZN(new_n730));
  INV_X1    g305(.A(G16), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(G286), .B2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G1966), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT94), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n734), .A2(new_n735), .ZN(new_n737));
  OAI221_X1 g312(.A(new_n726), .B1(new_n727), .B2(new_n729), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(G5), .A2(G16), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G171), .B2(G16), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n729), .A2(new_n727), .B1(new_n740), .B2(G1961), .ZN(new_n741));
  OR2_X1    g316(.A1(G29), .A2(G33), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n479), .A2(G103), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT25), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n478), .A2(G139), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n499), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n744), .B(new_n745), .C1(new_n746), .C2(new_n488), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n742), .B1(new_n747), .B2(new_n728), .ZN(new_n748));
  INV_X1    g323(.A(G2072), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n731), .A2(G19), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n553), .B2(new_n731), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G1341), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n732), .A2(new_n733), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n741), .A2(new_n750), .A3(new_n753), .A4(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n752), .A2(G1341), .ZN(new_n756));
  NOR3_X1   g331(.A1(new_n738), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  AND2_X1   g332(.A1(KEYINPUT24), .A2(G34), .ZN(new_n758));
  NOR2_X1   g333(.A1(KEYINPUT24), .A2(G34), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n728), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n485), .B2(new_n728), .ZN(new_n761));
  INV_X1    g336(.A(G2084), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OR2_X1    g338(.A1(G29), .A2(G32), .ZN(new_n764));
  NAND3_X1  g339(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT26), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n497), .B2(G129), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n479), .A2(G105), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n478), .A2(G141), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n764), .B1(new_n770), .B2(new_n728), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT27), .B(G1996), .ZN(new_n772));
  OAI221_X1 g347(.A(new_n763), .B1(G1961), .B2(new_n740), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT96), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n719), .A2(G1348), .A3(new_n720), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n723), .A2(new_n757), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT31), .B(G11), .ZN(new_n777));
  OAI221_X1 g352(.A(new_n777), .B1(new_n761), .B2(new_n762), .C1(G2078), .C2(new_n725), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n748), .A2(new_n749), .ZN(new_n779));
  OR2_X1    g354(.A1(KEYINPUT30), .A2(G28), .ZN(new_n780));
  NAND2_X1  g355(.A1(KEYINPUT30), .A2(G28), .ZN(new_n781));
  AOI21_X1  g356(.A(G29), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR4_X1   g357(.A1(new_n776), .A2(new_n778), .A3(new_n779), .A4(new_n782), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n731), .A2(KEYINPUT23), .A3(G20), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT23), .ZN(new_n785));
  INV_X1    g360(.A(G20), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(G16), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n784), .B(new_n787), .C1(new_n619), .C2(new_n731), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT97), .B(G1956), .Z(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n771), .A2(new_n772), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n728), .A2(G35), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G162), .B2(new_n728), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT29), .B(G2090), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n783), .A2(new_n790), .A3(new_n791), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n731), .A2(G6), .ZN(new_n797));
  AND4_X1   g372(.A1(new_n581), .A2(new_n590), .A3(new_n592), .A4(new_n582), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(new_n731), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT32), .B(G1981), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n731), .A2(G22), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G166), .B2(new_n731), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(G1971), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n803), .A2(G1971), .ZN(new_n805));
  NOR2_X1   g380(.A1(G16), .A2(G23), .ZN(new_n806));
  INV_X1    g381(.A(G288), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(G16), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT33), .B(G1976), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n801), .A2(new_n804), .A3(new_n805), .A4(new_n810), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n811), .A2(KEYINPUT34), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(KEYINPUT34), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n731), .A2(G24), .ZN(new_n814));
  INV_X1    g389(.A(G290), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n815), .B2(new_n731), .ZN(new_n816));
  INV_X1    g391(.A(G1986), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n497), .A2(G119), .B1(G131), .B2(new_n478), .ZN(new_n819));
  NOR2_X1   g394(.A1(G95), .A2(G2105), .ZN(new_n820));
  OAI21_X1  g395(.A(G2104), .B1(new_n488), .B2(G107), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  MUX2_X1   g397(.A(G25), .B(new_n822), .S(G29), .Z(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT35), .B(G1991), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n823), .B(new_n825), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n812), .A2(new_n813), .A3(new_n818), .A4(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT36), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT90), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n828), .A2(KEYINPUT90), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR3_X1   g407(.A1(new_n827), .A2(KEYINPUT90), .A3(new_n828), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT28), .ZN(new_n835));
  INV_X1    g410(.A(G26), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n836), .B2(G29), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n836), .A2(G29), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n478), .A2(G140), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT92), .ZN(new_n840));
  OR2_X1    g415(.A1(G104), .A2(G2105), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n841), .B(G2104), .C1(G116), .C2(new_n488), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT93), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(new_n497), .B2(G128), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n838), .B1(new_n845), .B2(G29), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n837), .B1(new_n846), .B2(new_n835), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(G2067), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n796), .A2(new_n834), .A3(new_n848), .ZN(G311));
  AND3_X1   g424(.A1(new_n783), .A2(new_n791), .A3(new_n795), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n832), .A2(new_n833), .ZN(new_n851));
  INV_X1    g426(.A(new_n848), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n850), .A2(new_n851), .A3(new_n852), .A4(new_n790), .ZN(G150));
  NAND2_X1  g428(.A1(G80), .A2(G543), .ZN(new_n854));
  INV_X1    g429(.A(G67), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n530), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G651), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT98), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n511), .B(G93), .C1(new_n513), .C2(new_n514), .ZN(new_n859));
  OAI211_X1 g434(.A(G55), .B(G543), .C1(new_n513), .C2(new_n514), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT98), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n856), .A2(new_n862), .A3(G651), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n858), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(G860), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT37), .Z(new_n866));
  AND2_X1   g441(.A1(new_n864), .A2(new_n553), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n864), .A2(new_n553), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XOR2_X1   g444(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n615), .A2(G559), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n866), .B1(new_n873), .B2(G860), .ZN(G145));
  XNOR2_X1  g449(.A(new_n822), .B(new_n770), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n631), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n845), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n840), .A2(new_n844), .A3(new_n631), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n747), .A2(G164), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n747), .A2(G164), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  AOI22_X1  g459(.A1(new_n878), .A2(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n497), .A2(G130), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT99), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n478), .A2(G142), .ZN(new_n888));
  NOR2_X1   g463(.A1(G106), .A2(G2105), .ZN(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(new_n488), .B2(G118), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NOR3_X1   g467(.A1(new_n884), .A2(new_n885), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n892), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n880), .A2(new_n883), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n878), .A2(new_n881), .A3(new_n882), .A4(new_n879), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n876), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n892), .B1(new_n884), .B2(new_n885), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n895), .A2(new_n894), .A3(new_n896), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n899), .A2(new_n875), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n644), .B(G160), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(G162), .ZN(new_n904));
  AOI21_X1  g479(.A(G37), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n904), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n898), .A2(new_n906), .A3(new_n901), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT100), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT100), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n898), .A2(new_n909), .A3(new_n901), .A4(new_n906), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n905), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g487(.A1(new_n864), .A2(new_n625), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n869), .B(KEYINPUT101), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(new_n627), .ZN(new_n915));
  INV_X1    g490(.A(new_n613), .ZN(new_n916));
  NAND2_X1  g491(.A1(G299), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n613), .B(new_n565), .C1(new_n571), .C2(new_n570), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(G299), .A2(new_n916), .A3(KEYINPUT102), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n915), .A2(KEYINPUT103), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n920), .A2(KEYINPUT41), .A3(new_n921), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT41), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n917), .A2(new_n918), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n915), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT103), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n915), .A2(new_n923), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n924), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT105), .ZN(new_n933));
  NAND2_X1  g508(.A1(G290), .A2(new_n807), .ZN(new_n934));
  NAND2_X1  g509(.A1(G303), .A2(KEYINPUT104), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n936));
  NAND2_X1  g511(.A1(G166), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n798), .ZN(new_n939));
  NAND3_X1  g514(.A1(G305), .A2(new_n935), .A3(new_n937), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n600), .A2(G288), .A3(new_n602), .ZN(new_n941));
  AND4_X1   g516(.A1(new_n934), .A2(new_n939), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  AOI22_X1  g517(.A1(new_n934), .A2(new_n941), .B1(new_n939), .B2(new_n940), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n933), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n934), .A2(new_n941), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n939), .A2(new_n940), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n934), .A2(new_n939), .A3(new_n940), .A4(new_n941), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n947), .A2(KEYINPUT105), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n944), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT42), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT42), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n952), .B1(new_n942), .B2(new_n943), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n932), .A2(new_n954), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n929), .A2(KEYINPUT103), .B1(new_n923), .B2(new_n915), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n953), .B(new_n951), .C1(new_n956), .C2(new_n924), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n913), .B1(new_n958), .B2(new_n625), .ZN(G295));
  OAI21_X1  g534(.A(new_n913), .B1(new_n958), .B2(new_n625), .ZN(G331));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n961));
  AOI21_X1  g536(.A(G286), .B1(G171), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(G301), .A2(KEYINPUT106), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n864), .A2(new_n553), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n624), .A2(new_n861), .A3(new_n858), .A4(new_n863), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n963), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI211_X1 g545(.A(KEYINPUT106), .B(G301), .C1(new_n867), .C2(new_n868), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n971), .A2(new_n962), .A3(new_n967), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n973), .B1(new_n927), .B2(new_n925), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n973), .A2(new_n922), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n950), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G37), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n922), .B1(new_n973), .B2(new_n926), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n917), .A2(new_n918), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n970), .A2(new_n972), .A3(KEYINPUT41), .A4(new_n979), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n978), .A2(new_n949), .A3(new_n944), .A4(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n976), .A2(new_n977), .A3(new_n981), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n982), .A2(KEYINPUT107), .A3(KEYINPUT43), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT107), .B1(new_n982), .B2(KEYINPUT43), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n928), .A2(new_n972), .A3(new_n970), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n973), .A2(new_n922), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n985), .A2(new_n949), .A3(new_n944), .A4(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT43), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n976), .A2(new_n987), .A3(new_n988), .A4(new_n977), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT44), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n983), .A2(new_n984), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n982), .A2(new_n988), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n976), .A2(new_n987), .A3(KEYINPUT43), .A4(new_n977), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT108), .B1(new_n991), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT108), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT107), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n982), .A2(KEYINPUT107), .A3(KEYINPUT43), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n998), .B(new_n995), .C1(new_n1003), .C2(new_n990), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n997), .A2(new_n1004), .ZN(G397));
  NAND2_X1  g580(.A1(new_n504), .A2(new_n505), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n488), .ZN(new_n1007));
  INV_X1    g582(.A(new_n509), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n500), .B1(new_n466), .B2(new_n471), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1007), .B(new_n1008), .C1(KEYINPUT4), .C2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G1384), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n474), .A2(G40), .A3(new_n484), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1996), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n770), .B(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G2067), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n845), .B(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1016), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g596(.A(new_n1021), .B(KEYINPUT109), .Z(new_n1022));
  NAND2_X1  g597(.A1(new_n815), .A2(new_n817), .ZN(new_n1023));
  NAND2_X1  g598(.A1(G290), .A2(G1986), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1016), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n822), .B(new_n825), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1026), .A2(new_n1016), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1022), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT50), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1010), .A2(new_n1031), .A3(new_n1011), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1030), .A2(new_n1032), .A3(new_n1014), .ZN(new_n1033));
  OR2_X1    g608(.A1(new_n1033), .A2(G1961), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1015), .B1(G164), .B2(G1384), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1010), .A2(KEYINPUT45), .A3(new_n1011), .ZN(new_n1036));
  INV_X1    g611(.A(G2078), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1014), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT120), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT120), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1038), .A2(new_n1042), .A3(new_n1039), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1034), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n1045));
  OR2_X1    g620(.A1(new_n1038), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1039), .B1(new_n1038), .B2(new_n1045), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(G171), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1050));
  XOR2_X1   g625(.A(new_n484), .B(KEYINPUT121), .Z(new_n1051));
  NOR2_X1   g626(.A1(new_n1051), .A2(new_n1039), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n474), .A2(G40), .A3(new_n1037), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1052), .A2(new_n1035), .A3(new_n1036), .A4(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1050), .A2(G301), .A3(new_n1034), .A4(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1049), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(G303), .A2(G8), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT110), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT111), .ZN(new_n1061));
  INV_X1    g636(.A(G8), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1062), .B1(new_n574), .B2(new_n575), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT111), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(new_n1064), .A3(KEYINPUT55), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1059), .A2(new_n1061), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1064), .B1(new_n1063), .B2(KEYINPUT55), .ZN(new_n1067));
  NOR4_X1   g642(.A1(G166), .A2(KEYINPUT111), .A3(new_n1058), .A4(new_n1062), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1063), .A2(KEYINPUT55), .ZN(new_n1069));
  OAI22_X1  g644(.A1(new_n1067), .A2(new_n1068), .B1(new_n1069), .B2(KEYINPUT110), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n1066), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G2090), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1035), .A2(new_n1014), .A3(new_n1036), .ZN(new_n1073));
  INV_X1    g648(.A(G1971), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1033), .A2(new_n1072), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1071), .B1(new_n1062), .B2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n577), .A2(new_n578), .A3(G1976), .A4(new_n579), .ZN(new_n1077));
  OAI211_X1 g652(.A(G8), .B(new_n1077), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1078));
  NAND2_X1  g653(.A1(KEYINPUT112), .A2(KEYINPUT52), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(G160), .A2(G40), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1079), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1081), .A2(G8), .A3(new_n1077), .A4(new_n1082), .ZN(new_n1083));
  OR3_X1    g658(.A1(new_n807), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1080), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n584), .A2(new_n713), .A3(new_n590), .A4(new_n592), .ZN(new_n1086));
  OAI21_X1  g661(.A(G1981), .B1(new_n583), .B2(new_n591), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT49), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1091), .A2(new_n1062), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1086), .A2(KEYINPUT49), .A3(new_n1087), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1090), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1085), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1030), .A2(new_n1032), .A3(new_n1014), .A4(new_n1072), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1062), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1066), .A2(new_n1070), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1076), .A2(new_n1095), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1076), .A2(new_n1095), .A3(KEYINPUT122), .A4(new_n1100), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n1029), .A2(new_n1056), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1030), .A2(new_n1032), .A3(new_n1014), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT116), .B(G1956), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n564), .A2(new_n563), .A3(new_n569), .A4(new_n566), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(KEYINPUT117), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n565), .B(KEYINPUT57), .C1(new_n570), .C2(new_n571), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT117), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1109), .A2(new_n1114), .A3(new_n1110), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1112), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  XOR2_X1   g691(.A(KEYINPUT56), .B(G2072), .Z(new_n1117));
  OAI211_X1 g692(.A(new_n1108), .B(new_n1116), .C1(new_n1073), .C2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1106), .A2(new_n722), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1091), .A2(new_n1019), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n613), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1108), .B1(new_n1073), .B2(new_n1117), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1116), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT58), .B(G1341), .ZN(new_n1126));
  OAI22_X1  g701(.A1(new_n1073), .A2(G1996), .B1(new_n1091), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n553), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT59), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1127), .A2(new_n1130), .A3(new_n553), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1125), .A2(KEYINPUT61), .A3(new_n1118), .ZN(new_n1133));
  OR2_X1    g708(.A1(new_n1118), .A2(KEYINPUT61), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n1119), .A2(new_n613), .A3(new_n1120), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT60), .B1(new_n1135), .B2(new_n1121), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1138), .A2(KEYINPUT60), .A3(new_n613), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1122), .B(new_n1125), .C1(new_n1137), .C2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1029), .B1(new_n1141), .B2(G301), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1034), .A2(new_n1041), .A3(new_n1043), .A4(new_n1054), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(G171), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(KEYINPUT123), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT123), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1143), .A2(new_n1146), .A3(G171), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1142), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1033), .A2(new_n762), .B1(new_n1073), .B2(new_n733), .ZN(new_n1149));
  NAND2_X1  g724(.A1(G286), .A2(G8), .ZN(new_n1150));
  OAI21_X1  g725(.A(KEYINPUT118), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1073), .A2(new_n733), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1030), .A2(new_n1032), .A3(new_n1014), .A4(new_n762), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT118), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1150), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1151), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT51), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1159), .B(G8), .C1(new_n1154), .C2(G286), .ZN(new_n1160));
  OAI211_X1 g735(.A(KEYINPUT51), .B(new_n1150), .C1(new_n1149), .C2(new_n1062), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1158), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1105), .A2(new_n1140), .A3(new_n1148), .A4(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1161), .A2(new_n1160), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1155), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1166));
  AOI211_X1 g741(.A(KEYINPUT118), .B(new_n1150), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1164), .B1(new_n1165), .B2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1158), .A2(KEYINPUT62), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1049), .ZN(new_n1173));
  AND4_X1   g748(.A1(KEYINPUT124), .A2(new_n1171), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1049), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1175));
  AOI21_X1  g750(.A(KEYINPUT124), .B1(new_n1175), .B2(new_n1172), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1163), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  AOI211_X1 g752(.A(new_n1062), .B(G286), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1076), .A2(new_n1095), .A3(new_n1100), .A4(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT63), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(KEYINPUT114), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT114), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1179), .A2(new_n1185), .A3(new_n1180), .ZN(new_n1186));
  INV_X1    g761(.A(G1976), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1094), .A2(new_n1187), .A3(new_n807), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(new_n1086), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT113), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1188), .A2(KEYINPUT113), .A3(new_n1086), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1191), .A2(new_n1092), .A3(new_n1192), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1095), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1186), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(KEYINPUT115), .B1(new_n1184), .B2(new_n1195), .ZN(new_n1196));
  AND2_X1   g771(.A1(new_n1186), .A2(new_n1194), .ZN(new_n1197));
  XNOR2_X1  g772(.A(new_n1071), .B(new_n1098), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1198), .A2(KEYINPUT63), .A3(new_n1095), .A4(new_n1178), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1199), .A2(KEYINPUT114), .A3(new_n1181), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT115), .ZN(new_n1201));
  NAND4_X1  g776(.A1(new_n1197), .A2(new_n1200), .A3(new_n1201), .A4(new_n1193), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1196), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1028), .B1(new_n1177), .B2(new_n1203), .ZN(new_n1204));
  OR3_X1    g779(.A1(new_n1022), .A2(new_n824), .A3(new_n822), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n840), .A2(new_n844), .A3(new_n1019), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1016), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n1016), .A2(G1996), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n1208), .B(KEYINPUT46), .ZN(new_n1209));
  INV_X1    g784(.A(new_n770), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1016), .B1(new_n1020), .B2(new_n1210), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  XNOR2_X1  g787(.A(new_n1212), .B(KEYINPUT125), .ZN(new_n1213));
  XNOR2_X1  g788(.A(new_n1213), .B(KEYINPUT47), .ZN(new_n1214));
  NOR2_X1   g789(.A1(new_n1023), .A2(new_n1016), .ZN(new_n1215));
  XNOR2_X1  g790(.A(new_n1215), .B(KEYINPUT48), .ZN(new_n1216));
  NOR3_X1   g791(.A1(new_n1022), .A2(new_n1027), .A3(new_n1216), .ZN(new_n1217));
  NOR3_X1   g792(.A1(new_n1207), .A2(new_n1214), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1204), .A2(new_n1218), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g794(.A1(new_n911), .A2(new_n676), .A3(new_n693), .ZN(new_n1221));
  NAND4_X1  g795(.A1(new_n992), .A2(G319), .A3(new_n715), .A4(new_n994), .ZN(new_n1222));
  INV_X1    g796(.A(KEYINPUT126), .ZN(new_n1223));
  OR3_X1    g797(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  OAI21_X1  g798(.A(new_n1223), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1225));
  NAND2_X1  g799(.A1(new_n1224), .A2(new_n1225), .ZN(G308));
  OR2_X1    g800(.A1(new_n1221), .A2(new_n1222), .ZN(G225));
endmodule


