

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581;

  XNOR2_X1 U322 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n377) );
  AND2_X1 U323 ( .A1(n451), .A2(n528), .ZN(n561) );
  XNOR2_X1 U324 ( .A(n365), .B(KEYINPUT65), .ZN(n366) );
  XOR2_X1 U325 ( .A(KEYINPUT90), .B(n479), .Z(n517) );
  XOR2_X1 U326 ( .A(n428), .B(n350), .Z(n290) );
  XOR2_X1 U327 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n291) );
  XOR2_X1 U328 ( .A(n386), .B(KEYINPUT91), .Z(n292) );
  XOR2_X1 U329 ( .A(KEYINPUT45), .B(n346), .Z(n293) );
  XNOR2_X1 U330 ( .A(KEYINPUT46), .B(KEYINPUT104), .ZN(n368) );
  XNOR2_X1 U331 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U332 ( .A(n316), .B(n315), .ZN(n325) );
  NOR2_X1 U333 ( .A1(n523), .A2(n544), .ZN(n527) );
  XNOR2_X1 U334 ( .A(n325), .B(n324), .ZN(n326) );
  NAND2_X1 U335 ( .A1(n481), .A2(n480), .ZN(n494) );
  NOR2_X1 U336 ( .A1(n416), .A2(n517), .ZN(n564) );
  XNOR2_X1 U337 ( .A(n367), .B(n366), .ZN(n457) );
  OR2_X1 U338 ( .A1(n496), .A2(n516), .ZN(n497) );
  XOR2_X1 U339 ( .A(n450), .B(n449), .Z(n528) );
  XOR2_X1 U340 ( .A(n391), .B(n390), .Z(n520) );
  XNOR2_X1 U341 ( .A(n452), .B(G190GAT), .ZN(n453) );
  XNOR2_X1 U342 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U343 ( .A(n454), .B(n453), .ZN(G1351GAT) );
  XOR2_X1 U344 ( .A(G113GAT), .B(G141GAT), .Z(n295) );
  XNOR2_X1 U345 ( .A(G169GAT), .B(G197GAT), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n295), .B(n294), .ZN(n310) );
  XNOR2_X1 U347 ( .A(G22GAT), .B(G15GAT), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n296), .B(G1GAT), .ZN(n339) );
  XOR2_X1 U349 ( .A(G29GAT), .B(n339), .Z(n298) );
  NAND2_X1 U350 ( .A1(G229GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U351 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U352 ( .A(n299), .B(G36GAT), .Z(n308) );
  XOR2_X1 U353 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n301) );
  XNOR2_X1 U354 ( .A(KEYINPUT29), .B(KEYINPUT30), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n301), .B(n300), .ZN(n306) );
  XOR2_X1 U356 ( .A(G43GAT), .B(G50GAT), .Z(n303) );
  XNOR2_X1 U357 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n302) );
  XNOR2_X1 U358 ( .A(n303), .B(n302), .ZN(n321) );
  XNOR2_X1 U359 ( .A(n321), .B(KEYINPUT67), .ZN(n304) );
  XNOR2_X1 U360 ( .A(n304), .B(G8GAT), .ZN(n305) );
  XNOR2_X1 U361 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U363 ( .A(n310), .B(n309), .Z(n565) );
  INV_X1 U364 ( .A(n565), .ZN(n560) );
  INV_X1 U365 ( .A(KEYINPUT106), .ZN(n362) );
  INV_X1 U366 ( .A(KEYINPUT36), .ZN(n329) );
  XOR2_X1 U367 ( .A(G92GAT), .B(KEYINPUT75), .Z(n312) );
  XNOR2_X1 U368 ( .A(G162GAT), .B(G106GAT), .ZN(n311) );
  XNOR2_X1 U369 ( .A(n312), .B(n311), .ZN(n327) );
  XOR2_X1 U370 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n314) );
  XOR2_X1 U371 ( .A(G29GAT), .B(G134GAT), .Z(n394) );
  XOR2_X1 U372 ( .A(G36GAT), .B(G190GAT), .Z(n383) );
  XNOR2_X1 U373 ( .A(n394), .B(n383), .ZN(n313) );
  XOR2_X1 U374 ( .A(n314), .B(n313), .Z(n316) );
  XNOR2_X1 U375 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n315) );
  XOR2_X1 U376 ( .A(KEYINPUT76), .B(KEYINPUT74), .Z(n318) );
  NAND2_X1 U377 ( .A1(G232GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U378 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U379 ( .A(n319), .B(KEYINPUT66), .Z(n323) );
  XNOR2_X1 U380 ( .A(G99GAT), .B(G85GAT), .ZN(n320) );
  XNOR2_X1 U381 ( .A(n320), .B(KEYINPUT72), .ZN(n357) );
  XNOR2_X1 U382 ( .A(n321), .B(n357), .ZN(n322) );
  XNOR2_X1 U383 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U384 ( .A(n327), .B(n326), .Z(n328) );
  XNOR2_X1 U385 ( .A(n329), .B(n328), .ZN(n579) );
  XOR2_X1 U386 ( .A(G64GAT), .B(G57GAT), .Z(n331) );
  XNOR2_X1 U387 ( .A(G127GAT), .B(G78GAT), .ZN(n330) );
  XNOR2_X1 U388 ( .A(n331), .B(n330), .ZN(n345) );
  XOR2_X1 U389 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n333) );
  XNOR2_X1 U390 ( .A(KEYINPUT15), .B(KEYINPUT77), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n333), .B(n332), .ZN(n338) );
  XNOR2_X1 U392 ( .A(G71GAT), .B(KEYINPUT70), .ZN(n334) );
  XNOR2_X1 U393 ( .A(n334), .B(KEYINPUT13), .ZN(n350) );
  XOR2_X1 U394 ( .A(n350), .B(KEYINPUT78), .Z(n336) );
  NAND2_X1 U395 ( .A1(G231GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U396 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U397 ( .A(n338), .B(n337), .ZN(n343) );
  XOR2_X1 U398 ( .A(G8GAT), .B(G183GAT), .Z(n387) );
  XOR2_X1 U399 ( .A(n387), .B(G155GAT), .Z(n341) );
  XNOR2_X1 U400 ( .A(n339), .B(G211GAT), .ZN(n340) );
  XNOR2_X1 U401 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U402 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n574) );
  NOR2_X1 U404 ( .A1(n579), .A2(n574), .ZN(n346) );
  XOR2_X1 U405 ( .A(G64GAT), .B(KEYINPUT73), .Z(n348) );
  XNOR2_X1 U406 ( .A(G204GAT), .B(G92GAT), .ZN(n347) );
  XNOR2_X1 U407 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U408 ( .A(G176GAT), .B(n349), .ZN(n390) );
  XOR2_X1 U409 ( .A(G106GAT), .B(G78GAT), .Z(n428) );
  NAND2_X1 U410 ( .A1(G230GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U411 ( .A(n290), .B(n351), .ZN(n355) );
  XOR2_X1 U412 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n353) );
  XNOR2_X1 U413 ( .A(KEYINPUT31), .B(KEYINPUT71), .ZN(n352) );
  XOR2_X1 U414 ( .A(n353), .B(n352), .Z(n354) );
  XNOR2_X1 U415 ( .A(n355), .B(n354), .ZN(n359) );
  XNOR2_X1 U416 ( .A(G120GAT), .B(G148GAT), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n356), .B(G57GAT), .ZN(n395) );
  XNOR2_X1 U418 ( .A(n395), .B(n357), .ZN(n358) );
  XOR2_X1 U419 ( .A(n359), .B(n358), .Z(n360) );
  XNOR2_X1 U420 ( .A(n390), .B(n360), .ZN(n367) );
  NOR2_X1 U421 ( .A1(n293), .A2(n367), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n362), .B(n361), .ZN(n363) );
  NOR2_X1 U423 ( .A1(n560), .A2(n363), .ZN(n364) );
  XOR2_X1 U424 ( .A(KEYINPUT107), .B(n364), .Z(n376) );
  INV_X1 U425 ( .A(KEYINPUT47), .ZN(n374) );
  INV_X1 U426 ( .A(KEYINPUT41), .ZN(n365) );
  NOR2_X1 U427 ( .A1(n457), .A2(n565), .ZN(n369) );
  INV_X1 U428 ( .A(n574), .ZN(n554) );
  NOR2_X1 U429 ( .A1(n370), .A2(n554), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n371), .B(KEYINPUT105), .ZN(n372) );
  NOR2_X1 U431 ( .A1(n372), .A2(n328), .ZN(n373) );
  XNOR2_X1 U432 ( .A(n374), .B(n373), .ZN(n375) );
  NOR2_X1 U433 ( .A1(n376), .A2(n375), .ZN(n378) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n545) );
  XOR2_X1 U435 ( .A(KEYINPUT81), .B(G218GAT), .Z(n380) );
  XNOR2_X1 U436 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n379) );
  XNOR2_X1 U437 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U438 ( .A(G197GAT), .B(n381), .Z(n418) );
  XNOR2_X1 U439 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n382) );
  XNOR2_X1 U440 ( .A(n291), .B(n382), .ZN(n448) );
  XOR2_X1 U441 ( .A(n383), .B(n448), .Z(n385) );
  NAND2_X1 U442 ( .A1(G226GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U443 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U444 ( .A(n387), .B(KEYINPUT92), .ZN(n388) );
  XNOR2_X1 U445 ( .A(n292), .B(n388), .ZN(n389) );
  XNOR2_X1 U446 ( .A(n418), .B(n389), .ZN(n391) );
  INV_X1 U447 ( .A(n520), .ZN(n466) );
  NOR2_X1 U448 ( .A1(n545), .A2(n466), .ZN(n393) );
  INV_X1 U449 ( .A(KEYINPUT54), .ZN(n392) );
  XNOR2_X1 U450 ( .A(n393), .B(n392), .ZN(n416) );
  XOR2_X1 U451 ( .A(n395), .B(n394), .Z(n397) );
  NAND2_X1 U452 ( .A1(G225GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U453 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U454 ( .A(n398), .B(KEYINPUT6), .Z(n402) );
  XOR2_X1 U455 ( .A(G127GAT), .B(KEYINPUT0), .Z(n400) );
  XNOR2_X1 U456 ( .A(G113GAT), .B(KEYINPUT79), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n447) );
  XNOR2_X1 U458 ( .A(G1GAT), .B(n447), .ZN(n401) );
  XNOR2_X1 U459 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U460 ( .A(KEYINPUT87), .B(KEYINPUT4), .Z(n404) );
  XNOR2_X1 U461 ( .A(G85GAT), .B(KEYINPUT86), .ZN(n403) );
  XNOR2_X1 U462 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U463 ( .A(n406), .B(n405), .Z(n415) );
  XNOR2_X1 U464 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n407), .B(KEYINPUT82), .ZN(n408) );
  XOR2_X1 U466 ( .A(n408), .B(KEYINPUT2), .Z(n410) );
  XNOR2_X1 U467 ( .A(G141GAT), .B(G162GAT), .ZN(n409) );
  XNOR2_X1 U468 ( .A(n410), .B(n409), .ZN(n417) );
  XOR2_X1 U469 ( .A(KEYINPUT88), .B(KEYINPUT1), .Z(n412) );
  XNOR2_X1 U470 ( .A(KEYINPUT5), .B(KEYINPUT89), .ZN(n411) );
  XNOR2_X1 U471 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n417), .B(n413), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n415), .B(n414), .ZN(n479) );
  XNOR2_X1 U474 ( .A(n418), .B(n417), .ZN(n432) );
  XOR2_X1 U475 ( .A(KEYINPUT22), .B(G204GAT), .Z(n420) );
  XNOR2_X1 U476 ( .A(G50GAT), .B(G22GAT), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U478 ( .A(KEYINPUT23), .B(KEYINPUT84), .Z(n422) );
  XNOR2_X1 U479 ( .A(KEYINPUT24), .B(G148GAT), .ZN(n421) );
  XNOR2_X1 U480 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U481 ( .A(n424), .B(n423), .Z(n430) );
  XOR2_X1 U482 ( .A(KEYINPUT85), .B(KEYINPUT83), .Z(n426) );
  NAND2_X1 U483 ( .A1(G228GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U484 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U485 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n472) );
  NAND2_X1 U488 ( .A1(n564), .A2(n472), .ZN(n435) );
  XOR2_X1 U489 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n433) );
  XNOR2_X1 U490 ( .A(KEYINPUT55), .B(n433), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n451) );
  XOR2_X1 U492 ( .A(G183GAT), .B(G176GAT), .Z(n437) );
  NAND2_X1 U493 ( .A1(G227GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U494 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U495 ( .A(n438), .B(G71GAT), .Z(n446) );
  XOR2_X1 U496 ( .A(G99GAT), .B(G134GAT), .Z(n440) );
  XNOR2_X1 U497 ( .A(G43GAT), .B(G190GAT), .ZN(n439) );
  XNOR2_X1 U498 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U499 ( .A(G120GAT), .B(KEYINPUT20), .Z(n442) );
  XNOR2_X1 U500 ( .A(G15GAT), .B(KEYINPUT80), .ZN(n441) );
  XNOR2_X1 U501 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U502 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U503 ( .A(n446), .B(n445), .ZN(n450) );
  XOR2_X1 U504 ( .A(n448), .B(n447), .Z(n449) );
  NAND2_X1 U505 ( .A1(n561), .A2(n328), .ZN(n454) );
  XOR2_X1 U506 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n452) );
  NAND2_X1 U507 ( .A1(n561), .A2(n554), .ZN(n456) );
  XNOR2_X1 U508 ( .A(KEYINPUT122), .B(G183GAT), .ZN(n455) );
  XNOR2_X1 U509 ( .A(n456), .B(n455), .ZN(G1350GAT) );
  XNOR2_X1 U510 ( .A(n457), .B(KEYINPUT101), .ZN(n533) );
  NAND2_X1 U511 ( .A1(n561), .A2(n533), .ZN(n463) );
  XOR2_X1 U512 ( .A(KEYINPUT121), .B(KEYINPUT120), .Z(n459) );
  XNOR2_X1 U513 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n458) );
  XOR2_X1 U514 ( .A(n459), .B(n458), .Z(n461) );
  XOR2_X1 U515 ( .A(G176GAT), .B(KEYINPUT119), .Z(n460) );
  XNOR2_X1 U516 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U517 ( .A(n463), .B(n462), .ZN(G1349GAT) );
  XOR2_X1 U518 ( .A(KEYINPUT97), .B(KEYINPUT34), .Z(n484) );
  INV_X1 U519 ( .A(n367), .ZN(n571) );
  NAND2_X1 U520 ( .A1(n560), .A2(n571), .ZN(n496) );
  NOR2_X1 U521 ( .A1(n328), .A2(n574), .ZN(n464) );
  XNOR2_X1 U522 ( .A(n464), .B(KEYINPUT16), .ZN(n482) );
  XOR2_X1 U523 ( .A(n472), .B(KEYINPUT28), .Z(n523) );
  XNOR2_X1 U524 ( .A(KEYINPUT27), .B(n520), .ZN(n475) );
  NAND2_X1 U525 ( .A1(n517), .A2(n475), .ZN(n544) );
  XOR2_X1 U526 ( .A(n527), .B(KEYINPUT93), .Z(n465) );
  INV_X1 U527 ( .A(n528), .ZN(n467) );
  NAND2_X1 U528 ( .A1(n465), .A2(n467), .ZN(n481) );
  NOR2_X1 U529 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U530 ( .A(KEYINPUT95), .B(n468), .ZN(n469) );
  NAND2_X1 U531 ( .A1(n469), .A2(n472), .ZN(n471) );
  XOR2_X1 U532 ( .A(KEYINPUT25), .B(KEYINPUT96), .Z(n470) );
  XNOR2_X1 U533 ( .A(n471), .B(n470), .ZN(n477) );
  XNOR2_X1 U534 ( .A(KEYINPUT94), .B(KEYINPUT26), .ZN(n474) );
  NOR2_X1 U535 ( .A1(n528), .A2(n472), .ZN(n473) );
  XNOR2_X1 U536 ( .A(n474), .B(n473), .ZN(n563) );
  NAND2_X1 U537 ( .A1(n475), .A2(n563), .ZN(n476) );
  NAND2_X1 U538 ( .A1(n477), .A2(n476), .ZN(n478) );
  NAND2_X1 U539 ( .A1(n479), .A2(n478), .ZN(n480) );
  NAND2_X1 U540 ( .A1(n482), .A2(n494), .ZN(n506) );
  NOR2_X1 U541 ( .A1(n496), .A2(n506), .ZN(n491) );
  NAND2_X1 U542 ( .A1(n491), .A2(n517), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U544 ( .A(G1GAT), .B(n485), .ZN(G1324GAT) );
  NAND2_X1 U545 ( .A1(n491), .A2(n520), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n486), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT35), .B(KEYINPUT99), .Z(n488) );
  NAND2_X1 U548 ( .A1(n491), .A2(n528), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(n490) );
  XOR2_X1 U550 ( .A(G15GAT), .B(KEYINPUT98), .Z(n489) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(G1326GAT) );
  NAND2_X1 U552 ( .A1(n491), .A2(n523), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n492), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U554 ( .A1(n554), .A2(n579), .ZN(n493) );
  NAND2_X1 U555 ( .A1(n494), .A2(n493), .ZN(n495) );
  XOR2_X1 U556 ( .A(KEYINPUT37), .B(n495), .Z(n516) );
  XOR2_X1 U557 ( .A(KEYINPUT38), .B(n497), .Z(n504) );
  NAND2_X1 U558 ( .A1(n517), .A2(n504), .ZN(n499) );
  XOR2_X1 U559 ( .A(KEYINPUT100), .B(KEYINPUT39), .Z(n498) );
  XNOR2_X1 U560 ( .A(G29GAT), .B(n500), .ZN(G1328GAT) );
  NAND2_X1 U561 ( .A1(n520), .A2(n504), .ZN(n501) );
  XNOR2_X1 U562 ( .A(G36GAT), .B(n501), .ZN(G1329GAT) );
  NAND2_X1 U563 ( .A1(n504), .A2(n528), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n502), .B(KEYINPUT40), .ZN(n503) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  NAND2_X1 U566 ( .A1(n504), .A2(n523), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n505), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n508) );
  NAND2_X1 U569 ( .A1(n565), .A2(n533), .ZN(n515) );
  NOR2_X1 U570 ( .A1(n515), .A2(n506), .ZN(n511) );
  NAND2_X1 U571 ( .A1(n517), .A2(n511), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n508), .B(n507), .ZN(G1332GAT) );
  NAND2_X1 U573 ( .A1(n511), .A2(n520), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n509), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U575 ( .A1(n511), .A2(n528), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n510), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT43), .B(KEYINPUT102), .Z(n513) );
  NAND2_X1 U578 ( .A1(n511), .A2(n523), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U580 ( .A(G78GAT), .B(n514), .ZN(G1335GAT) );
  XOR2_X1 U581 ( .A(G85GAT), .B(KEYINPUT103), .Z(n519) );
  NOR2_X1 U582 ( .A1(n516), .A2(n515), .ZN(n524) );
  NAND2_X1 U583 ( .A1(n524), .A2(n517), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n519), .B(n518), .ZN(G1336GAT) );
  NAND2_X1 U585 ( .A1(n524), .A2(n520), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n521), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U587 ( .A1(n524), .A2(n528), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n522), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U589 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n525), .B(KEYINPUT44), .ZN(n526) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  XOR2_X1 U592 ( .A(G113GAT), .B(KEYINPUT109), .Z(n532) );
  NAND2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U594 ( .A1(n545), .A2(n529), .ZN(n530) );
  XNOR2_X1 U595 ( .A(KEYINPUT108), .B(n530), .ZN(n540) );
  NAND2_X1 U596 ( .A1(n540), .A2(n560), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT111), .B(KEYINPUT49), .Z(n535) );
  NAND2_X1 U599 ( .A1(n540), .A2(n533), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n535), .B(n534), .ZN(n537) );
  XOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT110), .Z(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  NAND2_X1 U603 ( .A1(n540), .A2(n554), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n538), .B(KEYINPUT50), .ZN(n539) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n539), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT51), .B(KEYINPUT112), .Z(n542) );
  NAND2_X1 U607 ( .A1(n328), .A2(n540), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U609 ( .A(G134GAT), .B(n543), .ZN(G1343GAT) );
  NOR2_X1 U610 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U611 ( .A1(n546), .A2(n563), .ZN(n547) );
  XOR2_X1 U612 ( .A(n547), .B(KEYINPUT113), .Z(n551) );
  INV_X1 U613 ( .A(n551), .ZN(n557) );
  NAND2_X1 U614 ( .A1(n560), .A2(n557), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n548), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT52), .B(KEYINPUT114), .Z(n550) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n553) );
  NOR2_X1 U619 ( .A1(n457), .A2(n551), .ZN(n552) );
  XOR2_X1 U620 ( .A(n553), .B(n552), .Z(G1345GAT) );
  XOR2_X1 U621 ( .A(G155GAT), .B(KEYINPUT115), .Z(n556) );
  NAND2_X1 U622 ( .A1(n557), .A2(n554), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(G1346GAT) );
  NAND2_X1 U624 ( .A1(n557), .A2(n328), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(KEYINPUT116), .ZN(n559) );
  XNOR2_X1 U626 ( .A(G162GAT), .B(n559), .ZN(G1347GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(n562), .ZN(G1348GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n578) );
  NOR2_X1 U630 ( .A1(n565), .A2(n578), .ZN(n570) );
  XOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n567) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(KEYINPUT124), .B(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  NOR2_X1 U636 ( .A1(n571), .A2(n578), .ZN(n573) );
  XNOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n578), .ZN(n575) );
  XOR2_X1 U640 ( .A(G211GAT), .B(n575), .Z(G1354GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n577) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n581) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U645 ( .A(n581), .B(n580), .Z(G1355GAT) );
endmodule

