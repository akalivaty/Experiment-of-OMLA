//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 0 0 1 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 1 1 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n862, new_n863,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976;
  INV_X1    g000(.A(G227gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n207));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n207), .B1(new_n208), .B2(KEYINPUT65), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n210), .B(KEYINPUT23), .C1(G169gat), .C2(G176gat), .ZN(new_n211));
  AND2_X1   g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  AND2_X1   g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT24), .ZN(new_n214));
  AOI22_X1  g013(.A1(new_n213), .A2(new_n214), .B1(G169gat), .B2(G176gat), .ZN(new_n215));
  INV_X1    g014(.A(G183gat), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(KEYINPUT24), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n206), .B1(new_n212), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(KEYINPUT66), .A3(KEYINPUT25), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n209), .A2(new_n211), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(new_n220), .A3(new_n215), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n224), .B1(new_n226), .B2(new_n206), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT25), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n228), .B1(new_n226), .B2(new_n224), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n223), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n208), .A2(KEYINPUT26), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT26), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(G169gat), .B2(G176gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n213), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT28), .B1(new_n239), .B2(new_n217), .ZN(new_n240));
  OAI211_X1 g039(.A(KEYINPUT28), .B(new_n217), .C1(new_n237), .C2(new_n238), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n236), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT67), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n236), .B(new_n245), .C1(new_n240), .C2(new_n242), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n247), .ZN(new_n248));
  OR2_X1    g047(.A1(G127gat), .A2(G134gat), .ZN(new_n249));
  XOR2_X1   g048(.A(KEYINPUT68), .B(G127gat), .Z(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(G134gat), .ZN(new_n251));
  INV_X1    g050(.A(G120gat), .ZN(new_n252));
  OR2_X1    g051(.A1(new_n252), .A2(G113gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(G113gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(KEYINPUT69), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT69), .B1(new_n253), .B2(new_n254), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n249), .B(new_n251), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  XOR2_X1   g058(.A(KEYINPUT70), .B(G113gat), .Z(new_n260));
  OAI21_X1  g059(.A(new_n254), .B1(new_n260), .B2(new_n252), .ZN(new_n261));
  NAND2_X1  g060(.A1(G127gat), .A2(G134gat), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT1), .B1(new_n249), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n259), .A2(new_n264), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n230), .A2(new_n267), .A3(new_n247), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n205), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT71), .B1(new_n269), .B2(KEYINPUT33), .ZN(new_n270));
  XNOR2_X1  g069(.A(G71gat), .B(G99gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT72), .ZN(new_n272));
  XOR2_X1   g071(.A(G15gat), .B(G43gat), .Z(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n230), .A2(new_n267), .A3(new_n247), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n267), .B1(new_n230), .B2(new_n247), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n204), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n274), .B1(new_n277), .B2(KEYINPUT32), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT33), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n270), .A2(new_n278), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT73), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT73), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n270), .A2(new_n278), .A3(new_n284), .A4(new_n281), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n277), .A2(KEYINPUT32), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n274), .A2(new_n280), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT34), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n266), .A2(new_n268), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n293), .A2(new_n204), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT34), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n286), .A2(new_n295), .A3(new_n290), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n292), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n294), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n295), .B1(new_n286), .B2(new_n290), .ZN(new_n299));
  AOI211_X1 g098(.A(KEYINPUT34), .B(new_n289), .C1(new_n283), .C2(new_n285), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G78gat), .B(G106gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT31), .B(G50gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT78), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT2), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(G141gat), .B2(G148gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(G141gat), .A2(G148gat), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G155gat), .B(G162gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n306), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G141gat), .ZN(new_n314));
  INV_X1    g113(.A(G148gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n316), .A2(new_n307), .A3(new_n309), .ZN(new_n317));
  AND2_X1   g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(G155gat), .A2(G162gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n317), .A2(KEYINPUT78), .A3(new_n320), .ZN(new_n321));
  AND2_X1   g120(.A1(KEYINPUT79), .A2(G141gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(KEYINPUT79), .A2(G141gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT80), .B(G148gat), .ZN(new_n325));
  OAI22_X1  g124(.A1(new_n324), .A2(new_n315), .B1(new_n325), .B2(new_n314), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n319), .A2(new_n307), .ZN(new_n327));
  INV_X1    g126(.A(new_n318), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n313), .A2(new_n321), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(KEYINPUT74), .B(G211gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G218gat), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT22), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XOR2_X1   g134(.A(G211gat), .B(G218gat), .Z(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  XOR2_X1   g136(.A(G197gat), .B(G204gat), .Z(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n335), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT22), .B1(new_n332), .B2(G218gat), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n336), .B1(new_n341), .B2(new_n338), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT29), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n331), .B1(new_n343), .B2(KEYINPUT3), .ZN(new_n344));
  AND3_X1   g143(.A1(new_n344), .A2(G228gat), .A3(G233gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n340), .A2(new_n342), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n315), .A2(KEYINPUT80), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT80), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G148gat), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n314), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(new_n314), .ZN(new_n353));
  NAND2_X1  g152(.A1(KEYINPUT79), .A2(G141gat), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n315), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n329), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT3), .ZN(new_n357));
  NOR3_X1   g156(.A1(new_n311), .A2(new_n306), .A3(new_n312), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT78), .B1(new_n317), .B2(new_n320), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n356), .B(new_n357), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT81), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n313), .A2(new_n321), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n363), .A2(KEYINPUT81), .A3(new_n357), .A4(new_n356), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT29), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT83), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n347), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AOI211_X1 g166(.A(KEYINPUT83), .B(KEYINPUT29), .C1(new_n362), .C2(new_n364), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n345), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G228gat), .A2(G233gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n365), .A2(new_n346), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT82), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n340), .A2(new_n372), .A3(new_n342), .ZN(new_n373));
  OAI211_X1 g172(.A(KEYINPUT82), .B(new_n336), .C1(new_n341), .C2(new_n338), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n330), .B1(new_n376), .B2(new_n357), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n370), .B1(new_n371), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(G22gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n369), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n379), .B1(new_n369), .B2(new_n378), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n305), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT84), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g184(.A(KEYINPUT84), .B(new_n305), .C1(new_n381), .C2(new_n382), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT86), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n344), .A2(G228gat), .A3(G233gat), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT81), .B1(new_n330), .B2(new_n357), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n360), .A2(new_n361), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n375), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n346), .B1(new_n392), .B2(KEYINPUT83), .ZN(new_n393));
  INV_X1    g192(.A(new_n368), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n389), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n392), .A2(new_n347), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n376), .A2(new_n357), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n331), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n396), .A2(new_n398), .B1(G228gat), .B2(G233gat), .ZN(new_n399));
  OAI21_X1  g198(.A(G22gat), .B1(new_n395), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT85), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n400), .A2(new_n401), .A3(new_n380), .ZN(new_n402));
  OAI211_X1 g201(.A(KEYINPUT85), .B(G22gat), .C1(new_n395), .C2(new_n399), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n388), .B1(new_n404), .B2(new_n304), .ZN(new_n405));
  AOI211_X1 g204(.A(KEYINPUT86), .B(new_n305), .C1(new_n402), .C2(new_n403), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n387), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n297), .A2(new_n301), .A3(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G8gat), .B(G36gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(G92gat), .ZN(new_n410));
  XOR2_X1   g209(.A(KEYINPUT76), .B(G64gat), .Z(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT75), .ZN(new_n413));
  NAND2_X1  g212(.A1(G226gat), .A2(G233gat), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n230), .A2(new_n243), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n413), .B(new_n414), .C1(new_n415), .C2(KEYINPUT29), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT29), .B1(new_n230), .B2(new_n243), .ZN(new_n417));
  INV_X1    g216(.A(new_n414), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT75), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n248), .A2(new_n418), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n416), .A2(new_n346), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n418), .A2(KEYINPUT29), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n415), .A2(new_n418), .B1(new_n248), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n347), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n412), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT77), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n421), .A2(new_n424), .A3(new_n412), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n428), .B(KEYINPUT30), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n267), .B1(KEYINPUT3), .B2(new_n331), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n362), .A2(new_n364), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(G225gat), .A2(G233gat), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT4), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n435), .B1(new_n265), .B2(new_n331), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n267), .A2(KEYINPUT4), .A3(new_n330), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n433), .A2(new_n434), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT5), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n265), .B(new_n330), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n441), .A2(new_n434), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n437), .A2(new_n436), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n443), .B1(new_n432), .B2(new_n431), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n442), .B1(new_n444), .B2(new_n434), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n440), .B1(new_n445), .B2(new_n439), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT6), .ZN(new_n447));
  XNOR2_X1  g246(.A(G1gat), .B(G29gat), .ZN(new_n448));
  INV_X1    g247(.A(G85gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n448), .B(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT0), .B(G57gat), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n450), .B(new_n451), .Z(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n446), .A2(new_n447), .A3(new_n453), .ZN(new_n454));
  OAI211_X1 g253(.A(KEYINPUT90), .B(new_n440), .C1(new_n445), .C2(new_n439), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT90), .ZN(new_n456));
  INV_X1    g255(.A(new_n442), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n439), .B1(new_n438), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT5), .B1(new_n444), .B2(new_n434), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n456), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n455), .A2(new_n460), .A3(new_n452), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT6), .B1(new_n446), .B2(new_n453), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n454), .B1(new_n463), .B2(KEYINPUT91), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT91), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n461), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  AOI211_X1 g265(.A(KEYINPUT35), .B(new_n430), .C1(new_n464), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n408), .A2(new_n467), .ZN(new_n468));
  OR2_X1    g267(.A1(new_n446), .A2(new_n453), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n454), .B1(new_n462), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n470), .A2(new_n430), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n297), .A2(new_n301), .A3(new_n471), .A4(new_n407), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT35), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n461), .A2(KEYINPUT40), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n444), .A2(new_n434), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT39), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n452), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT89), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n441), .ZN(new_n482));
  INV_X1    g281(.A(new_n434), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n484), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT39), .B1(new_n486), .B2(new_n480), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n479), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n476), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT40), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n489), .B(new_n430), .C1(new_n490), .C2(new_n488), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n416), .A2(new_n347), .A3(new_n419), .A4(new_n420), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT37), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n493), .B1(new_n423), .B2(new_n346), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT38), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n412), .A2(new_n493), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n495), .B1(new_n425), .B2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(KEYINPUT92), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n464), .A2(new_n498), .A3(new_n428), .A4(new_n466), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n425), .A2(new_n496), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n493), .B1(new_n421), .B2(new_n424), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT38), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n502), .B(KEYINPUT93), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n407), .B(new_n491), .C1(new_n499), .C2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n471), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n380), .A2(new_n401), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n507), .A2(new_n382), .ZN(new_n508));
  INV_X1    g307(.A(new_n403), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n304), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT86), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n404), .A2(new_n388), .A3(new_n304), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT87), .B1(new_n513), .B2(new_n387), .ZN(new_n514));
  OAI211_X1 g313(.A(KEYINPUT87), .B(new_n387), .C1(new_n405), .C2(new_n406), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n506), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n297), .A2(new_n301), .A3(KEYINPUT36), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT36), .B1(new_n297), .B2(new_n301), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT88), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n505), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT36), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n294), .B1(new_n292), .B2(new_n296), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n299), .A2(new_n300), .A3(new_n298), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT87), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n407), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(new_n515), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n527), .A2(new_n518), .B1(new_n530), .B2(new_n506), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT88), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n475), .B1(new_n523), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G120gat), .B(G148gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(G176gat), .B(G204gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(G99gat), .ZN(new_n538));
  INV_X1    g337(.A(G106gat), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT8), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT7), .ZN(new_n541));
  INV_X1    g340(.A(G92gat), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n541), .B1(new_n449), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n540), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(KEYINPUT101), .B(G85gat), .Z(new_n546));
  AOI21_X1  g345(.A(new_n545), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G99gat), .B(G106gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT102), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n547), .A2(new_n548), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n551), .A2(KEYINPUT102), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT9), .ZN(new_n555));
  INV_X1    g354(.A(G71gat), .ZN(new_n556));
  INV_X1    g355(.A(G78gat), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n558), .A2(KEYINPUT100), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(KEYINPUT100), .ZN(new_n560));
  XNOR2_X1  g359(.A(G57gat), .B(G64gat), .ZN(new_n561));
  NOR3_X1   g360(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(G71gat), .B(G78gat), .Z(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n562), .A2(new_n564), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n554), .A2(KEYINPUT10), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n550), .A2(new_n567), .A3(new_n552), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n549), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n569), .B1(new_n572), .B2(KEYINPUT10), .ZN(new_n573));
  NAND2_X1  g372(.A1(G230gat), .A2(G233gat), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n574), .B(KEYINPUT104), .Z(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n570), .A2(new_n571), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n577), .A2(new_n574), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n537), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n579), .B(KEYINPUT105), .Z(new_n580));
  NAND2_X1  g379(.A1(new_n573), .A2(new_n574), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n581), .A2(new_n578), .A3(new_n537), .ZN(new_n582));
  AND2_X1   g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G15gat), .B(G22gat), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT16), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n584), .B1(new_n585), .B2(G1gat), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n586), .B1(G1gat), .B2(new_n584), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n587), .B(G8gat), .Z(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n568), .A2(KEYINPUT21), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n568), .A2(KEYINPUT21), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n592), .B1(new_n589), .B2(new_n590), .ZN(new_n593));
  NAND2_X1  g392(.A1(G231gat), .A2(G233gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(G183gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(G211gat), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n593), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G127gat), .B(G155gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n598), .B(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(G29gat), .A2(G36gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT14), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT95), .B(G36gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(G29gat), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n604), .B1(KEYINPUT97), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n607), .B1(KEYINPUT97), .B2(new_n606), .ZN(new_n608));
  XNOR2_X1  g407(.A(G43gat), .B(G50gat), .ZN(new_n609));
  OAI21_X1  g408(.A(KEYINPUT96), .B1(new_n609), .B2(KEYINPUT15), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(KEYINPUT15), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n604), .B1(G29gat), .B2(new_n605), .ZN(new_n613));
  OAI22_X1  g412(.A1(new_n608), .A2(new_n612), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT17), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n616), .B(KEYINPUT98), .Z(new_n617));
  OR2_X1    g416(.A1(new_n614), .A2(new_n615), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n553), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n554), .A2(new_n614), .ZN(new_n621));
  NAND3_X1  g420(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624));
  OAI22_X1  g423(.A1(new_n620), .A2(new_n623), .B1(KEYINPUT103), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(KEYINPUT103), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(G134gat), .B(G162gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n625), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n602), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n588), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n617), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G229gat), .A2(G233gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT99), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n589), .A2(new_n614), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT18), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n636), .A2(KEYINPUT18), .A3(new_n638), .A4(new_n639), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n614), .B(new_n588), .Z(new_n644));
  XOR2_X1   g443(.A(new_n638), .B(KEYINPUT13), .Z(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n642), .A2(new_n643), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G169gat), .B(G197gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(G113gat), .B(G141gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT94), .B(KEYINPUT11), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n652), .B(KEYINPUT12), .Z(new_n653));
  NAND2_X1  g452(.A1(new_n647), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n653), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n642), .A2(new_n655), .A3(new_n643), .A4(new_n646), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n583), .A2(new_n634), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(KEYINPUT106), .B1(new_n533), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n504), .B1(new_n531), .B2(KEYINPUT88), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n527), .A2(new_n518), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n661), .A2(KEYINPUT88), .A3(new_n517), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n474), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT106), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n654), .A2(new_n656), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n580), .A2(new_n582), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n663), .A2(new_n664), .A3(new_n667), .A4(new_n634), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n659), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n470), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g470(.A(KEYINPUT16), .B(G8gat), .Z(new_n672));
  NAND3_X1  g471(.A1(new_n669), .A2(new_n430), .A3(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(KEYINPUT42), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n669), .A2(new_n430), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n675), .B1(new_n676), .B2(G8gat), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n674), .B1(new_n673), .B2(new_n677), .ZN(G1325gat));
  NOR2_X1   g477(.A1(new_n525), .A2(new_n526), .ZN(new_n679));
  AOI21_X1  g478(.A(G15gat), .B1(new_n669), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n661), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n681), .A2(G15gat), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n680), .B1(new_n669), .B2(new_n682), .ZN(G1326gat));
  AOI21_X1  g482(.A(new_n379), .B1(new_n669), .B2(new_n530), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n669), .A2(new_n379), .A3(new_n530), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1327gat));
  INV_X1    g488(.A(new_n633), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n533), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n602), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n665), .A2(new_n666), .A3(new_n692), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(G29gat), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(new_n695), .A3(new_n470), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT108), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT44), .B1(new_n533), .B2(new_n690), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n504), .B(new_n517), .C1(new_n519), .C2(new_n520), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n474), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n633), .B(KEYINPUT109), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n700), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n693), .ZN(new_n708));
  INV_X1    g507(.A(new_n470), .ZN(new_n709));
  OAI21_X1  g508(.A(G29gat), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n696), .A2(KEYINPUT108), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n696), .A2(KEYINPUT108), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n711), .A2(new_n712), .A3(KEYINPUT45), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n699), .A2(new_n710), .A3(new_n713), .ZN(G1328gat));
  INV_X1    g513(.A(new_n430), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(new_n605), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n691), .A2(new_n693), .A3(new_n716), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(KEYINPUT46), .Z(new_n718));
  OAI21_X1  g517(.A(new_n605), .B1(new_n708), .B2(new_n715), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n718), .A2(KEYINPUT110), .A3(new_n719), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(G1329gat));
  OAI21_X1  g523(.A(G43gat), .B1(new_n708), .B2(new_n661), .ZN(new_n725));
  INV_X1    g524(.A(G43gat), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n694), .A2(new_n726), .A3(new_n679), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT47), .B1(new_n727), .B2(KEYINPUT111), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1330gat));
  INV_X1    g529(.A(new_n530), .ZN(new_n731));
  OAI21_X1  g530(.A(G50gat), .B1(new_n708), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n731), .A2(G50gat), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n694), .A2(new_n733), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n708), .A2(new_n407), .ZN(new_n736));
  INV_X1    g535(.A(G50gat), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n734), .A2(KEYINPUT48), .ZN(new_n739));
  OAI22_X1  g538(.A1(new_n735), .A2(KEYINPUT48), .B1(new_n738), .B2(new_n739), .ZN(G1331gat));
  NOR2_X1   g539(.A1(new_n583), .A2(new_n657), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n741), .A2(new_n634), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n702), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n470), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g545(.A1(new_n743), .A2(new_n715), .ZN(new_n747));
  NOR2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  AND2_X1   g547(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(new_n747), .B2(new_n748), .ZN(G1333gat));
  NAND3_X1  g550(.A1(new_n744), .A2(G71gat), .A3(new_n681), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n743), .A2(new_n526), .A3(new_n525), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n753), .B2(G71gat), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g554(.A1(new_n743), .A2(new_n731), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(new_n557), .ZN(G1335gat));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n602), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n758), .B1(new_n700), .B2(new_n706), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(new_n709), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n692), .A2(new_n657), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n702), .A2(new_n633), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AOI211_X1 g565(.A(new_n765), .B(new_n690), .C1(new_n701), .C2(new_n474), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT51), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n690), .B1(new_n701), .B2(new_n474), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n762), .B1(new_n770), .B2(KEYINPUT112), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n771), .A2(new_n772), .A3(new_n767), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n666), .A2(new_n470), .A3(new_n546), .ZN(new_n775));
  OAI22_X1  g574(.A1(new_n761), .A2(new_n546), .B1(new_n774), .B2(new_n775), .ZN(G1336gat));
  INV_X1    g575(.A(new_n758), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n703), .B1(new_n663), .B2(new_n633), .ZN(new_n778));
  INV_X1    g577(.A(new_n706), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n430), .B(new_n777), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G92gat), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n583), .A2(G92gat), .A3(new_n715), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n783), .B1(new_n769), .B2(new_n773), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n781), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n782), .B1(new_n781), .B2(new_n784), .ZN(new_n786));
  INV_X1    g585(.A(new_n783), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n766), .A2(KEYINPUT51), .A3(new_n768), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n772), .B1(new_n771), .B2(new_n767), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT52), .B1(new_n790), .B2(KEYINPUT113), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n785), .A2(new_n786), .A3(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n793), .B1(new_n784), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n542), .B1(new_n759), .B2(new_n430), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT114), .B1(new_n796), .B2(new_n790), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n781), .A2(new_n784), .A3(new_n782), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n795), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n792), .A2(new_n799), .ZN(G1337gat));
  OAI21_X1  g599(.A(G99gat), .B1(new_n760), .B2(new_n661), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n679), .A2(new_n538), .A3(new_n666), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(new_n774), .B2(new_n802), .ZN(G1338gat));
  INV_X1    g602(.A(new_n407), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n804), .A2(new_n666), .A3(new_n539), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n774), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(KEYINPUT53), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT115), .B1(new_n759), .B2(new_n804), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n759), .A2(KEYINPUT115), .A3(new_n804), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G106gat), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n807), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n539), .B1(new_n759), .B2(new_n530), .ZN(new_n812));
  OAI21_X1  g611(.A(KEYINPUT53), .B1(new_n806), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(G1339gat));
  NAND3_X1  g613(.A1(new_n583), .A2(new_n665), .A3(new_n634), .ZN(new_n815));
  XOR2_X1   g614(.A(new_n815), .B(KEYINPUT116), .Z(new_n816));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n536), .B1(new_n576), .B2(KEYINPUT54), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n820), .B1(new_n573), .B2(new_n574), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n822));
  INV_X1    g621(.A(new_n575), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n569), .B(new_n823), .C1(new_n572), .C2(KEYINPUT10), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n821), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n822), .B1(new_n821), .B2(new_n824), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n819), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n582), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n821), .A2(new_n824), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT117), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n818), .B1(new_n832), .B2(new_n825), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(KEYINPUT55), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n817), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n582), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n836), .B1(new_n833), .B2(KEYINPUT55), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n828), .A2(new_n829), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n837), .A2(KEYINPUT118), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n638), .B1(new_n636), .B2(new_n639), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n644), .A2(new_n645), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n652), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n840), .A2(new_n656), .A3(new_n705), .A4(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n666), .A2(new_n656), .A3(new_n843), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n846), .B1(new_n840), .B2(new_n657), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n844), .B1(new_n847), .B2(new_n705), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n816), .B1(new_n848), .B2(new_n602), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n709), .A2(new_n430), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n850), .A2(new_n679), .A3(new_n731), .A4(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(G113gat), .B1(new_n852), .B2(new_n665), .ZN(new_n853));
  INV_X1    g652(.A(new_n408), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n851), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n665), .A2(new_n260), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n853), .B1(new_n856), .B2(new_n857), .ZN(G1340gat));
  OAI21_X1  g657(.A(G120gat), .B1(new_n852), .B2(new_n583), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n666), .A2(new_n252), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n859), .B1(new_n856), .B2(new_n860), .ZN(G1341gat));
  INV_X1    g660(.A(new_n250), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n852), .A2(new_n862), .A3(new_n602), .ZN(new_n863));
  INV_X1    g662(.A(new_n856), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n692), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n863), .B1(new_n862), .B2(new_n865), .ZN(G1342gat));
  OR3_X1    g665(.A1(new_n856), .A2(G134gat), .A3(new_n690), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n867), .A2(KEYINPUT56), .ZN(new_n868));
  OAI21_X1  g667(.A(G134gat), .B1(new_n852), .B2(new_n690), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(KEYINPUT56), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(G1343gat));
  NAND2_X1  g670(.A1(new_n661), .A2(new_n851), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n849), .A2(new_n407), .A3(new_n872), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n873), .A2(new_n314), .A3(new_n657), .ZN(new_n874));
  OR3_X1    g673(.A1(new_n849), .A2(KEYINPUT57), .A3(new_n407), .ZN(new_n875));
  INV_X1    g674(.A(new_n872), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n833), .A2(KEYINPUT119), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n829), .B1(new_n833), .B2(KEYINPUT119), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n657), .B(new_n837), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n879), .A2(new_n845), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n844), .B1(new_n880), .B2(new_n633), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n816), .B1(new_n881), .B2(new_n602), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT57), .B1(new_n882), .B2(new_n731), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n875), .A2(new_n657), .A3(new_n876), .A4(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n874), .B1(new_n884), .B2(new_n324), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n886), .B1(new_n884), .B2(new_n324), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n885), .A2(new_n887), .A3(KEYINPUT58), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT58), .ZN(new_n889));
  AOI221_X4 g688(.A(new_n874), .B1(new_n886), .B2(new_n889), .C1(new_n884), .C2(new_n324), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n888), .A2(new_n890), .ZN(G1344gat));
  INV_X1    g690(.A(new_n325), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n873), .A2(new_n892), .A3(new_n666), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n875), .A2(new_n876), .A3(new_n883), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n894), .A2(new_n583), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n895), .A2(KEYINPUT59), .A3(new_n892), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT57), .B1(new_n849), .B2(new_n407), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n731), .A2(KEYINPUT57), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n633), .B1(new_n879), .B2(new_n845), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n633), .A2(new_n656), .A3(new_n843), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n830), .A2(new_n901), .A3(new_n834), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n602), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n903), .A2(new_n904), .A3(new_n815), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n903), .B2(new_n815), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n899), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n872), .A2(KEYINPUT121), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n583), .B1(new_n876), .B2(new_n909), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n898), .A2(new_n907), .A3(new_n908), .A4(new_n910), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n911), .A2(KEYINPUT123), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n315), .B1(new_n911), .B2(KEYINPUT123), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n897), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n893), .B1(new_n896), .B2(new_n914), .ZN(G1345gat));
  NAND2_X1  g714(.A1(new_n692), .A2(G155gat), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT124), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n894), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(G155gat), .B1(new_n873), .B2(new_n692), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(G1346gat));
  INV_X1    g719(.A(G162gat), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n894), .A2(new_n921), .A3(new_n704), .ZN(new_n922));
  AOI21_X1  g721(.A(G162gat), .B1(new_n873), .B2(new_n633), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n922), .A2(new_n923), .ZN(G1347gat));
  NAND2_X1  g723(.A1(new_n731), .A2(new_n679), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n715), .A2(new_n470), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n849), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(G169gat), .B1(new_n929), .B2(new_n665), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n855), .A2(new_n926), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n665), .A2(G169gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(G1348gat));
  INV_X1    g732(.A(new_n931), .ZN(new_n934));
  AOI21_X1  g733(.A(G176gat), .B1(new_n934), .B2(new_n666), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n666), .A2(G176gat), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n935), .B1(new_n928), .B2(new_n936), .ZN(G1349gat));
  NAND3_X1  g736(.A1(new_n934), .A2(new_n239), .A3(new_n692), .ZN(new_n938));
  OAI21_X1  g737(.A(G183gat), .B1(new_n929), .B2(new_n602), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g740(.A1(new_n934), .A2(new_n217), .A3(new_n705), .ZN(new_n942));
  OAI21_X1  g741(.A(G190gat), .B1(new_n929), .B2(new_n690), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n943), .A2(KEYINPUT61), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n943), .A2(KEYINPUT61), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(G1351gat));
  INV_X1    g745(.A(G197gat), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n898), .A2(new_n907), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n681), .A2(new_n927), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n947), .B1(new_n950), .B2(new_n657), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n849), .A2(new_n407), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(new_n949), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n953), .A2(G197gat), .A3(new_n665), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n951), .A2(new_n954), .ZN(G1352gat));
  OR2_X1    g754(.A1(new_n583), .A2(G204gat), .ZN(new_n956));
  OR3_X1    g755(.A1(new_n953), .A2(KEYINPUT62), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(KEYINPUT62), .B1(new_n953), .B2(new_n956), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n948), .A2(new_n666), .A3(new_n949), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT125), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g760(.A(G204gat), .B1(new_n959), .B2(new_n960), .ZN(new_n962));
  OAI211_X1 g761(.A(new_n957), .B(new_n958), .C1(new_n961), .C2(new_n962), .ZN(G1353gat));
  OR3_X1    g762(.A1(new_n953), .A2(new_n332), .A3(new_n602), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n898), .A2(new_n907), .A3(new_n692), .A4(new_n949), .ZN(new_n965));
  AND3_X1   g764(.A1(new_n965), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n966));
  AOI21_X1  g765(.A(KEYINPUT63), .B1(new_n965), .B2(G211gat), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n964), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT126), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI211_X1 g769(.A(KEYINPUT126), .B(new_n964), .C1(new_n966), .C2(new_n967), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(G1354gat));
  NAND2_X1  g771(.A1(new_n633), .A2(G218gat), .ZN(new_n973));
  XOR2_X1   g772(.A(new_n973), .B(KEYINPUT127), .Z(new_n974));
  NAND3_X1  g773(.A1(new_n952), .A2(new_n705), .A3(new_n949), .ZN(new_n975));
  INV_X1    g774(.A(G218gat), .ZN(new_n976));
  AOI22_X1  g775(.A1(new_n950), .A2(new_n974), .B1(new_n975), .B2(new_n976), .ZN(G1355gat));
endmodule


