//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1248, new_n1249,
    new_n1250, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n208), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(new_n201), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  INV_X1    g0025(.A(G244), .ZN(new_n226));
  INV_X1    g0026(.A(G107), .ZN(new_n227));
  INV_X1    g0027(.A(G264), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n225), .B1(new_n203), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n210), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n213), .B1(new_n216), .B2(new_n218), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT65), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT66), .ZN(new_n243));
  XOR2_X1   g0043(.A(G58), .B(G77), .Z(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n245), .B(new_n249), .ZN(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n214), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT8), .B(G58), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n208), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G150), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  OAI22_X1  g0057(.A1(new_n253), .A2(new_n254), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n208), .B1(new_n201), .B2(new_n202), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n252), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n260), .A2(KEYINPUT67), .B1(new_n202), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n252), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n261), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n265), .A2(KEYINPUT68), .B1(new_n207), .B2(G20), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(KEYINPUT68), .B2(new_n265), .ZN(new_n267));
  OAI221_X1 g0067(.A(new_n263), .B1(KEYINPUT67), .B2(new_n260), .C1(new_n267), .C2(new_n202), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT9), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT69), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT10), .ZN(new_n272));
  INV_X1    g0072(.A(G274), .ZN(new_n273));
  AND2_X1   g0073(.A1(G1), .A2(G13), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n274), .A2(new_n275), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n277), .ZN(new_n281));
  INV_X1    g0081(.A(G226), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n279), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT3), .B(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G222), .A2(G1698), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(G223), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n284), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(KEYINPUT3), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT3), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n280), .B1(new_n293), .B2(new_n203), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n283), .B1(new_n288), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G190), .ZN(new_n296));
  INV_X1    g0096(.A(G200), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n296), .B1(new_n297), .B2(new_n295), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n298), .B1(new_n268), .B2(new_n269), .ZN(new_n299));
  AND3_X1   g0099(.A1(new_n271), .A2(new_n272), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n272), .B1(new_n271), .B2(new_n299), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n295), .A2(G169), .ZN(new_n304));
  INV_X1    g0104(.A(G179), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n304), .B1(new_n305), .B2(new_n295), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n268), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT18), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT16), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT7), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(new_n284), .B2(G20), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n293), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n220), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT73), .ZN(new_n315));
  INV_X1    g0115(.A(G159), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n315), .B1(new_n257), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n256), .A2(KEYINPUT73), .A3(G159), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G58), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(new_n220), .ZN(new_n321));
  OAI21_X1  g0121(.A(G20), .B1(new_n321), .B2(new_n201), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n310), .B1(new_n314), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT72), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n289), .B2(KEYINPUT3), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n291), .A2(KEYINPUT72), .A3(G33), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n290), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n208), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n220), .B1(new_n329), .B2(KEYINPUT7), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(new_n311), .A3(new_n208), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n323), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n252), .B(new_n324), .C1(new_n334), .C2(new_n310), .ZN(new_n335));
  INV_X1    g0135(.A(new_n253), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n336), .A2(new_n262), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n337), .B1(new_n267), .B2(new_n336), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G232), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n279), .B1(new_n281), .B2(new_n341), .ZN(new_n342));
  AND2_X1   g0142(.A1(G33), .A2(G41), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n343), .A2(new_n214), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n282), .A2(G1698), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(G223), .B2(G1698), .ZN(new_n346));
  OAI22_X1  g0146(.A1(new_n328), .A2(new_n346), .B1(new_n289), .B2(new_n222), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n342), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G179), .ZN(new_n349));
  INV_X1    g0149(.A(G169), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n349), .B1(new_n350), .B2(new_n348), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n309), .B1(new_n340), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n342), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n347), .A2(new_n344), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n297), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G190), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n357), .A2(KEYINPUT74), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n357), .A2(KEYINPUT74), .ZN(new_n359));
  OR2_X1    g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n356), .B1(new_n348), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n335), .A2(new_n361), .A3(new_n339), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT17), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n340), .A2(new_n351), .A3(new_n309), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n362), .A2(new_n363), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n353), .A2(new_n364), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n256), .A2(G50), .B1(G20), .B2(new_n220), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n203), .B2(new_n254), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n252), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT11), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n369), .A2(KEYINPUT11), .A3(new_n252), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(KEYINPUT70), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n265), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n220), .B1(new_n207), .B2(G20), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT12), .B1(new_n261), .B2(G68), .ZN(new_n377));
  OR3_X1    g0177(.A1(new_n261), .A2(KEYINPUT12), .A3(G68), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n375), .A2(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT70), .B1(new_n372), .B2(new_n373), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n279), .B1(new_n281), .B2(new_n221), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT13), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n341), .A2(G1698), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n284), .B(new_n386), .C1(G226), .C2(G1698), .ZN(new_n387));
  NAND2_X1  g0187(.A1(G33), .A2(G97), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n384), .B(new_n385), .C1(new_n389), .C2(new_n280), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n280), .B1(new_n387), .B2(new_n388), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT13), .B1(new_n391), .B2(new_n383), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT14), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(new_n394), .A3(G169), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT71), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n350), .B1(new_n390), .B2(new_n392), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n398), .A2(KEYINPUT71), .A3(new_n394), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n398), .A2(new_n394), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n393), .A2(new_n305), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n382), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n382), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n393), .A2(new_n357), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n297), .B1(new_n390), .B2(new_n392), .ZN(new_n407));
  NOR3_X1   g0207(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n203), .B1(new_n207), .B2(G20), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n375), .A2(new_n410), .B1(new_n203), .B2(new_n262), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n253), .A2(new_n257), .B1(new_n208), .B2(new_n203), .ZN(new_n412));
  XNOR2_X1  g0212(.A(KEYINPUT15), .B(G87), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n413), .A2(new_n254), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n252), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n279), .B1(new_n281), .B2(new_n226), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n284), .A2(G238), .A3(G1698), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n284), .A2(G232), .A3(new_n286), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n418), .B(new_n419), .C1(new_n227), .C2(new_n284), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n417), .B1(new_n420), .B2(new_n344), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n416), .B1(new_n421), .B2(G190), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n297), .B2(new_n421), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n305), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n424), .B(new_n416), .C1(G169), .C2(new_n421), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n409), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NOR3_X1   g0226(.A1(new_n308), .A2(new_n367), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(G45), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(G1), .ZN(new_n429));
  NAND2_X1  g0229(.A1(KEYINPUT5), .A2(G41), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(KEYINPUT5), .A2(G41), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n429), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n433), .A2(G264), .A3(new_n280), .ZN(new_n434));
  OAI21_X1  g0234(.A(G274), .B1(new_n343), .B2(new_n214), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n433), .A2(new_n435), .A3(KEYINPUT76), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT76), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n207), .A2(G45), .ZN(new_n438));
  OR2_X1    g0238(.A1(KEYINPUT5), .A2(G41), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n438), .B1(new_n439), .B2(new_n430), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n437), .B1(new_n440), .B2(new_n276), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n434), .B1(new_n436), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(G250), .A2(G1698), .ZN(new_n443));
  INV_X1    g0243(.A(G257), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n443), .B1(new_n444), .B2(G1698), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n445), .A2(new_n290), .A3(new_n326), .A4(new_n327), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G33), .A2(G294), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n280), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT82), .B1(new_n442), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT76), .B1(new_n433), .B2(new_n435), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n440), .A2(new_n437), .A3(new_n276), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n439), .A2(new_n430), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n344), .B1(new_n429), .B2(new_n452), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n450), .A2(new_n451), .B1(new_n453), .B2(G264), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT82), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n444), .A2(G1698), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(G250), .B2(G1698), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n447), .B1(new_n328), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n344), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n454), .A2(new_n455), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n449), .A2(G169), .A3(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n442), .A2(new_n448), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G179), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n261), .A2(G107), .ZN(new_n465));
  XNOR2_X1  g0265(.A(new_n465), .B(KEYINPUT25), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n207), .A2(G33), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n264), .A2(KEYINPUT75), .A3(new_n261), .A4(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n261), .A2(new_n467), .A3(new_n214), .A4(new_n251), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT75), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n466), .B1(new_n472), .B2(new_n227), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT81), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT81), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n466), .B(new_n475), .C1(new_n472), .C2(new_n227), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT22), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n208), .A2(G87), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n478), .B1(new_n293), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G116), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(G20), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT23), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n208), .B2(G107), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n227), .A2(KEYINPUT23), .A3(G20), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n326), .A2(new_n327), .A3(new_n208), .A4(new_n290), .ZN(new_n487));
  NAND2_X1  g0287(.A1(KEYINPUT22), .A2(G87), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n480), .B(new_n486), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT24), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n264), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n487), .A2(new_n488), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n492), .A2(KEYINPUT24), .A3(new_n480), .A4(new_n486), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n477), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n464), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT83), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(G238), .A2(G1698), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n499), .B1(new_n226), .B2(G1698), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n500), .A2(new_n290), .A3(new_n326), .A4(new_n327), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n280), .B1(new_n501), .B2(new_n481), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n438), .A2(G250), .ZN(new_n503));
  OAI22_X1  g0303(.A1(new_n435), .A2(new_n438), .B1(new_n344), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(G200), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT19), .ZN(new_n506));
  INV_X1    g0306(.A(G97), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n222), .A2(new_n507), .A3(new_n227), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n388), .A2(new_n208), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AND4_X1   g0310(.A1(new_n506), .A2(new_n208), .A3(G33), .A4(G97), .ZN(new_n511));
  OAI22_X1  g0311(.A1(new_n510), .A2(new_n511), .B1(new_n487), .B2(new_n220), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n512), .A2(new_n252), .B1(new_n262), .B2(new_n413), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n468), .A2(new_n471), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G87), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n226), .A2(G1698), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(G238), .B2(G1698), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n481), .B1(new_n328), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n344), .ZN(new_n519));
  INV_X1    g0319(.A(new_n504), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(G190), .A3(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n505), .A2(new_n513), .A3(new_n515), .A4(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n487), .A2(new_n220), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n508), .A2(new_n509), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n511), .B1(new_n524), .B2(KEYINPUT19), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n252), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n413), .A2(new_n262), .ZN(new_n527));
  INV_X1    g0327(.A(new_n413), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n468), .A2(new_n471), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n350), .B1(new_n502), .B2(new_n504), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n504), .B1(new_n518), .B2(new_n344), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n305), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n522), .A2(new_n534), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n442), .A2(KEYINPUT82), .A3(new_n448), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n455), .B1(new_n454), .B2(new_n459), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n357), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n454), .A2(new_n459), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n297), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n474), .A2(new_n476), .B1(new_n491), .B2(new_n493), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n535), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n227), .B1(new_n312), .B2(new_n313), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n256), .A2(G77), .ZN(new_n545));
  NAND2_X1  g0345(.A1(KEYINPUT6), .A2(G97), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n546), .A2(G107), .ZN(new_n547));
  XNOR2_X1  g0347(.A(G97), .B(G107), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT6), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n545), .B1(new_n550), .B2(new_n208), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n252), .B1(new_n544), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n514), .A2(G97), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n262), .A2(new_n507), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n326), .A2(new_n290), .A3(new_n327), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n226), .A2(G1698), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT4), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n290), .A2(new_n292), .A3(G250), .A4(G1698), .ZN(new_n559));
  AND2_X1   g0359(.A1(KEYINPUT4), .A2(G244), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n290), .A2(new_n292), .A3(new_n560), .A4(new_n286), .ZN(new_n561));
  NAND2_X1  g0361(.A1(G33), .A2(G283), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n559), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n344), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n450), .A2(new_n451), .B1(new_n453), .B2(G257), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n305), .A3(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n563), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT4), .ZN(new_n568));
  INV_X1    g0368(.A(new_n557), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n568), .B1(new_n328), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n280), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n433), .A2(new_n280), .ZN(new_n572));
  OAI22_X1  g0372(.A1(new_n436), .A2(new_n441), .B1(new_n444), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n350), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n555), .A2(new_n566), .A3(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(KEYINPUT77), .B1(new_n571), .B2(new_n573), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT77), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n564), .A2(new_n577), .A3(new_n565), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(G200), .A3(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n571), .A2(new_n573), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n555), .B1(G190), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n575), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n461), .A2(new_n463), .B1(new_n477), .B2(new_n494), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT83), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n498), .A2(new_n543), .A3(new_n582), .A4(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(G116), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n251), .A2(new_n214), .B1(G20), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(G20), .B1(G33), .B2(G283), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n289), .A2(G97), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n588), .A2(new_n589), .A3(KEYINPUT78), .ZN(new_n590));
  AOI21_X1  g0390(.A(KEYINPUT78), .B1(new_n588), .B2(new_n589), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n587), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  XOR2_X1   g0392(.A(KEYINPUT79), .B(KEYINPUT20), .Z(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(KEYINPUT79), .A2(KEYINPUT20), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n587), .B(new_n595), .C1(new_n590), .C2(new_n591), .ZN(new_n596));
  MUX2_X1   g0396(.A(new_n261), .B(new_n469), .S(G116), .Z(new_n597));
  NAND3_X1  g0397(.A1(new_n594), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n228), .A2(G1698), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(G257), .B2(G1698), .ZN(new_n600));
  INV_X1    g0400(.A(G303), .ZN(new_n601));
  OAI22_X1  g0401(.A1(new_n328), .A2(new_n600), .B1(new_n601), .B2(new_n284), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n344), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n450), .A2(new_n451), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n453), .A2(G270), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n598), .A2(new_n606), .A3(G169), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT21), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n606), .A2(G200), .ZN(new_n610));
  INV_X1    g0410(.A(new_n598), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n450), .A2(new_n451), .B1(new_n453), .B2(G270), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n612), .A2(new_n360), .A3(new_n603), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n598), .A2(G179), .A3(new_n603), .A4(new_n612), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n598), .A2(new_n606), .A3(KEYINPUT21), .A4(G169), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n609), .A2(new_n614), .A3(new_n615), .A4(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT80), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n616), .A2(new_n615), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT80), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n619), .A2(new_n620), .A3(new_n609), .A4(new_n614), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n585), .A2(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n427), .A2(new_n623), .ZN(G372));
  INV_X1    g0424(.A(new_n307), .ZN(new_n625));
  XNOR2_X1  g0425(.A(new_n362), .B(KEYINPUT17), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n408), .A2(new_n425), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n626), .B1(new_n404), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n365), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n629), .A2(new_n352), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n625), .B1(new_n303), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n580), .A2(G190), .ZN(new_n634));
  INV_X1    g0434(.A(new_n555), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n579), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(G190), .B1(new_n449), .B2(new_n460), .ZN(new_n637));
  INV_X1    g0437(.A(new_n540), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n542), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n555), .A2(new_n574), .A3(new_n566), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n522), .A2(new_n534), .ZN(new_n641));
  AND4_X1   g0441(.A1(new_n636), .A2(new_n639), .A3(new_n640), .A4(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n609), .A2(new_n615), .A3(new_n616), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n496), .ZN(new_n645));
  AOI21_X1  g0445(.A(KEYINPUT84), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n639), .A2(new_n636), .A3(new_n640), .A4(new_n641), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n583), .A2(new_n643), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT84), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT85), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n641), .A2(new_n575), .A3(KEYINPUT26), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT26), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(new_n535), .B2(new_n640), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n651), .B1(new_n655), .B2(new_n534), .ZN(new_n656));
  INV_X1    g0456(.A(new_n534), .ZN(new_n657));
  AOI211_X1 g0457(.A(KEYINPUT85), .B(new_n657), .C1(new_n652), .C2(new_n654), .ZN(new_n658));
  OAI22_X1  g0458(.A1(new_n646), .A2(new_n650), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n633), .B1(new_n427), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT86), .ZN(G369));
  XNOR2_X1  g0461(.A(new_n583), .B(new_n497), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G213), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G343), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n644), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n662), .A2(new_n639), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n668), .B(KEYINPUT89), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n583), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(G330), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n618), .A2(new_n621), .ZN(new_n676));
  INV_X1    g0476(.A(new_n668), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n611), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT87), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n644), .A2(new_n679), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n680), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n678), .B1(new_n618), .B2(new_n621), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT87), .B1(new_n685), .B2(new_n682), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n675), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n662), .B(new_n639), .C1(new_n542), .C2(new_n677), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n583), .A2(new_n668), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(KEYINPUT88), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n691), .A2(KEYINPUT88), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n674), .B1(new_n693), .B2(new_n694), .ZN(G399));
  INV_X1    g0495(.A(new_n211), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G41), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n508), .A2(G116), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(G1), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n218), .B2(new_n698), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT28), .ZN(new_n702));
  AOI21_X1  g0502(.A(KEYINPUT26), .B1(new_n641), .B2(new_n575), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n535), .A2(new_n640), .A3(new_n653), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n534), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT85), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n655), .A2(new_n651), .A3(new_n534), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n645), .A2(new_n543), .A3(new_n582), .A4(KEYINPUT84), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n649), .B1(new_n647), .B2(new_n648), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n706), .A2(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n671), .ZN(new_n711));
  OAI21_X1  g0511(.A(KEYINPUT90), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT90), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n659), .A2(new_n713), .A3(new_n671), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT29), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n712), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n498), .A2(new_n584), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n642), .B1(new_n717), .B2(new_n643), .ZN(new_n718));
  XOR2_X1   g0518(.A(new_n534), .B(KEYINPUT91), .Z(new_n719));
  AOI21_X1  g0519(.A(new_n719), .B1(new_n654), .B2(new_n652), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n668), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n721), .A2(new_n715), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n662), .A2(new_n642), .A3(new_n676), .A4(new_n671), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  INV_X1    g0524(.A(new_n532), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n539), .A2(new_n725), .A3(new_n606), .A4(new_n305), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n580), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n532), .A2(new_n459), .A3(new_n434), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n603), .A2(new_n604), .A3(G179), .A4(new_n605), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n728), .A2(new_n730), .A3(new_n580), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT30), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n532), .A2(new_n459), .A3(new_n434), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(new_n729), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT30), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n734), .A2(new_n735), .A3(new_n580), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n727), .B1(new_n732), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n724), .B1(new_n737), .B2(new_n677), .ZN(new_n738));
  AND4_X1   g0538(.A1(new_n735), .A2(new_n728), .A3(new_n730), .A4(new_n580), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n735), .B1(new_n734), .B2(new_n580), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n739), .A2(new_n740), .B1(new_n580), .B2(new_n726), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(KEYINPUT31), .A3(new_n711), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n723), .A2(new_n738), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G330), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n716), .A2(new_n722), .A3(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n702), .B1(new_n746), .B2(G1), .ZN(G364));
  AOI21_X1  g0547(.A(new_n214), .B1(G20), .B2(new_n350), .ZN(new_n748));
  INV_X1    g0548(.A(new_n360), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n208), .A2(new_n305), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G200), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(new_n297), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(G190), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n752), .A2(G50), .B1(G77), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G179), .A2(G200), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n208), .B1(new_n756), .B2(G190), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G97), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n208), .A2(G179), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n760), .A2(new_n357), .A3(G200), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n755), .B(new_n759), .C1(new_n227), .C2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n760), .A2(G190), .A3(G200), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n222), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n293), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n751), .A2(G190), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n749), .A2(new_n753), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n765), .B1(new_n220), .B2(new_n767), .C1(new_n769), .C2(new_n320), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n756), .A2(G20), .A3(new_n357), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n316), .ZN(new_n772));
  XNOR2_X1  g0572(.A(KEYINPUT93), .B(KEYINPUT32), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n762), .A2(new_n770), .A3(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G322), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n769), .A2(new_n776), .B1(new_n601), .B2(new_n763), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n752), .A2(G326), .ZN(new_n778));
  INV_X1    g0578(.A(G311), .ZN(new_n779));
  INV_X1    g0579(.A(new_n754), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  XOR2_X1   g0581(.A(KEYINPUT33), .B(G317), .Z(new_n782));
  INV_X1    g0582(.A(G283), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n767), .A2(new_n782), .B1(new_n783), .B2(new_n761), .ZN(new_n784));
  INV_X1    g0584(.A(new_n771), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n284), .B1(new_n785), .B2(G329), .ZN(new_n786));
  INV_X1    g0586(.A(G294), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n786), .B1(new_n787), .B2(new_n757), .ZN(new_n788));
  NOR4_X1   g0588(.A1(new_n777), .A2(new_n781), .A3(new_n784), .A4(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n748), .B1(new_n775), .B2(new_n789), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n208), .A2(G13), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n207), .B1(new_n791), .B2(G45), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n697), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n211), .A2(G355), .A3(new_n284), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n245), .A2(new_n428), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n696), .A2(new_n556), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(G45), .B2(new_n218), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n796), .B1(G116), .B2(new_n211), .C1(new_n797), .C2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G13), .A2(G33), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT92), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(G20), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n748), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n795), .B1(new_n800), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n684), .A2(new_n686), .ZN(new_n806));
  INV_X1    g0606(.A(new_n803), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n790), .B(new_n805), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n806), .A2(G330), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n795), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n806), .A2(G330), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(G396));
  NAND2_X1  g0612(.A1(new_n416), .A2(new_n668), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n423), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n425), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n425), .A2(new_n668), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n671), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n659), .A2(new_n820), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n712), .A2(new_n714), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n822), .B2(new_n818), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n794), .B1(new_n823), .B2(new_n744), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n744), .B2(new_n823), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n748), .A2(new_n801), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n794), .B1(G77), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n328), .B1(G132), .B2(new_n785), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n768), .A2(G143), .B1(G150), .B2(new_n766), .ZN(new_n830));
  INV_X1    g0630(.A(G137), .ZN(new_n831));
  INV_X1    g0631(.A(new_n752), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n830), .B1(new_n831), .B2(new_n832), .C1(new_n316), .C2(new_n780), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT34), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n829), .B1(new_n320), .B2(new_n757), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  INV_X1    g0636(.A(new_n761), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(G68), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n202), .B2(new_n763), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT94), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n763), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n754), .A2(G116), .B1(new_n842), .B2(G107), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n843), .B1(new_n832), .B2(new_n601), .C1(new_n787), .C2(new_n769), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n766), .A2(G283), .B1(new_n837), .B2(G87), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n284), .B1(new_n785), .B2(G311), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n845), .A2(new_n759), .A3(new_n846), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n835), .A2(new_n841), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n828), .B1(new_n848), .B2(new_n748), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n818), .B2(new_n802), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n825), .A2(new_n850), .ZN(G384));
  XOR2_X1   g0651(.A(new_n550), .B(KEYINPUT95), .Z(new_n852));
  INV_X1    g0652(.A(KEYINPUT35), .ZN(new_n853));
  OAI211_X1 g0653(.A(G116), .B(new_n215), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(new_n853), .B2(new_n852), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT36), .ZN(new_n856));
  OR3_X1    g0656(.A1(new_n218), .A2(new_n203), .A3(new_n321), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n202), .A2(G68), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n207), .B(G13), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT38), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT37), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n340), .A2(new_n351), .ZN(new_n863));
  INV_X1    g0663(.A(new_n666), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n340), .A2(new_n864), .ZN(new_n865));
  AND4_X1   g0665(.A1(new_n862), .A2(new_n863), .A3(new_n865), .A4(new_n362), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n334), .A2(new_n310), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n323), .B1(new_n330), .B2(new_n331), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n264), .B1(new_n868), .B2(KEYINPUT16), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n339), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n871), .A2(KEYINPUT97), .A3(new_n864), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT97), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n338), .B1(new_n867), .B2(new_n869), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n873), .B1(new_n874), .B2(new_n666), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n871), .A2(new_n351), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n872), .A2(new_n875), .A3(new_n876), .A4(new_n362), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n866), .B1(KEYINPUT37), .B2(new_n877), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n630), .A2(new_n626), .B1(new_n875), .B2(new_n872), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n861), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n872), .A2(new_n875), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n367), .A2(new_n881), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n877), .A2(KEYINPUT37), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n882), .B(KEYINPUT38), .C1(new_n883), .C2(new_n866), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n405), .A2(new_n668), .ZN(new_n886));
  INV_X1    g0686(.A(new_n408), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n402), .B(new_n401), .C1(new_n397), .C2(new_n399), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n886), .B(new_n887), .C1(new_n888), .C2(new_n382), .ZN(new_n889));
  INV_X1    g0689(.A(new_n886), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n404), .B2(new_n408), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT96), .B1(new_n821), .B2(new_n816), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT96), .ZN(new_n894));
  INV_X1    g0694(.A(new_n816), .ZN(new_n895));
  AOI211_X1 g0695(.A(new_n894), .B(new_n895), .C1(new_n659), .C2(new_n820), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n885), .B(new_n892), .C1(new_n893), .C2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n404), .A2(new_n677), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n880), .A2(new_n884), .A3(KEYINPUT39), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n863), .A2(new_n865), .A3(new_n362), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(new_n862), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n865), .B1(new_n630), .B2(new_n626), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n861), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n904), .A2(new_n884), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n899), .B(new_n900), .C1(new_n905), .C2(KEYINPUT39), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n666), .B1(new_n629), .B2(new_n352), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n897), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n716), .A2(new_n722), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n633), .B1(new_n909), .B2(new_n427), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n908), .B(new_n910), .Z(new_n911));
  NAND3_X1  g0711(.A1(new_n741), .A2(KEYINPUT31), .A3(new_n668), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n738), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n723), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n427), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n817), .B1(new_n889), .B2(new_n891), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n914), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT40), .B1(new_n905), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n917), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT40), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n919), .A2(new_n885), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n915), .A2(new_n918), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n904), .A2(new_n884), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n920), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n916), .A2(new_n920), .A3(new_n914), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n884), .B2(new_n880), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n427), .B(new_n914), .C1(new_n924), .C2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n922), .A2(G330), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n911), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n207), .B2(new_n791), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n911), .A2(new_n928), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n860), .B1(new_n930), .B2(new_n931), .ZN(G367));
  OAI21_X1  g0732(.A(new_n804), .B1(new_n211), .B2(new_n413), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n798), .A2(new_n240), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n794), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n752), .A2(G143), .ZN(new_n936));
  OAI221_X1 g0736(.A(new_n936), .B1(new_n203), .B2(new_n761), .C1(new_n769), .C2(new_n255), .ZN(new_n937));
  AOI22_X1  g0737(.A1(G50), .A2(new_n754), .B1(new_n766), .B2(G159), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT102), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n284), .B1(new_n757), .B2(new_n220), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n763), .A2(new_n320), .B1(new_n831), .B2(new_n771), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT103), .ZN(new_n942));
  NOR4_X1   g0742(.A1(new_n937), .A2(new_n939), .A3(new_n940), .A4(new_n942), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n754), .A2(G283), .B1(new_n837), .B2(G97), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n944), .B1(new_n787), .B2(new_n767), .C1(new_n832), .C2(new_n779), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n556), .B1(G317), .B2(new_n785), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n946), .B1(new_n227), .B2(new_n757), .C1(new_n769), .C2(new_n601), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n763), .A2(new_n586), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT46), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n945), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n943), .A2(new_n950), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n951), .B(KEYINPUT47), .Z(new_n952));
  AOI21_X1  g0752(.A(new_n935), .B1(new_n952), .B2(new_n748), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n677), .B1(new_n513), .B2(new_n515), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n534), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n641), .B2(new_n954), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT98), .Z(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n953), .B1(new_n807), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n670), .B1(new_n690), .B2(new_n669), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n687), .A2(KEYINPUT100), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n687), .A2(KEYINPUT100), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n962), .A2(new_n960), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n965), .A2(new_n746), .A3(KEYINPUT101), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT44), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n636), .B(new_n640), .C1(new_n635), .C2(new_n671), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n575), .A2(new_n711), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n968), .A2(KEYINPUT99), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT99), .B1(new_n968), .B2(new_n969), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n967), .B1(new_n674), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n673), .A2(KEYINPUT44), .A3(new_n972), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n674), .A2(KEYINPUT45), .A3(new_n973), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT45), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n673), .B2(new_n972), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n976), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n694), .B2(new_n693), .ZN(new_n982));
  INV_X1    g0782(.A(new_n694), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n983), .A2(new_n976), .A3(new_n980), .A4(new_n692), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT101), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n963), .A2(new_n964), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n986), .B1(new_n987), .B2(new_n745), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n966), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n746), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n697), .B(KEYINPUT41), .Z(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n793), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n972), .A2(new_n670), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT42), .Z(new_n996));
  NAND2_X1  g0796(.A1(new_n973), .A2(new_n717), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n711), .B1(new_n997), .B2(new_n640), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n994), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1000), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n1002), .B(new_n994), .C1(new_n996), .C2(new_n998), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NOR3_X1   g0804(.A1(new_n693), .A2(new_n694), .A3(new_n972), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1004), .B(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n959), .B1(new_n993), .B2(new_n1007), .ZN(G387));
  NAND2_X1  g0808(.A1(new_n966), .A2(new_n988), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1009), .B(new_n697), .C1(new_n746), .C2(new_n965), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n688), .A2(new_n689), .A3(new_n803), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n748), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n768), .A2(G317), .B1(G303), .B2(new_n754), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n779), .B2(new_n767), .C1(new_n776), .C2(new_n832), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT48), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n842), .A2(G294), .B1(new_n758), .B2(G283), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT49), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n761), .A2(new_n586), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n556), .B(new_n1023), .C1(G326), .C2(new_n785), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n780), .A2(new_n220), .B1(new_n413), .B2(new_n757), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n203), .A2(new_n763), .B1(new_n761), .B2(new_n507), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n768), .A2(G50), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n752), .A2(G159), .B1(new_n336), .B2(new_n766), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n328), .B1(G150), .B2(new_n785), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1012), .B1(new_n1025), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n798), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n237), .B2(G45), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n699), .B(new_n428), .C1(new_n220), .C2(new_n203), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT104), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1039));
  OAI21_X1  g0839(.A(KEYINPUT50), .B1(new_n253), .B2(G50), .ZN(new_n1040));
  OR3_X1    g0840(.A1(new_n253), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1035), .B1(new_n1038), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n211), .A2(new_n284), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1043), .B1(G107), .B2(new_n211), .C1(new_n699), .C2(new_n1044), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n795), .B(new_n1033), .C1(new_n804), .C2(new_n1045), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n965), .A2(new_n793), .B1(new_n1011), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1010), .A2(new_n1047), .ZN(G393));
  NAND2_X1  g0848(.A1(new_n985), .A2(new_n793), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1034), .A2(new_n249), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n804), .B1(new_n507), .B2(new_n211), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n794), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G150), .A2(new_n752), .B1(new_n768), .B2(G159), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT51), .Z(new_n1054));
  NOR2_X1   g0854(.A1(new_n757), .A2(new_n203), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n780), .B2(new_n253), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G50), .B2(new_n766), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n220), .A2(new_n763), .B1(new_n761), .B2(new_n222), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n328), .B(new_n1059), .C1(G143), .C2(new_n785), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1054), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G311), .A2(new_n768), .B1(new_n752), .B2(G317), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT52), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n293), .B1(new_n771), .B2(new_n776), .C1(new_n761), .C2(new_n227), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n780), .A2(new_n787), .B1(new_n763), .B2(new_n783), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n766), .A2(G303), .B1(G116), .B2(new_n758), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1064), .B(new_n1065), .C1(KEYINPUT105), .C2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(KEYINPUT105), .B2(new_n1066), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1061), .B1(new_n1063), .B2(new_n1068), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT106), .Z(new_n1070));
  AOI21_X1  g0870(.A(new_n1052), .B1(new_n1070), .B2(new_n748), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n807), .B2(new_n973), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n989), .A2(new_n697), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n985), .B1(new_n966), .B2(new_n988), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1049), .B(new_n1072), .C1(new_n1073), .C2(new_n1074), .ZN(G390));
  AND2_X1   g0875(.A1(new_n768), .A2(G132), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n293), .B(new_n1076), .C1(G125), .C2(new_n785), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n763), .A2(new_n255), .ZN(new_n1078));
  XOR2_X1   g0878(.A(KEYINPUT109), .B(KEYINPUT53), .Z(new_n1079));
  XNOR2_X1  g0879(.A(new_n1078), .B(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(KEYINPUT54), .B(G143), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n780), .A2(new_n1081), .B1(new_n202), .B2(new_n761), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(G128), .B2(new_n752), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n766), .A2(G137), .B1(G159), .B2(new_n758), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1077), .A2(new_n1080), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G116), .A2(new_n768), .B1(new_n752), .B2(G283), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n284), .B(new_n764), .C1(G294), .C2(new_n785), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1086), .A2(new_n838), .A3(new_n1056), .A4(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G97), .A2(new_n754), .B1(new_n766), .B2(G107), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT110), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1085), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1012), .B1(new_n1091), .B2(KEYINPUT111), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(KEYINPUT111), .B2(new_n1091), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1093), .B(new_n794), .C1(new_n336), .C2(new_n827), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n900), .B1(new_n905), .B2(KEYINPUT39), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n802), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n675), .B1(new_n913), .B2(new_n723), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n916), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n880), .A2(new_n884), .A3(KEYINPUT39), .ZN(new_n1101));
  AOI21_X1  g0901(.A(KEYINPUT39), .B1(new_n904), .B2(new_n884), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n892), .B1(new_n893), .B2(new_n896), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1103), .B1(new_n1104), .B2(new_n898), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n895), .B1(new_n721), .B2(new_n815), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n892), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n923), .B(new_n898), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1100), .B1(new_n1105), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n706), .A2(new_n707), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n708), .A2(new_n709), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n819), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n894), .B1(new_n1113), .B2(new_n895), .ZN(new_n1114));
  OAI211_X1 g0914(.A(KEYINPUT96), .B(new_n816), .C1(new_n710), .C2(new_n819), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1107), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1095), .B1(new_n1116), .B2(new_n899), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n743), .A2(new_n892), .A3(G330), .A4(new_n818), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1117), .A2(new_n1108), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1110), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1097), .B1(new_n1121), .B2(new_n793), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n893), .A2(new_n896), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n743), .A2(G330), .A3(new_n818), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1124), .A2(new_n1107), .B1(new_n916), .B2(new_n1098), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n817), .B1(new_n1098), .B2(KEYINPUT107), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT107), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n738), .A2(new_n912), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n623), .B2(new_n671), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1127), .B1(new_n1129), .B2(new_n675), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n892), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1118), .A2(new_n1106), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n1123), .A2(new_n1125), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n427), .A2(new_n1098), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1133), .A2(new_n910), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n698), .B1(new_n1120), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n909), .A2(new_n427), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1137), .A2(new_n632), .A3(new_n1134), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1131), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1132), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1125), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1139), .A2(new_n1140), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1138), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1144), .A2(new_n1110), .A3(new_n1119), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n1136), .A2(KEYINPUT108), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT108), .B1(new_n1136), .B2(new_n1145), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1122), .B1(new_n1146), .B2(new_n1147), .ZN(G378));
  AOI21_X1  g0948(.A(new_n675), .B1(new_n918), .B2(new_n921), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n908), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(G330), .B1(new_n924), .B2(new_n926), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1151), .A2(new_n906), .A3(new_n907), .A4(new_n897), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n268), .A2(new_n864), .ZN(new_n1153));
  XOR2_X1   g0953(.A(new_n1153), .B(KEYINPUT112), .Z(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n303), .A2(new_n307), .A3(new_n1155), .ZN(new_n1156));
  XOR2_X1   g0956(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1157));
  NAND2_X1  g0957(.A1(new_n308), .A2(new_n1154), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1157), .B1(new_n1158), .B2(new_n1156), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1150), .A2(new_n1152), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1161), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1163));
  OAI21_X1  g0963(.A(KEYINPUT57), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n1117), .A2(new_n1108), .A3(new_n1118), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1099), .B1(new_n1117), .B2(new_n1108), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n1165), .A2(new_n1166), .A3(new_n1135), .ZN(new_n1167));
  OAI21_X1  g0967(.A(KEYINPUT113), .B1(new_n1167), .B2(new_n1138), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT113), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1138), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1145), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1164), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(KEYINPUT114), .B1(new_n1172), .B2(new_n698), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT57), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1163), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1150), .A2(new_n1152), .A3(new_n1161), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1174), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1145), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1169), .B1(new_n1145), .B2(new_n1170), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1177), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT114), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n1181), .A3(new_n697), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n1178), .A2(new_n1179), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n1174), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1173), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n793), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1161), .A2(new_n1096), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n556), .A2(G41), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n769), .A2(new_n227), .B1(new_n413), .B2(new_n780), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n767), .A2(new_n507), .B1(new_n320), .B2(new_n761), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n758), .A2(G68), .B1(new_n785), .B2(G283), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n752), .A2(G116), .B1(G77), .B2(new_n842), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1193), .A2(new_n1188), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1190), .B1(new_n1197), .B2(KEYINPUT58), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(KEYINPUT58), .B2(new_n1197), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G125), .A2(new_n752), .B1(new_n768), .B2(G128), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n754), .A2(G137), .B1(G150), .B2(new_n758), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1081), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n766), .A2(G132), .B1(new_n842), .B2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1200), .A2(new_n1201), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n837), .A2(G159), .ZN(new_n1206));
  AOI211_X1 g1006(.A(G33), .B(G41), .C1(new_n785), .C2(G124), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n748), .B1(new_n1199), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n795), .B1(new_n202), .B2(new_n826), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1187), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1186), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1185), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT115), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1215), .B(new_n1216), .ZN(G375));
  XOR2_X1   g1017(.A(new_n792), .B(KEYINPUT116), .Z(new_n1218));
  NOR2_X1   g1018(.A1(new_n1143), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1107), .A2(new_n801), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n794), .B1(G68), .B2(new_n827), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n1221), .B(KEYINPUT117), .Z(new_n1222));
  OAI22_X1  g1022(.A1(new_n783), .A2(new_n769), .B1(new_n832), .B2(new_n787), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n767), .A2(new_n586), .B1(new_n780), .B2(new_n227), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n293), .B1(new_n771), .B2(new_n601), .C1(new_n761), .C2(new_n203), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n763), .A2(new_n507), .B1(new_n757), .B2(new_n413), .ZN(new_n1226));
  OR4_X1    g1026(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n780), .A2(new_n255), .B1(new_n202), .B2(new_n757), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G159), .B2(new_n842), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n328), .B1(G128), .B2(new_n785), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n768), .A2(G137), .B1(G58), .B2(new_n837), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n752), .A2(G132), .B1(new_n766), .B2(new_n1202), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1227), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1222), .B1(new_n1234), .B2(new_n748), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1219), .B1(new_n1220), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1135), .A2(new_n992), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1170), .A2(new_n1133), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1236), .B1(new_n1237), .B2(new_n1238), .ZN(G381));
  NAND2_X1  g1039(.A1(new_n1136), .A2(new_n1145), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1240), .A2(new_n1122), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(G381), .A2(G384), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(G393), .A2(G396), .ZN(new_n1244));
  INV_X1    g1044(.A(G390), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  OR4_X1    g1046(.A1(G387), .A2(G375), .A3(new_n1242), .A4(new_n1246), .ZN(G407));
  NAND2_X1  g1047(.A1(new_n667), .A2(G213), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1241), .A2(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(G407), .B(G213), .C1(G375), .C2(new_n1250), .ZN(G409));
  NAND2_X1  g1051(.A1(G387), .A2(new_n1245), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(KEYINPUT122), .ZN(new_n1253));
  OR2_X1    g1053(.A1(new_n993), .A2(new_n1007), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1254), .A2(KEYINPUT121), .A3(new_n959), .A4(G390), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT122), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(G387), .A2(new_n1245), .A3(new_n1256), .ZN(new_n1257));
  OAI211_X1 g1057(.A(G390), .B(new_n959), .C1(new_n993), .C2(new_n1007), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT121), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1253), .A2(new_n1255), .A3(new_n1257), .A4(new_n1260), .ZN(new_n1261));
  XOR2_X1   g1061(.A(G393), .B(G396), .Z(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1262), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(new_n1252), .A3(new_n1258), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT61), .B1(new_n1263), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1249), .A2(G2897), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1238), .B1(KEYINPUT60), .B2(new_n1135), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1138), .A2(new_n1143), .A3(KEYINPUT60), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n697), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1236), .B1(new_n1269), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(G384), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT119), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1274), .B(new_n1275), .ZN(new_n1276));
  OAI211_X1 g1076(.A(G384), .B(new_n1236), .C1(new_n1269), .C2(new_n1271), .ZN(new_n1277));
  XOR2_X1   g1077(.A(new_n1277), .B(KEYINPUT118), .Z(new_n1278));
  OAI21_X1  g1078(.A(new_n1268), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1274), .B(KEYINPUT119), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1277), .B(KEYINPUT118), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1280), .A2(new_n1281), .A3(new_n1267), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1279), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1185), .A2(G378), .A3(new_n1214), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1285));
  OAI221_X1 g1085(.A(new_n1213), .B1(new_n1285), .B2(new_n1218), .C1(new_n1183), .C2(new_n991), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1241), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1249), .B1(new_n1284), .B2(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1266), .B1(new_n1283), .B2(new_n1288), .ZN(new_n1289));
  XOR2_X1   g1089(.A(KEYINPUT120), .B(KEYINPUT63), .Z(new_n1290));
  NOR2_X1   g1090(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1290), .B1(new_n1288), .B2(new_n1291), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1289), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT123), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1284), .A2(new_n1287), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1294), .B1(new_n1295), .B2(new_n1248), .ZN(new_n1296));
  AOI211_X1 g1096(.A(KEYINPUT123), .B(new_n1249), .C1(new_n1284), .C2(new_n1287), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1291), .A2(KEYINPUT63), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1296), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1293), .B1(new_n1299), .B2(KEYINPUT124), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1295), .A2(new_n1248), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(KEYINPUT123), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1288), .A2(new_n1294), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1298), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1302), .A2(new_n1303), .A3(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT124), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  OAI21_X1  g1107(.A(KEYINPUT125), .B1(new_n1300), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1299), .A2(KEYINPUT124), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT125), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1309), .A2(new_n1310), .A3(new_n1311), .A4(new_n1293), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1308), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT126), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1283), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1314), .B1(new_n1315), .B2(KEYINPUT61), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT61), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1318));
  OAI211_X1 g1118(.A(KEYINPUT126), .B(new_n1317), .C1(new_n1318), .C2(new_n1283), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1302), .A2(KEYINPUT62), .A3(new_n1303), .A4(new_n1291), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT62), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1291), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1321), .B1(new_n1301), .B2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1320), .A2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1316), .A2(new_n1319), .A3(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1313), .A2(new_n1328), .ZN(G405));
  INV_X1    g1129(.A(KEYINPUT127), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1284), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1331), .B1(G375), .B2(new_n1241), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1322), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1333), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1332), .A2(new_n1322), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1330), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  OR2_X1    g1136(.A1(new_n1332), .A2(new_n1322), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1337), .A2(KEYINPUT127), .A3(new_n1333), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1336), .A2(new_n1338), .A3(new_n1326), .ZN(new_n1339));
  OAI211_X1 g1139(.A(new_n1330), .B(new_n1327), .C1(new_n1334), .C2(new_n1335), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1339), .A2(new_n1340), .ZN(G402));
endmodule


