//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 1 1 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1007, new_n1008, new_n1009, new_n1010, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G113), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT5), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n189), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(KEYINPUT66), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT66), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G116), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n196), .A3(G119), .ZN(new_n197));
  INV_X1    g011(.A(new_n191), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n193), .B1(new_n199), .B2(new_n192), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G116), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n191), .B1(new_n201), .B2(G119), .ZN(new_n202));
  XOR2_X1   g016(.A(KEYINPUT2), .B(G113), .Z(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(G107), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(G107), .ZN(new_n208));
  AOI22_X1  g022(.A1(new_n206), .A2(new_n207), .B1(new_n208), .B2(KEYINPUT81), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  INV_X1    g024(.A(G107), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G104), .ZN(new_n212));
  INV_X1    g026(.A(new_n207), .ZN(new_n213));
  NOR2_X1   g027(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT81), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(new_n205), .A3(G107), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n209), .A2(new_n210), .A3(new_n215), .A4(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n210), .B1(new_n212), .B2(new_n208), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n200), .A2(new_n204), .A3(new_n218), .A4(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n207), .A2(G104), .A3(new_n211), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT81), .B1(new_n211), .B2(G104), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n223), .A3(new_n217), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT80), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n227), .A2(new_n207), .B1(G104), .B2(new_n211), .ZN(new_n228));
  OAI21_X1  g042(.A(G101), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n218), .A2(new_n229), .A3(KEYINPUT4), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n231), .B(G101), .C1(new_n224), .C2(new_n228), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n202), .A2(new_n203), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n203), .A2(new_n197), .A3(new_n198), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n221), .B1(new_n230), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(G110), .B(G122), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n237), .B(new_n221), .C1(new_n230), .C2(new_n235), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(KEYINPUT6), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G953), .ZN(new_n242));
  INV_X1    g056(.A(G143), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G146), .ZN(new_n244));
  INV_X1    g058(.A(G128), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n244), .B1(KEYINPUT1), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(G143), .B(G146), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n246), .B1(new_n247), .B2(KEYINPUT1), .ZN(new_n248));
  INV_X1    g062(.A(G146), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G143), .ZN(new_n250));
  AOI21_X1  g064(.A(G128), .B1(new_n250), .B2(new_n244), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(G125), .B1(new_n248), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G125), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n243), .A2(G146), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n249), .A2(G143), .ZN(new_n256));
  NAND2_X1  g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(KEYINPUT0), .A2(G128), .ZN(new_n259));
  OAI22_X1  g073(.A1(new_n255), .A2(new_n256), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n250), .A2(new_n244), .A3(new_n257), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n254), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OAI211_X1 g076(.A(G224), .B(new_n242), .C1(new_n253), .C2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(KEYINPUT1), .B1(new_n250), .B2(new_n244), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT1), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n265), .A2(G128), .B1(new_n243), .B2(G146), .ZN(new_n266));
  OAI22_X1  g080(.A1(new_n264), .A2(new_n266), .B1(G128), .B2(new_n247), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n254), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n260), .A2(new_n261), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G125), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n242), .A2(G224), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n268), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n263), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n236), .A2(new_n274), .A3(new_n238), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n241), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n237), .B(KEYINPUT8), .ZN(new_n277));
  INV_X1    g091(.A(new_n221), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n200), .A2(new_n204), .B1(new_n218), .B2(new_n220), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OR2_X1    g094(.A1(new_n272), .A2(KEYINPUT7), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT7), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n271), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n263), .A2(new_n272), .A3(new_n283), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n280), .A2(new_n240), .A3(new_n281), .A4(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G902), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n188), .B1(new_n276), .B2(new_n287), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n285), .A2(new_n286), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n241), .A2(new_n273), .A3(new_n275), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(new_n290), .A3(new_n187), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G475), .ZN(new_n293));
  NOR2_X1   g107(.A1(G237), .A2(G953), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G214), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(KEYINPUT85), .A3(G143), .ZN(new_n296));
  OR2_X1    g110(.A1(KEYINPUT85), .A2(G143), .ZN(new_n297));
  NAND2_X1  g111(.A1(KEYINPUT85), .A2(G143), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n297), .A2(G214), .A3(new_n294), .A4(new_n298), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n296), .A2(G131), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(G131), .B1(new_n296), .B2(new_n299), .ZN(new_n301));
  NOR3_X1   g115(.A1(new_n300), .A2(new_n301), .A3(KEYINPUT17), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n296), .A2(new_n299), .A3(KEYINPUT17), .A4(G131), .ZN(new_n303));
  INV_X1    g117(.A(G140), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G125), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n254), .A2(G140), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT16), .ZN(new_n307));
  OR3_X1    g121(.A1(new_n254), .A2(KEYINPUT16), .A3(G140), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n249), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n307), .A2(new_n308), .A3(G146), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n303), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT86), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n313), .B1(new_n296), .B2(new_n299), .ZN(new_n314));
  NAND2_X1  g128(.A1(KEYINPUT18), .A2(G131), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n305), .A2(new_n306), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G146), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n305), .A2(new_n306), .A3(new_n249), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n321), .B1(new_n314), .B2(new_n315), .ZN(new_n322));
  OAI22_X1  g136(.A1(new_n302), .A2(new_n312), .B1(new_n317), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(G113), .B(G122), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(new_n205), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n303), .A2(new_n310), .A3(new_n311), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n296), .A2(new_n299), .ZN(new_n329));
  INV_X1    g143(.A(G131), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT17), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n296), .A2(G131), .A3(new_n299), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n328), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n329), .A2(KEYINPUT86), .ZN(new_n336));
  INV_X1    g150(.A(new_n315), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(new_n316), .A3(new_n321), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n335), .A2(new_n339), .A3(new_n325), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n327), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n293), .B1(new_n341), .B2(new_n286), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT19), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT19), .B1(new_n305), .B2(new_n306), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n249), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n345), .B(new_n311), .C1(new_n300), .C2(new_n301), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n346), .B1(new_n317), .B2(new_n322), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n326), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n340), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT20), .ZN(new_n350));
  NOR2_X1   g164(.A1(G475), .A2(G902), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n350), .B1(new_n349), .B2(new_n351), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT87), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n349), .A2(KEYINPUT87), .A3(new_n350), .A4(new_n351), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n342), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(G214), .B1(G237), .B2(G902), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(KEYINPUT84), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G478), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(KEYINPUT15), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n243), .A2(G128), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n245), .A2(KEYINPUT88), .A3(G143), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT88), .B1(new_n245), .B2(G143), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G134), .ZN(new_n368));
  INV_X1    g182(.A(G134), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n369), .B(new_n364), .C1(new_n365), .C2(new_n366), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n201), .A2(KEYINPUT14), .A3(G122), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n194), .A2(new_n196), .A3(G122), .ZN(new_n373));
  OR2_X1    g187(.A1(new_n190), .A2(G122), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g189(.A(G107), .B(new_n372), .C1(new_n375), .C2(KEYINPUT14), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n373), .A2(new_n211), .A3(new_n374), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n371), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT13), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n379), .B1(new_n365), .B2(new_n366), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n367), .A2(new_n380), .A3(G134), .ZN(new_n381));
  OAI221_X1 g195(.A(new_n364), .B1(new_n379), .B2(new_n369), .C1(new_n365), .C2(new_n366), .ZN(new_n382));
  INV_X1    g196(.A(new_n377), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n211), .B1(new_n373), .B2(new_n374), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n381), .B(new_n382), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(KEYINPUT9), .B(G234), .ZN(new_n386));
  INV_X1    g200(.A(G217), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n386), .A2(new_n387), .A3(G953), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n378), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n388), .B1(new_n378), .B2(new_n385), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n286), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT89), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT89), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n393), .B(new_n286), .C1(new_n389), .C2(new_n390), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n363), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n242), .A2(G952), .ZN(new_n396));
  NAND2_X1  g210(.A1(G234), .A2(G237), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n397), .A2(G902), .A3(G953), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(KEYINPUT21), .B(G898), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n399), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n378), .A2(new_n385), .ZN(new_n404));
  INV_X1    g218(.A(new_n388), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n378), .A2(new_n385), .A3(new_n388), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(new_n286), .A3(new_n363), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NOR3_X1   g224(.A1(new_n395), .A2(new_n403), .A3(new_n410), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n292), .A2(new_n357), .A3(new_n360), .A4(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(G221), .B1(new_n386), .B2(G902), .ZN(new_n413));
  XNOR2_X1  g227(.A(G110), .B(G140), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n242), .A2(G227), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n414), .B(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n218), .A2(new_n229), .A3(KEYINPUT4), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(new_n269), .A3(new_n232), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n219), .B1(new_n248), .B2(new_n252), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n420), .A2(KEYINPUT10), .A3(new_n218), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n218), .A2(new_n267), .A3(new_n220), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n419), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT11), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n426), .B1(new_n369), .B2(G137), .ZN(new_n427));
  INV_X1    g241(.A(G137), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(KEYINPUT11), .A3(G134), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n369), .A2(G137), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n427), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G131), .ZN(new_n432));
  AOI21_X1  g246(.A(G131), .B1(new_n369), .B2(G137), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n427), .A2(new_n433), .A3(new_n429), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n425), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n435), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n419), .A2(new_n437), .A3(new_n421), .A4(new_n424), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n417), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n417), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT83), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n265), .B1(new_n255), .B2(new_n256), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n251), .B1(new_n442), .B2(new_n246), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n224), .A2(new_n228), .A3(G101), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n443), .B1(new_n444), .B2(new_n219), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n422), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(KEYINPUT12), .A3(new_n435), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT12), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n218), .A2(new_n220), .ZN(new_n449));
  AOI22_X1  g263(.A1(new_n449), .A2(new_n443), .B1(new_n420), .B2(new_n218), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n448), .B1(new_n450), .B2(new_n437), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n440), .A2(new_n441), .B1(new_n447), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n438), .A2(KEYINPUT83), .A3(new_n417), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n439), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n454), .A2(G469), .A3(G902), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n451), .A2(new_n447), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n438), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n416), .ZN(new_n458));
  INV_X1    g272(.A(new_n440), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n436), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n458), .A2(G469), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G469), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(new_n286), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n413), .B1(new_n455), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n412), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G210), .ZN(new_n469));
  NOR3_X1   g283(.A1(new_n469), .A2(G237), .A3(G953), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT27), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(KEYINPUT26), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(new_n210), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT28), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n369), .A2(G137), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n428), .A2(G134), .ZN(new_n477));
  OAI21_X1  g291(.A(G131), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n478), .A2(new_n434), .A3(KEYINPUT67), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT67), .B1(new_n478), .B2(new_n434), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n267), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT68), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT68), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n483), .B(new_n267), .C1(new_n479), .C2(new_n480), .ZN(new_n484));
  INV_X1    g298(.A(new_n203), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n199), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n204), .A2(new_n486), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n432), .A2(new_n434), .B1(new_n260), .B2(new_n261), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n482), .A2(new_n484), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT0), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n245), .ZN(new_n492));
  AOI22_X1  g306(.A1(new_n250), .A2(new_n244), .B1(new_n492), .B2(new_n257), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n250), .A2(new_n244), .A3(new_n257), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT64), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT64), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n260), .A2(new_n496), .A3(new_n261), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n435), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT65), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n478), .A2(new_n434), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n499), .B1(new_n443), .B2(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n267), .A2(KEYINPUT65), .A3(new_n434), .A4(new_n478), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n498), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n487), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n475), .B1(new_n490), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT28), .B1(new_n489), .B2(new_n481), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n474), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT70), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT70), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n474), .B(new_n509), .C1(new_n505), .C2(new_n506), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT30), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n488), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n482), .A2(new_n484), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n503), .A2(new_n512), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n487), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(new_n490), .A3(new_n473), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT69), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT31), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT31), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n516), .A2(new_n520), .A3(new_n490), .A4(new_n473), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n518), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n517), .A2(KEYINPUT31), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n511), .A2(new_n519), .A3(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(G472), .A2(G902), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(KEYINPUT32), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n516), .A2(new_n490), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n528), .A2(new_n473), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT29), .ZN(new_n530));
  AOI21_X1  g344(.A(G902), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OR2_X1    g345(.A1(new_n505), .A2(new_n506), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n473), .B1(new_n532), .B2(KEYINPUT29), .ZN(new_n533));
  INV_X1    g347(.A(new_n488), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n482), .A2(new_n484), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n487), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n490), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT28), .ZN(new_n538));
  XOR2_X1   g352(.A(new_n506), .B(KEYINPUT73), .Z(new_n539));
  AOI21_X1  g353(.A(new_n530), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n531), .B1(new_n533), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(G472), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n527), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT72), .ZN(new_n544));
  INV_X1    g358(.A(new_n526), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n508), .A2(new_n510), .B1(new_n522), .B2(new_n523), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n545), .B1(new_n546), .B2(new_n519), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT71), .B(KEYINPUT32), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n544), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n525), .A2(new_n526), .ZN(new_n550));
  INV_X1    g364(.A(new_n548), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(KEYINPUT72), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n543), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n242), .A2(G221), .A3(G234), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT22), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n428), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n554), .A2(KEYINPUT22), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n554), .A2(KEYINPUT22), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n557), .A2(G137), .A3(new_n558), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT74), .ZN(new_n562));
  INV_X1    g376(.A(G119), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n563), .A3(G128), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n245), .A2(G119), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  XOR2_X1   g380(.A(KEYINPUT24), .B(G110), .Z(new_n567));
  OAI21_X1  g381(.A(KEYINPUT74), .B1(new_n245), .B2(G119), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n566), .A2(KEYINPUT75), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT75), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(new_n564), .A3(new_n565), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT24), .B(G110), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n307), .A2(G146), .A3(new_n308), .ZN(new_n574));
  AOI21_X1  g388(.A(G146), .B1(new_n307), .B2(new_n308), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n569), .B(new_n573), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(G110), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT23), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n563), .B2(G128), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n245), .A2(KEYINPUT23), .A3(G119), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n563), .A2(G128), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT76), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n577), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n579), .A2(new_n580), .A3(KEYINPUT76), .A4(new_n581), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n576), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n311), .A2(new_n320), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n579), .A2(new_n580), .A3(new_n577), .A4(new_n581), .ZN(new_n589));
  AOI22_X1  g403(.A1(KEYINPUT77), .A2(new_n589), .B1(new_n571), .B2(new_n572), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n589), .A2(KEYINPUT77), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n561), .B1(new_n587), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n590), .A2(new_n591), .ZN(new_n594));
  INV_X1    g408(.A(new_n588), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n596), .B(new_n560), .C1(new_n586), .C2(new_n576), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n593), .A2(new_n286), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT25), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT25), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n593), .A2(new_n600), .A3(new_n597), .A4(new_n286), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n387), .B1(G234), .B2(new_n286), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n593), .A2(new_n597), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n602), .A2(G902), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT78), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n603), .A2(KEYINPUT78), .A3(new_n606), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(KEYINPUT79), .B1(new_n553), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g426(.A1(new_n547), .A2(KEYINPUT32), .B1(G472), .B2(new_n541), .ZN(new_n613));
  AOI21_X1  g427(.A(KEYINPUT72), .B1(new_n550), .B2(new_n551), .ZN(new_n614));
  AOI211_X1 g428(.A(new_n544), .B(new_n548), .C1(new_n525), .C2(new_n526), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT79), .ZN(new_n617));
  INV_X1    g431(.A(new_n611), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n468), .B1(new_n612), .B2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(new_n210), .ZN(G3));
  NAND2_X1  g435(.A1(new_n525), .A2(new_n286), .ZN(new_n622));
  AOI22_X1  g436(.A1(new_n622), .A2(G472), .B1(new_n526), .B2(new_n525), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n466), .A2(new_n611), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n359), .B1(new_n288), .B2(new_n291), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n393), .B1(new_n408), .B2(new_n286), .ZN(new_n627));
  INV_X1    g441(.A(new_n394), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n361), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT33), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n630), .B1(new_n389), .B2(new_n390), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n406), .A2(KEYINPUT33), .A3(new_n407), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n286), .A2(G478), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n629), .B(KEYINPUT90), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT90), .ZN(new_n636));
  AOI21_X1  g450(.A(G478), .B1(new_n392), .B2(new_n394), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n633), .A2(new_n634), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n357), .ZN(new_n641));
  INV_X1    g455(.A(new_n403), .ZN(new_n642));
  AND4_X1   g456(.A1(new_n626), .A2(new_n640), .A3(new_n641), .A4(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n625), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT34), .B(G104), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  AND3_X1   g460(.A1(new_n335), .A2(new_n339), .A3(new_n325), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n325), .B1(new_n339), .B2(new_n346), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n351), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(KEYINPUT20), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n352), .ZN(new_n651));
  INV_X1    g465(.A(new_n342), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n651), .B(new_n652), .C1(new_n395), .C2(new_n410), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n403), .B(KEYINPUT91), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g469(.A(KEYINPUT92), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n362), .B1(new_n627), .B2(new_n628), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n409), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n342), .B1(new_n650), .B2(new_n352), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT92), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n658), .A2(new_n659), .A3(new_n660), .A4(new_n654), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n656), .A2(new_n626), .A3(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT93), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n656), .A2(KEYINPUT93), .A3(new_n661), .A4(new_n626), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n625), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT35), .B(G107), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G9));
  INV_X1    g483(.A(KEYINPUT36), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n556), .A2(new_n670), .A3(new_n559), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n672), .B1(new_n587), .B2(new_n592), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n596), .B(new_n671), .C1(new_n586), .C2(new_n576), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n673), .A2(new_n605), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(KEYINPUT94), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT94), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n673), .A2(new_n677), .A3(new_n674), .A4(new_n605), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n679), .A2(KEYINPUT95), .A3(new_n603), .ZN(new_n680));
  AOI21_X1  g494(.A(KEYINPUT95), .B1(new_n679), .B2(new_n603), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT96), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT95), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n676), .A2(new_n678), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n679), .A2(KEYINPUT95), .A3(new_n603), .ZN(new_n688));
  AOI21_X1  g502(.A(KEYINPUT96), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n623), .A2(new_n690), .A3(new_n467), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT37), .B(G110), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G12));
  INV_X1    g507(.A(new_n653), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n398), .B1(G900), .B2(new_n400), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n682), .B1(new_n680), .B2(new_n681), .ZN(new_n698));
  INV_X1    g512(.A(new_n413), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n438), .A2(KEYINPUT83), .A3(new_n417), .ZN(new_n700));
  AOI21_X1  g514(.A(KEYINPUT83), .B1(new_n438), .B2(new_n417), .ZN(new_n701));
  AOI21_X1  g515(.A(KEYINPUT12), .B1(new_n446), .B2(new_n435), .ZN(new_n702));
  AOI211_X1 g516(.A(new_n448), .B(new_n437), .C1(new_n445), .C2(new_n422), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n700), .A2(new_n701), .A3(new_n704), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n462), .B(new_n286), .C1(new_n705), .C2(new_n439), .ZN(new_n706));
  AOI22_X1  g520(.A1(new_n457), .A2(new_n416), .B1(new_n459), .B2(new_n436), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n463), .B1(new_n707), .B2(G469), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n699), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n687), .A2(KEYINPUT96), .A3(new_n688), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n698), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n626), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n616), .A2(new_n697), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G128), .ZN(G30));
  AOI21_X1  g529(.A(new_n473), .B1(new_n536), .B2(new_n490), .ZN(new_n716));
  OR2_X1    g530(.A1(new_n716), .A2(KEYINPUT97), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(KEYINPUT97), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n717), .A2(new_n517), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(G472), .B1(new_n719), .B2(G902), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n527), .B(new_n720), .C1(new_n614), .C2(new_n615), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n721), .A2(KEYINPUT98), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(KEYINPUT98), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n695), .B(KEYINPUT39), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n709), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(KEYINPUT99), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT40), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n292), .B(KEYINPUT38), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n687), .A2(new_n688), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n395), .A2(new_n410), .ZN(new_n731));
  NOR4_X1   g545(.A1(new_n730), .A2(new_n359), .A3(new_n357), .A4(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n724), .A2(new_n728), .A3(new_n729), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G143), .ZN(G45));
  NAND2_X1  g548(.A1(new_n355), .A2(new_n356), .ZN(new_n735));
  AOI22_X1  g549(.A1(new_n635), .A2(new_n639), .B1(new_n735), .B2(new_n652), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n695), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n553), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n713), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G146), .ZN(G48));
  OAI21_X1  g554(.A(G469), .B1(new_n454), .B2(G902), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(KEYINPUT100), .A3(new_n706), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT100), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n743), .B(G469), .C1(new_n454), .C2(G902), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n699), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n643), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n616), .A3(new_n618), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT101), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT101), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n746), .A2(new_n616), .A3(new_n749), .A4(new_n618), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(KEYINPUT41), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G113), .ZN(G15));
  NAND4_X1  g567(.A1(new_n666), .A2(new_n616), .A3(new_n618), .A4(new_n745), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G116), .ZN(G18));
  AND4_X1   g569(.A1(new_n357), .A2(new_n698), .A3(new_n411), .A4(new_n710), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n745), .A2(KEYINPUT102), .A3(new_n626), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT102), .B1(new_n745), .B2(new_n626), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n616), .B(new_n756), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G119), .ZN(G21));
  NAND2_X1  g574(.A1(new_n622), .A2(G472), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n473), .B1(new_n538), .B2(new_n539), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n523), .A2(new_n521), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n526), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AND4_X1   g578(.A1(new_n603), .A2(new_n761), .A3(new_n606), .A4(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n745), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n655), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n357), .A2(new_n359), .A3(new_n731), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n292), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT103), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n768), .A2(KEYINPUT103), .A3(new_n292), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n765), .A2(new_n767), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G122), .ZN(G24));
  INV_X1    g589(.A(new_n737), .ZN(new_n776));
  AOI21_X1  g590(.A(G902), .B1(new_n546), .B2(new_n519), .ZN(new_n777));
  INV_X1    g591(.A(G472), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n764), .B(new_n730), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n776), .B(new_n780), .C1(new_n757), .C2(new_n758), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G125), .ZN(G27));
  OR2_X1    g596(.A1(new_n547), .A2(KEYINPUT32), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n607), .B1(new_n783), .B2(new_n613), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n289), .A2(new_n290), .A3(new_n187), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n187), .B1(new_n289), .B2(new_n290), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n785), .A2(new_n786), .A3(new_n359), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n736), .A2(new_n709), .A3(new_n695), .A4(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n784), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n624), .A2(new_n787), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(KEYINPUT42), .ZN(new_n792));
  AOI22_X1  g606(.A1(KEYINPUT42), .A2(new_n790), .B1(new_n738), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G131), .ZN(G33));
  NAND4_X1  g608(.A1(new_n616), .A2(new_n624), .A3(new_n697), .A4(new_n787), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G134), .ZN(G36));
  XNOR2_X1  g610(.A(new_n357), .B(KEYINPUT106), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(KEYINPUT43), .A3(new_n640), .ZN(new_n798));
  XNOR2_X1  g612(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n799));
  INV_X1    g613(.A(new_n640), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n799), .B1(new_n800), .B2(new_n641), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n761), .A2(new_n550), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n803), .A2(KEYINPUT107), .A3(new_n730), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT107), .B1(new_n803), .B2(new_n730), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n802), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT44), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n288), .A2(new_n360), .A3(new_n291), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n707), .A2(KEYINPUT45), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n707), .A2(KEYINPUT45), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(G469), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT104), .ZN(new_n814));
  OR2_X1    g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n813), .A2(new_n814), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n463), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n817), .A2(KEYINPUT46), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n706), .B1(new_n817), .B2(KEYINPUT46), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n413), .B(new_n725), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n809), .A2(new_n810), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n821), .B1(new_n808), .B2(new_n807), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(G137), .ZN(G39));
  OAI21_X1  g637(.A(new_n413), .B1(new_n818), .B2(new_n819), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(KEYINPUT47), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT47), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n826), .B(new_n413), .C1(new_n818), .C2(new_n819), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n553), .A2(new_n611), .A3(new_n776), .A4(new_n787), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n825), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT108), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT108), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n825), .A2(new_n832), .A3(new_n827), .A4(new_n829), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(G140), .ZN(G42));
  NOR2_X1   g649(.A1(G952), .A2(G953), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT119), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n754), .A2(new_n759), .A3(new_n774), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n838), .A2(new_n751), .A3(new_n793), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n360), .B(new_n654), .C1(new_n785), .C2(new_n786), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n800), .A2(new_n357), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n625), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n357), .A2(new_n658), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n841), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n624), .A2(new_n550), .A3(new_n761), .A4(new_n845), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n691), .A2(KEYINPUT110), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT110), .B1(new_n691), .B2(new_n846), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n843), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n620), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n779), .A2(new_n788), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n711), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT111), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n731), .A2(new_n659), .A3(new_n695), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n810), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n731), .A2(new_n659), .A3(KEYINPUT111), .A4(new_n695), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT112), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n657), .A2(new_n409), .A3(new_n695), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n651), .A2(new_n652), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n854), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(new_n787), .A3(new_n857), .A4(KEYINPUT112), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n853), .B1(new_n858), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n852), .B1(new_n864), .B2(new_n553), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n553), .A2(new_n696), .A3(new_n791), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT113), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n861), .A2(new_n787), .A3(new_n857), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT112), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n711), .B1(new_n870), .B2(new_n862), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n851), .B1(new_n871), .B2(new_n616), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT113), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n872), .A2(new_n795), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n839), .A2(new_n840), .A3(new_n850), .A4(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n620), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n691), .A2(new_n846), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT110), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n691), .A2(new_n846), .A3(KEYINPUT110), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n880), .A2(new_n881), .B1(new_n625), .B2(new_n842), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n872), .A2(new_n873), .A3(new_n795), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n873), .B1(new_n872), .B2(new_n795), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n877), .B(new_n882), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n838), .A2(new_n751), .A3(new_n793), .ZN(new_n886));
  OAI21_X1  g700(.A(KEYINPUT114), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n616), .B(new_n713), .C1(new_n697), .C2(new_n776), .ZN(new_n888));
  AND4_X1   g702(.A1(new_n603), .A2(new_n709), .A3(new_n679), .A4(new_n695), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n721), .A2(new_n773), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n888), .A2(new_n781), .A3(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT52), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n888), .A2(new_n781), .A3(new_n890), .A4(KEYINPUT52), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n876), .A2(new_n887), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT53), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n895), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n754), .A2(new_n759), .A3(new_n774), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n750), .B2(new_n748), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n901), .A2(new_n875), .A3(new_n793), .A4(new_n850), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n899), .B1(new_n902), .B2(KEYINPUT114), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT53), .B1(new_n903), .B2(new_n876), .ZN(new_n904));
  OAI21_X1  g718(.A(KEYINPUT54), .B1(new_n898), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n896), .A2(new_n897), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n886), .A2(KEYINPUT115), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT115), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n838), .A2(new_n751), .A3(new_n908), .A4(new_n793), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n895), .A2(KEYINPUT53), .A3(new_n850), .A4(new_n875), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n906), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n905), .B1(KEYINPUT54), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n766), .A2(new_n810), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n916), .A2(new_n618), .A3(new_n399), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n724), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(new_n357), .A3(new_n800), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n398), .B1(new_n798), .B2(new_n801), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n920), .A2(new_n780), .A3(new_n916), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT117), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n920), .A2(new_n765), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n766), .A2(new_n729), .A3(new_n360), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT50), .Z(new_n927));
  AND2_X1   g741(.A1(new_n924), .A2(new_n787), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT116), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n742), .A2(new_n744), .ZN(new_n930));
  AOI22_X1  g744(.A1(new_n825), .A2(new_n827), .B1(new_n699), .B2(new_n930), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n923), .A2(KEYINPUT51), .A3(new_n927), .A4(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n920), .A2(new_n784), .A3(new_n916), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT48), .ZN(new_n935));
  OR3_X1    g749(.A1(new_n934), .A2(KEYINPUT118), .A3(new_n935), .ZN(new_n936));
  XNOR2_X1  g750(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n924), .B1(new_n758), .B2(new_n757), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n936), .A2(new_n396), .A3(new_n938), .A4(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n736), .B2(new_n918), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n932), .A2(new_n927), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n942), .A2(new_n922), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n933), .B(new_n941), .C1(new_n943), .C2(KEYINPUT51), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n837), .B1(new_n915), .B2(new_n944), .ZN(new_n945));
  NOR4_X1   g759(.A1(new_n800), .A2(new_n607), .A3(new_n699), .A4(new_n359), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT49), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n946), .B(new_n797), .C1(new_n947), .C2(new_n930), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT109), .Z(new_n949));
  AOI21_X1  g763(.A(new_n729), .B1(new_n947), .B2(new_n930), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n945), .B1(new_n724), .B2(new_n951), .ZN(G75));
  NOR2_X1   g766(.A1(new_n242), .A2(G952), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT120), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT56), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n914), .A2(G902), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n956), .B1(new_n957), .B2(new_n469), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n241), .A2(new_n275), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(new_n273), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT55), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n961), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n956), .B(new_n963), .C1(new_n957), .C2(new_n469), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n955), .B1(new_n962), .B2(new_n964), .ZN(G51));
  XNOR2_X1  g779(.A(new_n463), .B(KEYINPUT57), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n914), .A2(KEYINPUT54), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n912), .B1(new_n896), .B2(new_n897), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT54), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n966), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n440), .A2(new_n441), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n972), .A2(new_n453), .A3(new_n456), .ZN(new_n973));
  INV_X1    g787(.A(new_n439), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n914), .A2(G902), .A3(new_n816), .A4(new_n815), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n953), .B1(new_n976), .B2(new_n977), .ZN(G54));
  NAND2_X1  g792(.A1(KEYINPUT58), .A2(G475), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n957), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n980), .A2(new_n349), .ZN(new_n981));
  INV_X1    g795(.A(new_n349), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n957), .A2(new_n982), .A3(new_n979), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n981), .A2(new_n953), .A3(new_n983), .ZN(G60));
  INV_X1    g798(.A(new_n633), .ZN(new_n985));
  NAND2_X1  g799(.A1(G478), .A2(G902), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT59), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n985), .B(new_n987), .C1(new_n967), .C2(new_n970), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n954), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n985), .B1(new_n915), .B2(new_n987), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n989), .A2(new_n990), .ZN(G63));
  AND2_X1   g805(.A1(new_n673), .A2(new_n674), .ZN(new_n992));
  NAND2_X1  g806(.A1(G217), .A2(G902), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT60), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n992), .B(new_n995), .C1(new_n904), .C2(new_n912), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(KEYINPUT122), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT122), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n914), .A2(new_n998), .A3(new_n992), .A4(new_n995), .ZN(new_n999));
  INV_X1    g813(.A(new_n604), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n1000), .B1(new_n968), .B2(new_n994), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n997), .A2(new_n954), .A3(new_n999), .A4(new_n1001), .ZN(new_n1002));
  XOR2_X1   g816(.A(KEYINPUT121), .B(KEYINPUT61), .Z(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n1001), .A2(new_n996), .A3(KEYINPUT61), .A4(new_n954), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(G66));
  NAND2_X1  g820(.A1(new_n901), .A2(new_n850), .ZN(new_n1007));
  NAND2_X1  g821(.A1(G224), .A2(G953), .ZN(new_n1008));
  OAI22_X1  g822(.A1(new_n1007), .A2(G953), .B1(new_n402), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n959), .B1(G898), .B2(new_n242), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1009), .B(new_n1010), .Z(G69));
  NAND2_X1  g825(.A1(new_n514), .A2(new_n515), .ZN(new_n1012));
  OR2_X1    g826(.A1(new_n343), .A2(new_n344), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n784), .A2(new_n773), .ZN(new_n1016));
  OR2_X1    g830(.A1(new_n820), .A2(new_n1016), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n888), .A2(new_n781), .ZN(new_n1018));
  AND4_X1   g832(.A1(new_n793), .A2(new_n1017), .A3(new_n795), .A4(new_n1018), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n834), .A2(new_n1019), .A3(new_n822), .ZN(new_n1020));
  AND2_X1   g834(.A1(new_n1020), .A2(new_n242), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n242), .A2(G900), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1015), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n242), .B1(G227), .B2(G900), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1024), .B(KEYINPUT125), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n733), .A2(new_n1018), .ZN(new_n1026));
  OR2_X1    g840(.A1(new_n1026), .A2(KEYINPUT62), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n612), .A2(new_n619), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n844), .B1(new_n800), .B2(new_n357), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n1028), .A2(new_n727), .A3(new_n787), .A4(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n1030), .B(KEYINPUT124), .ZN(new_n1031));
  AND4_X1   g845(.A1(new_n822), .A2(new_n1027), .A3(new_n834), .A4(new_n1031), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1026), .A2(KEYINPUT62), .ZN(new_n1033));
  XNOR2_X1  g847(.A(new_n1033), .B(KEYINPUT123), .ZN(new_n1034));
  AOI21_X1  g848(.A(G953), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g849(.A(new_n1023), .B(new_n1025), .C1(new_n1035), .C2(new_n1015), .ZN(new_n1036));
  INV_X1    g850(.A(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1038), .A2(new_n242), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1039), .A2(new_n1014), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1025), .B1(new_n1040), .B2(new_n1023), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n1037), .A2(new_n1041), .ZN(G72));
  INV_X1    g856(.A(new_n529), .ZN(new_n1043));
  INV_X1    g857(.A(new_n1007), .ZN(new_n1044));
  NAND4_X1  g858(.A1(new_n834), .A2(new_n1019), .A3(new_n822), .A4(new_n1044), .ZN(new_n1045));
  NAND2_X1  g859(.A1(G472), .A2(G902), .ZN(new_n1046));
  XOR2_X1   g860(.A(new_n1046), .B(KEYINPUT63), .Z(new_n1047));
  AOI21_X1  g861(.A(new_n1043), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g862(.A(KEYINPUT126), .ZN(new_n1049));
  OR3_X1    g863(.A1(new_n1048), .A2(new_n1049), .A3(new_n953), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1049), .B1(new_n1048), .B2(new_n953), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n1047), .B1(new_n1038), .B2(new_n1007), .ZN(new_n1053));
  NAND3_X1  g867(.A1(new_n1053), .A2(new_n473), .A3(new_n528), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n528), .A2(new_n473), .ZN(new_n1055));
  NAND3_X1  g869(.A1(new_n1043), .A2(new_n1047), .A3(new_n1055), .ZN(new_n1056));
  XOR2_X1   g870(.A(new_n1056), .B(KEYINPUT127), .Z(new_n1057));
  OAI21_X1  g871(.A(new_n1057), .B1(new_n898), .B2(new_n904), .ZN(new_n1058));
  AND3_X1   g872(.A1(new_n1052), .A2(new_n1054), .A3(new_n1058), .ZN(G57));
endmodule


