//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1199, new_n1200, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT65), .Z(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n207), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n210), .B1(new_n214), .B2(new_n216), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  NAND2_X1  g0044(.A1(G33), .A2(G41), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n245), .A2(G1), .A3(G13), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT3), .B(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n247), .A2(G222), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(G1698), .ZN(new_n250));
  INV_X1    g0050(.A(G223), .ZN(new_n251));
  OAI221_X1 g0051(.A(new_n249), .B1(new_n203), .B2(new_n247), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n246), .B1(new_n252), .B2(KEYINPUT66), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n253), .B1(KEYINPUT66), .B2(new_n252), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n246), .A2(G274), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n246), .A2(new_n257), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n258), .B1(G226), .B2(new_n260), .ZN(new_n261));
  AND2_X1   g0061(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G190), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT71), .B(G200), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n264), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(KEYINPUT10), .B1(new_n266), .B2(KEYINPUT73), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n256), .A2(G13), .A3(G20), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT67), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n256), .A2(KEYINPUT67), .A3(G13), .A4(G20), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n211), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n256), .A2(G20), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(G50), .A3(new_n276), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT8), .B(G58), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n212), .A2(G33), .ZN(new_n279));
  INV_X1    g0079(.A(G150), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G20), .A2(G33), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI22_X1  g0082(.A1(new_n278), .A2(new_n279), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n212), .B1(new_n201), .B2(new_n202), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n274), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n270), .A2(new_n271), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n277), .B(new_n285), .C1(G50), .C2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n289), .B(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n266), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n267), .A2(new_n292), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n266), .B(new_n291), .C1(KEYINPUT73), .C2(KEYINPUT10), .ZN(new_n294));
  INV_X1    g0094(.A(G179), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n262), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n287), .B1(new_n262), .B2(G169), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n293), .A2(new_n294), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n257), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n300), .A2(new_n246), .A3(G274), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n301), .B1(new_n219), .B2(new_n259), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G33), .A2(G97), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n230), .A2(G1698), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(G226), .B2(G1698), .ZN(new_n305));
  AND2_X1   g0105(.A1(KEYINPUT3), .A2(G33), .ZN(new_n306));
  NOR2_X1   g0106(.A1(KEYINPUT3), .A2(G33), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n303), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  OR2_X1    g0109(.A1(new_n309), .A2(KEYINPUT74), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n246), .B1(new_n309), .B2(KEYINPUT74), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n302), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT13), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n313), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G169), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT14), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT14), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n316), .A2(new_n319), .A3(G169), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n318), .B(new_n320), .C1(new_n295), .C2(new_n316), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n272), .A2(new_n218), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT12), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n275), .A2(G68), .A3(new_n276), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n323), .A2(KEYINPUT75), .A3(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n282), .A2(new_n202), .ZN(new_n326));
  OAI22_X1  g0126(.A1(new_n279), .A2(new_n203), .B1(new_n212), .B2(G68), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n274), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n328), .B(KEYINPUT11), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(KEYINPUT75), .B1(new_n323), .B2(new_n324), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n321), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n316), .A2(G200), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n314), .A2(G190), .A3(new_n315), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n332), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n247), .A2(G232), .A3(new_n248), .ZN(new_n339));
  INV_X1    g0139(.A(G107), .ZN(new_n340));
  OAI221_X1 g0140(.A(new_n339), .B1(new_n340), .B2(new_n247), .C1(new_n250), .C2(new_n219), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n258), .B1(G244), .B2(new_n260), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT68), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n343), .A2(KEYINPUT68), .A3(new_n344), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OR2_X1    g0149(.A1(new_n349), .A2(new_n263), .ZN(new_n350));
  INV_X1    g0150(.A(new_n274), .ZN(new_n351));
  XOR2_X1   g0151(.A(new_n278), .B(KEYINPUT69), .Z(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n281), .B(KEYINPUT70), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT15), .B(G87), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n279), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n357), .A2(new_n358), .B1(G20), .B2(G77), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n351), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n203), .B1(new_n256), .B2(G20), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n275), .A2(new_n361), .B1(new_n203), .B2(new_n272), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n350), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n349), .A2(new_n265), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n364), .ZN(new_n368));
  INV_X1    g0168(.A(G169), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n347), .A2(new_n369), .A3(new_n348), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n368), .B(new_n370), .C1(new_n349), .C2(G179), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n251), .A2(new_n248), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n247), .B(new_n373), .C1(G226), .C2(new_n248), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G33), .A2(G87), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n246), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n301), .B1(new_n230), .B2(new_n259), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(G169), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n295), .B2(new_n378), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT7), .B1(new_n308), .B2(new_n212), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT3), .ZN(new_n382));
  INV_X1    g0182(.A(G33), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(KEYINPUT3), .A2(G33), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n384), .A2(KEYINPUT7), .A3(new_n212), .A4(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(G68), .B1(new_n381), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g0188(.A(G58), .B(G68), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n389), .A2(G20), .B1(G159), .B2(new_n281), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT16), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n388), .A2(KEYINPUT16), .A3(new_n390), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(new_n394), .A3(new_n274), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n278), .B1(new_n256), .B2(G20), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n275), .A2(new_n396), .B1(new_n272), .B2(new_n278), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT18), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n380), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n399), .B1(new_n380), .B2(new_n398), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT76), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n380), .A2(new_n398), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT18), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT76), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n380), .A2(new_n398), .A3(new_n399), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G200), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n374), .A2(new_n375), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n342), .ZN(new_n411));
  INV_X1    g0211(.A(new_n377), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n376), .A2(new_n377), .A3(new_n263), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n415), .A2(new_n395), .A3(new_n397), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT78), .ZN(new_n417));
  XOR2_X1   g0217(.A(KEYINPUT77), .B(KEYINPUT17), .Z(new_n418));
  NAND3_X1  g0218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n415), .A2(new_n395), .A3(new_n397), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n420), .A2(KEYINPUT17), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n415), .A2(new_n395), .A3(new_n397), .A4(new_n418), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT78), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n419), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n408), .A2(new_n425), .ZN(new_n426));
  NOR4_X1   g0226(.A1(new_n299), .A2(new_n338), .A3(new_n372), .A4(new_n426), .ZN(new_n427));
  XOR2_X1   g0227(.A(KEYINPUT85), .B(KEYINPUT25), .Z(new_n428));
  NAND3_X1  g0228(.A1(new_n272), .A2(new_n340), .A3(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(KEYINPUT85), .B(KEYINPUT25), .C1(new_n286), .C2(G107), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT79), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n256), .B2(G33), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n383), .A2(KEYINPUT79), .A3(G1), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n286), .A2(new_n435), .A3(new_n351), .ZN(new_n436));
  OR2_X1    g0236(.A1(new_n436), .A2(new_n340), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n431), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n247), .A2(new_n212), .A3(G87), .ZN(new_n439));
  AND2_X1   g0239(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n440));
  NOR2_X1   g0240(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n247), .A2(new_n212), .A3(G87), .A4(new_n440), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT23), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n445), .B1(new_n212), .B2(G107), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n340), .A2(KEYINPUT23), .A3(G20), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n358), .A2(G116), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n443), .A2(new_n444), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT24), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n449), .A2(KEYINPUT84), .A3(new_n450), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n451), .A2(new_n274), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n449), .A2(KEYINPUT84), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT84), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n443), .A2(new_n454), .A3(new_n444), .A4(new_n448), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(KEYINPUT24), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n438), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(G250), .B(new_n248), .C1(new_n306), .C2(new_n307), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT86), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT86), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n247), .A2(new_n461), .A3(G250), .A4(new_n248), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G294), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n247), .A2(G257), .A3(G1698), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n460), .A2(new_n462), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n342), .ZN(new_n466));
  INV_X1    g0266(.A(G45), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(G1), .ZN(new_n468));
  AND2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  NOR2_X1   g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AND3_X1   g0271(.A1(new_n471), .A2(G264), .A3(new_n246), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT88), .B1(new_n466), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT88), .ZN(new_n475));
  AOI211_X1 g0275(.A(new_n475), .B(new_n472), .C1(new_n465), .C2(new_n342), .ZN(new_n476));
  XNOR2_X1  g0276(.A(KEYINPUT5), .B(G41), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n477), .A2(G274), .A3(new_n246), .A4(new_n468), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NOR4_X1   g0279(.A1(new_n474), .A2(new_n476), .A3(new_n295), .A4(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT87), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n466), .A2(new_n473), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(new_n479), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n472), .B1(new_n465), .B2(new_n342), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(KEYINPUT87), .A3(new_n478), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n369), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n458), .B1(new_n480), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n474), .A2(new_n476), .ZN(new_n488));
  AOI21_X1  g0288(.A(G200), .B1(new_n488), .B2(new_n478), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n484), .A2(KEYINPUT87), .A3(new_n478), .ZN(new_n490));
  AOI21_X1  g0290(.A(KEYINPUT87), .B1(new_n484), .B2(new_n478), .ZN(new_n491));
  NOR3_X1   g0291(.A1(new_n490), .A2(new_n491), .A3(G190), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n457), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G283), .ZN(new_n495));
  INV_X1    g0295(.A(G97), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n495), .B(new_n212), .C1(G33), .C2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(G116), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G20), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n274), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT20), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT82), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n274), .A2(new_n499), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT82), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n503), .A2(new_n504), .A3(new_n497), .A4(KEYINPUT20), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n500), .A2(new_n501), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n502), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(G116), .B1(new_n270), .B2(new_n271), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n508), .B1(new_n436), .B2(G116), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT81), .ZN(new_n511));
  OAI211_X1 g0311(.A(G264), .B(G1698), .C1(new_n306), .C2(new_n307), .ZN(new_n512));
  OAI211_X1 g0312(.A(G257), .B(new_n248), .C1(new_n306), .C2(new_n307), .ZN(new_n513));
  INV_X1    g0313(.A(G303), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n512), .B(new_n513), .C1(new_n514), .C2(new_n247), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n515), .A2(new_n342), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n471), .A2(new_n246), .ZN(new_n517));
  INV_X1    g0317(.A(G270), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n478), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n511), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n519), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n515), .A2(new_n342), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(KEYINPUT81), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n510), .B1(new_n525), .B2(new_n263), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n526), .B1(G200), .B2(new_n525), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT21), .ZN(new_n528));
  OAI21_X1  g0328(.A(G169), .B1(new_n507), .B2(new_n509), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n528), .B1(new_n524), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n509), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n502), .A2(new_n505), .A3(new_n506), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n369), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n533), .A2(KEYINPUT21), .A3(new_n520), .A4(new_n523), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n521), .A2(G179), .A3(new_n522), .ZN(new_n535));
  OR2_X1    g0335(.A1(new_n510), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n530), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n527), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n471), .A2(G257), .A3(new_n246), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n478), .ZN(new_n540));
  OAI211_X1 g0340(.A(G244), .B(new_n248), .C1(new_n306), .C2(new_n307), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT4), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n247), .A2(KEYINPUT4), .A3(G244), .A4(new_n248), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n247), .A2(G250), .A3(G1698), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n495), .A4(new_n545), .ZN(new_n546));
  AOI211_X1 g0346(.A(new_n263), .B(new_n540), .C1(new_n546), .C2(new_n342), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n282), .A2(new_n203), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n340), .A2(KEYINPUT6), .A3(G97), .ZN(new_n550));
  XNOR2_X1  g0350(.A(G97), .B(G107), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT6), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n549), .B1(new_n553), .B2(new_n212), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n384), .A2(new_n212), .A3(new_n385), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT7), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n340), .B1(new_n557), .B2(new_n386), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n274), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n272), .A2(new_n496), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n286), .A2(new_n435), .A3(new_n351), .A4(G97), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n547), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n546), .A2(new_n342), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT80), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n546), .A2(KEYINPUT80), .A3(new_n342), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n540), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n564), .B1(new_n569), .B2(new_n409), .ZN(new_n570));
  INV_X1    g0370(.A(new_n540), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n572), .A2(new_n369), .B1(new_n559), .B2(new_n562), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n546), .A2(KEYINPUT80), .A3(new_n342), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT80), .B1(new_n546), .B2(new_n342), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n295), .B(new_n571), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(G238), .B(new_n248), .C1(new_n306), .C2(new_n307), .ZN(new_n578));
  OAI211_X1 g0378(.A(G244), .B(G1698), .C1(new_n306), .C2(new_n307), .ZN(new_n579));
  NAND2_X1  g0379(.A1(G33), .A2(G116), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n342), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n256), .A2(G45), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G250), .ZN(new_n584));
  OAI22_X1  g0384(.A1(new_n255), .A2(new_n583), .B1(new_n342), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n265), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT19), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n212), .B1(new_n303), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(G97), .A2(G107), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n220), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n212), .B(G68), .C1(new_n306), .C2(new_n307), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n589), .B1(new_n279), .B2(new_n496), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n274), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n272), .A2(new_n356), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n286), .A2(new_n435), .A3(new_n351), .A4(G87), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n582), .A2(new_n586), .A3(G190), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n588), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n582), .A2(new_n586), .A3(new_n295), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n286), .A2(new_n435), .A3(new_n351), .A4(new_n357), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n597), .A2(new_n598), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n585), .B1(new_n342), .B2(new_n581), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n603), .B(new_n605), .C1(G169), .C2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n570), .A2(new_n577), .A3(new_n609), .ZN(new_n610));
  AND4_X1   g0410(.A1(new_n427), .A2(new_n494), .A3(new_n538), .A4(new_n610), .ZN(G372));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n493), .ZN(new_n612));
  OAI21_X1  g0412(.A(G169), .B1(new_n490), .B2(new_n491), .ZN(new_n613));
  INV_X1    g0413(.A(new_n474), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n484), .A2(KEYINPUT88), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n614), .A2(G179), .A3(new_n478), .A4(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n457), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n617), .A2(new_n537), .ZN(new_n618));
  OR3_X1    g0418(.A1(new_n612), .A2(new_n618), .A3(KEYINPUT89), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n540), .B1(new_n546), .B2(new_n342), .ZN(new_n620));
  OAI21_X1  g0420(.A(G107), .B1(new_n381), .B2(new_n387), .ZN(new_n621));
  AND2_X1   g0421(.A1(G97), .A2(G107), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n552), .B1(new_n622), .B2(new_n591), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n340), .A2(KEYINPUT6), .A3(G97), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n548), .B1(new_n625), .B2(G20), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n351), .B1(new_n621), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n560), .A2(new_n561), .ZN(new_n628));
  OAI22_X1  g0428(.A1(new_n620), .A2(G169), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(new_n569), .B2(new_n295), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT26), .B1(new_n630), .B2(new_n609), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT26), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n577), .A2(new_n632), .A3(new_n608), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n607), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(KEYINPUT89), .B1(new_n612), .B2(new_n618), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n619), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n427), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n298), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n400), .A2(new_n401), .ZN(new_n641));
  INV_X1    g0441(.A(new_n371), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n321), .A2(new_n333), .B1(new_n337), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n641), .B1(new_n643), .B2(new_n424), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n293), .A2(new_n294), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n640), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n639), .A2(new_n646), .ZN(G369));
  NAND3_X1  g0447(.A1(new_n256), .A2(new_n212), .A3(G13), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n649));
  XOR2_X1   g0449(.A(new_n649), .B(KEYINPUT90), .Z(new_n650));
  INV_X1    g0450(.A(G213), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n653));
  XOR2_X1   g0453(.A(new_n653), .B(KEYINPUT91), .Z(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(new_n510), .ZN(new_n658));
  MUX2_X1   g0458(.A(new_n538), .B(new_n537), .S(new_n658), .Z(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(G330), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n494), .B1(new_n457), .B2(new_n657), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n487), .B2(new_n657), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n530), .A2(new_n534), .A3(new_n536), .ZN(new_n664));
  INV_X1    g0464(.A(new_n657), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n494), .A2(new_n666), .B1(new_n617), .B2(new_n657), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n663), .A2(new_n667), .ZN(G399));
  INV_X1    g0468(.A(new_n208), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT92), .B1(new_n669), .B2(G41), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n669), .A2(KEYINPUT92), .A3(G41), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n591), .A2(new_n220), .A3(new_n498), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n673), .A2(new_n256), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n216), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(new_n673), .ZN(new_n677));
  XOR2_X1   g0477(.A(new_n677), .B(KEYINPUT28), .Z(new_n678));
  INV_X1    g0478(.A(G330), .ZN(new_n679));
  XNOR2_X1  g0479(.A(KEYINPUT93), .B(KEYINPUT31), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n657), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n572), .A2(new_n535), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n614), .A2(new_n615), .A3(new_n606), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(KEYINPUT94), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n683), .A2(KEYINPUT94), .ZN(new_n686));
  OAI211_X1 g0486(.A(KEYINPUT30), .B(new_n682), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n569), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n525), .A2(new_n295), .A3(new_n688), .A4(new_n587), .ZN(new_n689));
  NOR3_X1   g0489(.A1(new_n474), .A2(new_n476), .A3(new_n479), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n682), .B1(new_n685), .B2(new_n686), .ZN(new_n692));
  XOR2_X1   g0492(.A(KEYINPUT95), .B(KEYINPUT30), .Z(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n691), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT96), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n687), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n689), .A2(new_n690), .ZN(new_n698));
  INV_X1    g0498(.A(new_n682), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n683), .A2(KEYINPUT94), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n699), .B1(new_n700), .B2(new_n684), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n698), .B1(new_n701), .B2(new_n693), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(KEYINPUT96), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n681), .B1(new_n697), .B2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n538), .A2(new_n494), .A3(new_n610), .A4(new_n657), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT31), .ZN(new_n706));
  INV_X1    g0506(.A(new_n687), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n665), .B1(new_n702), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n679), .B1(new_n704), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(KEYINPUT98), .B1(new_n612), .B2(new_n618), .ZN(new_n711));
  OAI211_X1 g0511(.A(KEYINPUT97), .B(new_n632), .C1(new_n577), .C2(new_n608), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n607), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT97), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n713), .B1(new_n634), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n487), .A2(new_n664), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT98), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n716), .A2(new_n717), .A3(new_n493), .A4(new_n610), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n711), .A2(new_n715), .A3(new_n718), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n719), .A2(KEYINPUT99), .A3(new_n657), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT99), .B1(new_n719), .B2(new_n657), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT29), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n638), .A2(new_n657), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT29), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n710), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n678), .B1(new_n726), .B2(G1), .ZN(G364));
  NAND2_X1  g0527(.A1(new_n212), .A2(G13), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n256), .B1(new_n729), .B2(G45), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n673), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n660), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(G330), .B2(new_n659), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n669), .A2(new_n308), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G355), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(G116), .B2(new_n208), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n240), .A2(new_n467), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n669), .A2(new_n247), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n740), .B1(new_n467), .B2(new_n676), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n737), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G13), .A2(G33), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n211), .B1(G20), .B2(new_n369), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n732), .B1(new_n742), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n212), .A2(new_n263), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n295), .A2(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n212), .A2(G190), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G179), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI22_X1  g0557(.A1(G322), .A2(new_n753), .B1(new_n757), .B2(G329), .ZN(new_n758));
  INV_X1    g0558(.A(G311), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n754), .A2(new_n751), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n758), .B(new_n308), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n755), .A2(G190), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n761), .B1(G294), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n265), .A2(new_n295), .A3(new_n754), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n265), .A2(new_n295), .A3(new_n750), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(G283), .A2(new_n766), .B1(new_n768), .B2(G303), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n212), .A2(new_n295), .A3(new_n409), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n770), .A2(KEYINPUT101), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(KEYINPUT101), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n263), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n771), .A2(new_n263), .A3(new_n772), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(KEYINPUT33), .B(G317), .ZN(new_n777));
  AOI22_X1  g0577(.A1(G326), .A2(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n764), .A2(new_n769), .A3(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G159), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n756), .A2(new_n780), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT32), .Z(new_n782));
  AOI211_X1 g0582(.A(new_n308), .B(new_n782), .C1(G97), .C2(new_n763), .ZN(new_n783));
  INV_X1    g0583(.A(new_n774), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n783), .B1(new_n218), .B2(new_n775), .C1(new_n202), .C2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G58), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n752), .A2(new_n786), .B1(new_n760), .B2(new_n203), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT100), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n768), .A2(G87), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n788), .B(new_n789), .C1(new_n340), .C2(new_n765), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n779), .B1(new_n785), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT102), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n746), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(new_n791), .B2(new_n792), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n749), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n745), .B(KEYINPUT103), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n796), .B1(new_n659), .B2(new_n797), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n734), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(G396));
  INV_X1    g0600(.A(KEYINPUT104), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n665), .A2(new_n368), .ZN(new_n802));
  AND3_X1   g0602(.A1(new_n371), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n802), .B1(new_n371), .B2(new_n801), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n367), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n723), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n805), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n638), .A2(new_n807), .A3(new_n657), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n710), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n732), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n710), .A2(new_n806), .A3(new_n808), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n766), .A2(G68), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n308), .B1(new_n757), .B2(G132), .ZN(new_n814));
  INV_X1    g0614(.A(new_n763), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n813), .B(new_n814), .C1(new_n786), .C2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n760), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n753), .A2(G143), .B1(new_n817), .B2(G159), .ZN(new_n818));
  INV_X1    g0618(.A(G137), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n818), .B1(new_n280), .B2(new_n775), .C1(new_n784), .C2(new_n819), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT34), .Z(new_n821));
  AOI211_X1 g0621(.A(new_n816), .B(new_n821), .C1(G50), .C2(new_n768), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G303), .A2(new_n774), .B1(new_n776), .B2(G283), .ZN(new_n823));
  INV_X1    g0623(.A(G294), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n308), .B1(new_n752), .B2(new_n824), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n760), .A2(new_n498), .B1(new_n756), .B2(new_n759), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n825), .B(new_n826), .C1(G97), .C2(new_n763), .ZN(new_n827));
  AOI22_X1  g0627(.A1(G87), .A2(new_n766), .B1(new_n768), .B2(G107), .ZN(new_n828));
  AND3_X1   g0628(.A1(new_n823), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n746), .B1(new_n822), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n732), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n746), .A2(new_n743), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n831), .B1(new_n203), .B2(new_n832), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n830), .B(new_n833), .C1(new_n807), .C2(new_n744), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n812), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(G384));
  AND2_X1   g0636(.A1(new_n625), .A2(KEYINPUT35), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n625), .A2(KEYINPUT35), .ZN(new_n838));
  NOR4_X1   g0638(.A1(new_n837), .A2(new_n214), .A3(new_n838), .A4(new_n498), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT36), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n676), .B(G77), .C1(new_n786), .C2(new_n218), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n202), .A2(G68), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n256), .B(G13), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n371), .A2(new_n665), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n808), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n655), .B1(new_n395), .B2(new_n397), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n849), .A2(new_n403), .A3(new_n420), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n849), .A2(KEYINPUT105), .A3(new_n420), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT37), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n416), .A2(new_n848), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n854), .B(new_n403), .C1(KEYINPUT105), .C2(KEYINPUT37), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n424), .B1(new_n402), .B2(new_n407), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n856), .B(KEYINPUT38), .C1(new_n857), .C2(new_n849), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT106), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n426), .A2(new_n848), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n861), .A2(KEYINPUT106), .A3(KEYINPUT38), .A4(new_n856), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT38), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n849), .B1(new_n408), .B2(new_n425), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n853), .A2(new_n855), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n860), .A2(new_n862), .A3(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n334), .B(new_n337), .C1(new_n332), .C2(new_n657), .ZN(new_n868));
  INV_X1    g0668(.A(new_n337), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n333), .B(new_n665), .C1(new_n321), .C2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n847), .A2(new_n867), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n655), .B1(new_n400), .B2(new_n401), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n321), .A2(new_n333), .A3(new_n657), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n867), .A2(KEYINPUT39), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n849), .B1(new_n425), .B2(new_n641), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n863), .B1(new_n878), .B2(new_n865), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n879), .A2(new_n858), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT39), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n874), .B1(new_n876), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n722), .A2(new_n427), .A3(new_n725), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n646), .ZN(new_n886));
  XOR2_X1   g0686(.A(new_n884), .B(new_n886), .Z(new_n887));
  INV_X1    g0687(.A(new_n680), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n708), .A2(new_n705), .A3(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT31), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n890), .B(new_n665), .C1(new_n702), .C2(new_n707), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT40), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n805), .B1(new_n868), .B2(new_n870), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n867), .A2(new_n892), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(new_n891), .A3(new_n889), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT40), .B1(new_n896), .B2(new_n880), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n892), .A2(new_n427), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n679), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n899), .B2(new_n898), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n887), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n256), .B2(new_n729), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n887), .A2(new_n901), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n844), .B1(new_n903), .B2(new_n904), .ZN(G367));
  NAND2_X1  g0705(.A1(new_n236), .A2(new_n739), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n748), .B1(new_n669), .B2(new_n357), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n831), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n657), .A2(new_n600), .ZN(new_n909));
  MUX2_X1   g0709(.A(new_n609), .B(new_n635), .S(new_n909), .Z(new_n910));
  AOI22_X1  g0710(.A1(G143), .A2(new_n774), .B1(new_n776), .B2(G159), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n763), .A2(G68), .ZN(new_n912));
  OAI22_X1  g0712(.A1(new_n752), .A2(new_n280), .B1(new_n756), .B2(new_n819), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n308), .B(new_n913), .C1(G50), .C2(new_n817), .ZN(new_n914));
  AOI22_X1  g0714(.A1(G58), .A2(new_n768), .B1(new_n766), .B2(G77), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n911), .A2(new_n912), .A3(new_n914), .A4(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n767), .A2(new_n498), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n774), .A2(G311), .B1(KEYINPUT46), .B2(new_n917), .ZN(new_n918));
  OAI221_X1 g0718(.A(new_n918), .B1(KEYINPUT46), .B2(new_n917), .C1(new_n824), .C2(new_n775), .ZN(new_n919));
  INV_X1    g0719(.A(G283), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n308), .B1(new_n760), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(G317), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n752), .A2(new_n514), .B1(new_n756), .B2(new_n922), .ZN(new_n923));
  AOI211_X1 g0723(.A(new_n921), .B(new_n923), .C1(G107), .C2(new_n763), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n496), .B2(new_n765), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n916), .B1(new_n919), .B2(new_n925), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n926), .B(KEYINPUT47), .Z(new_n927));
  OAI221_X1 g0727(.A(new_n908), .B1(new_n910), .B2(new_n797), .C1(new_n927), .C2(new_n794), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n665), .A2(new_n563), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(new_n577), .A3(new_n570), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n665), .A2(new_n630), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n667), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT107), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n934), .A2(KEYINPUT44), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(KEYINPUT44), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n667), .A2(new_n932), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n937), .B(KEYINPUT45), .Z(new_n938));
  NAND3_X1  g0738(.A1(new_n935), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n663), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n939), .A2(KEYINPUT108), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(KEYINPUT108), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n935), .A2(new_n936), .A3(new_n942), .A4(new_n938), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n494), .A2(new_n666), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n662), .B2(new_n666), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(new_n660), .Z(new_n947));
  OAI21_X1  g0747(.A(new_n726), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n673), .B(KEYINPUT41), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n731), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n932), .A2(new_n494), .A3(new_n666), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n951), .A2(KEYINPUT42), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n577), .B1(new_n930), .B2(new_n487), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n951), .A2(KEYINPUT42), .B1(new_n657), .B2(new_n953), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n952), .A2(new_n954), .B1(KEYINPUT43), .B2(new_n910), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n910), .A2(KEYINPUT43), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n955), .B(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n940), .A2(new_n932), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n957), .B(new_n958), .Z(new_n959));
  OAI21_X1  g0759(.A(new_n928), .B1(new_n950), .B2(new_n959), .ZN(G387));
  INV_X1    g0760(.A(new_n673), .ZN(new_n961));
  INV_X1    g0761(.A(new_n947), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n961), .B1(new_n962), .B2(new_n726), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n726), .B2(new_n962), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n753), .A2(G317), .B1(new_n817), .B2(G303), .ZN(new_n965));
  INV_X1    g0765(.A(G322), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n965), .B1(new_n759), .B2(new_n775), .C1(new_n784), .C2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT48), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n768), .A2(G294), .B1(G283), .B2(new_n763), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT49), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(new_n973), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n765), .A2(new_n498), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n247), .B(new_n976), .C1(G326), .C2(new_n757), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n974), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n774), .A2(G159), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT109), .Z(new_n980));
  INV_X1    g0780(.A(new_n278), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n776), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n815), .A2(new_n356), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n247), .B1(new_n760), .B2(new_n218), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n752), .A2(new_n202), .B1(new_n756), .B2(new_n280), .ZN(new_n985));
  NOR3_X1   g0785(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  AOI22_X1  g0786(.A1(G77), .A2(new_n768), .B1(new_n766), .B2(G97), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n980), .A2(new_n982), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n794), .B1(new_n978), .B2(new_n988), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n735), .A2(new_n674), .B1(new_n340), .B2(new_n669), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n353), .A2(new_n202), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT50), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n467), .B1(new_n218), .B2(new_n203), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n992), .A2(new_n674), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n739), .B1(new_n233), .B2(new_n467), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n990), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n831), .B(new_n989), .C1(new_n747), .C2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT110), .Z(new_n998));
  OR2_X1    g0798(.A1(new_n662), .A2(new_n797), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n998), .A2(new_n999), .B1(new_n731), .B2(new_n962), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n964), .A2(new_n1000), .ZN(G393));
  XNOR2_X1  g0801(.A(new_n939), .B(new_n663), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n731), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n930), .A2(new_n745), .A3(new_n931), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT111), .Z(new_n1005));
  OAI221_X1 g0805(.A(new_n308), .B1(new_n756), .B2(new_n966), .C1(new_n824), .C2(new_n760), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(G116), .B2(new_n763), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(G107), .A2(new_n766), .B1(new_n768), .B2(G283), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1007), .B(new_n1008), .C1(new_n514), .C2(new_n775), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n774), .A2(G317), .B1(G311), .B2(new_n753), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT52), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n774), .A2(G150), .B1(G159), .B2(new_n753), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT51), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n353), .A2(new_n817), .B1(new_n768), .B2(G68), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n308), .B1(new_n757), .B2(G143), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n203), .B2(new_n815), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G87), .B2(new_n766), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1014), .B(new_n1017), .C1(new_n202), .C2(new_n775), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n1009), .A2(new_n1011), .B1(new_n1013), .B2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT112), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n746), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n747), .B1(new_n496), .B2(new_n208), .C1(new_n243), .C2(new_n740), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1005), .A2(new_n1021), .A3(new_n732), .A4(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1003), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n962), .A2(new_n726), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n944), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1026), .A2(new_n961), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1002), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n1025), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1024), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(G390));
  AOI21_X1  g0831(.A(new_n876), .B1(new_n847), .B2(new_n871), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n883), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n871), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n807), .B1(new_n720), .B2(new_n721), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1035), .B1(new_n1036), .B2(new_n846), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT113), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n880), .A2(new_n876), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  NOR3_X1   g0840(.A1(new_n1037), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n719), .A2(new_n657), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT99), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n719), .A2(KEYINPUT99), .A3(new_n657), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n805), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n871), .B1(new_n1046), .B2(new_n845), .ZN(new_n1047));
  AOI21_X1  g0847(.A(KEYINPUT113), .B1(new_n1047), .B2(new_n1039), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1034), .B1(new_n1041), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT114), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n894), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n889), .A2(new_n891), .ZN(new_n1052));
  NOR3_X1   g0852(.A1(new_n1051), .A2(new_n1052), .A3(new_n679), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1049), .A2(new_n1050), .A3(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1038), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n845), .B1(new_n1056), .B2(new_n807), .ZN(new_n1057));
  OAI211_X1 g0857(.A(KEYINPUT113), .B(new_n1039), .C1(new_n1057), .C2(new_n1035), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1033), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1053), .ZN(new_n1060));
  OAI21_X1  g0860(.A(KEYINPUT114), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n710), .A2(new_n807), .A3(new_n871), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1054), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n871), .B1(new_n710), .B2(new_n807), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n847), .B1(new_n1065), .B2(new_n1053), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n889), .A2(new_n807), .A3(G330), .A4(new_n891), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n1035), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1057), .A2(new_n1062), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n892), .A2(new_n427), .A3(G330), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n885), .A2(new_n646), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT115), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n885), .A2(new_n646), .A3(KEYINPUT115), .A4(new_n1071), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1070), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1064), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1076), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1054), .A2(new_n1061), .A3(new_n1063), .A4(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1077), .A2(new_n673), .A3(new_n1079), .ZN(new_n1080));
  AND3_X1   g0880(.A1(new_n1054), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n877), .A2(new_n743), .A3(new_n882), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n832), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n732), .B1(new_n981), .B2(new_n1083), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(KEYINPUT54), .B(G143), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n753), .A2(G132), .B1(new_n817), .B2(new_n1086), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1087), .B1(new_n780), .B2(new_n815), .C1(new_n775), .C2(new_n819), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(G128), .B2(new_n774), .ZN(new_n1089));
  INV_X1    g0889(.A(G125), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n247), .B1(new_n1090), .B2(new_n756), .C1(new_n765), .C2(new_n202), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT116), .Z(new_n1092));
  NOR2_X1   g0892(.A1(new_n767), .A2(new_n280), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT53), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1089), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT117), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G283), .A2(new_n774), .B1(new_n776), .B2(G107), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n308), .B1(new_n760), .B2(new_n496), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n752), .A2(new_n498), .B1(new_n756), .B2(new_n824), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1099), .B(new_n1100), .C1(G77), .C2(new_n763), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1098), .A2(new_n789), .A3(new_n813), .A4(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1097), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1084), .B1(new_n1104), .B2(new_n746), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1081), .A2(new_n731), .B1(new_n1082), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1080), .A2(new_n1106), .ZN(G378));
  NAND2_X1  g0907(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1079), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n898), .A2(G330), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n299), .A2(new_n287), .A3(new_n656), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n656), .A2(new_n287), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n293), .A2(new_n294), .A3(new_n298), .A4(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n1112), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1115), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1111), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1118), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n898), .A2(G330), .A3(new_n1120), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n1119), .A2(new_n884), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n884), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT57), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1110), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n673), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1124), .ZN(new_n1129));
  AOI21_X1  g0929(.A(KEYINPUT57), .B1(new_n1110), .B2(new_n1129), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1118), .A2(new_n743), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n732), .B1(G50), .B2(new_n1083), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n784), .A2(new_n498), .B1(new_n496), .B2(new_n775), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n247), .A2(G41), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n752), .A2(new_n340), .B1(new_n760), .B2(new_n356), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1135), .B(new_n1136), .C1(G283), .C2(new_n757), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n768), .A2(G77), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1137), .A2(new_n912), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n766), .A2(G58), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT118), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n1134), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1144));
  INV_X1    g0944(.A(G41), .ZN(new_n1145));
  AOI21_X1  g0945(.A(G50), .B1(new_n383), .B2(new_n1145), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1143), .A2(new_n1144), .B1(new_n1135), .B2(new_n1146), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n753), .A2(G128), .B1(new_n817), .B2(G137), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n280), .B2(new_n815), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n768), .B2(new_n1086), .ZN(new_n1150));
  INV_X1    g0950(.A(G132), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1150), .B1(new_n1090), .B2(new_n784), .C1(new_n1151), .C2(new_n775), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1152), .A2(KEYINPUT59), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(KEYINPUT59), .ZN(new_n1154));
  AOI211_X1 g0954(.A(G33), .B(G41), .C1(new_n757), .C2(G124), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n780), .B2(new_n765), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT120), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1147), .B1(new_n1144), .B2(new_n1143), .C1(new_n1153), .C2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1133), .B1(new_n1159), .B2(new_n746), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n1129), .A2(new_n731), .B1(new_n1132), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1131), .A2(new_n1161), .ZN(G375));
  INV_X1    g0962(.A(new_n1070), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1108), .A2(new_n1163), .A3(KEYINPUT122), .ZN(new_n1164));
  AOI21_X1  g0964(.A(KEYINPUT122), .B1(new_n1108), .B2(new_n1163), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n949), .B(KEYINPUT121), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1166), .A2(new_n1076), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1070), .A2(new_n731), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT123), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1169), .B(new_n1170), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n784), .A2(new_n824), .B1(new_n498), .B2(new_n775), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(G107), .A2(new_n817), .B1(new_n757), .B2(G303), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1173), .B(new_n308), .C1(new_n920), .C2(new_n752), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n203), .A2(new_n765), .B1(new_n767), .B2(new_n496), .ZN(new_n1175));
  NOR4_X1   g0975(.A1(new_n1172), .A2(new_n983), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n784), .A2(new_n1151), .B1(new_n775), .B2(new_n1085), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n247), .B1(new_n760), .B2(new_n280), .ZN(new_n1178));
  INV_X1    g0978(.A(G128), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n752), .A2(new_n819), .B1(new_n756), .B2(new_n1179), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1178), .B(new_n1180), .C1(G50), .C2(new_n763), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n780), .B2(new_n767), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n1177), .A2(new_n1182), .A3(new_n1141), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n746), .B1(new_n1176), .B2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1184), .B(new_n732), .C1(G68), .C2(new_n1083), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT124), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n871), .B2(new_n744), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n1171), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1168), .A2(new_n1188), .ZN(G381));
  NOR2_X1   g0989(.A1(G393), .A2(G396), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n835), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT125), .Z(new_n1192));
  NOR4_X1   g0992(.A1(new_n1192), .A2(G387), .A3(G390), .A4(G381), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1082), .A2(new_n1105), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n1064), .B2(new_n730), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n961), .B1(new_n1064), .B2(new_n1076), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1195), .B1(new_n1079), .B2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1193), .A2(new_n1197), .A3(new_n1131), .A4(new_n1161), .ZN(G407));
  NOR2_X1   g0998(.A1(new_n651), .A2(G343), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  OAI211_X1 g1000(.A(G407), .B(G213), .C1(G375), .C2(new_n1200), .ZN(G409));
  INV_X1    g1001(.A(KEYINPUT126), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1108), .A2(new_n1163), .A3(KEYINPUT60), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n673), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1076), .A2(KEYINPUT60), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1204), .B1(new_n1166), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1171), .A2(new_n1187), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n835), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1205), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n1209), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1188), .B(G384), .C1(new_n1210), .C2(new_n1204), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1208), .A2(new_n1211), .ZN(new_n1212));
  OAI211_X1 g1012(.A(G378), .B(new_n1161), .C1(new_n1128), .C2(new_n1130), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1161), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1167), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1215), .B(new_n1124), .C1(new_n1079), .C2(new_n1109), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1197), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1199), .B(new_n1212), .C1(new_n1213), .C2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1202), .B1(new_n1218), .B2(KEYINPUT63), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1213), .A2(new_n1217), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1212), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1199), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT63), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1223), .A2(KEYINPUT126), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1218), .A2(KEYINPUT63), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(G387), .A2(new_n1030), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(G387), .A2(new_n1030), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n799), .B1(new_n964), .B2(new_n1000), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n1228), .A2(new_n1229), .B1(new_n1190), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1229), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1190), .A2(new_n1230), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1232), .A2(new_n1233), .A3(new_n1227), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT61), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1231), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1199), .A2(G2897), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1212), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1208), .A2(new_n1211), .A3(new_n1238), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1236), .B1(new_n1237), .B2(new_n1242), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1219), .A2(new_n1225), .A3(new_n1226), .A4(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1223), .A2(KEYINPUT62), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(KEYINPUT127), .B(KEYINPUT61), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1199), .B1(new_n1213), .B2(new_n1217), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1246), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT62), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n1247), .B2(new_n1221), .ZN(new_n1251));
  NOR3_X1   g1051(.A1(new_n1245), .A2(new_n1249), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1231), .A2(new_n1234), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1244), .B1(new_n1252), .B2(new_n1254), .ZN(G405));
  NAND2_X1  g1055(.A1(G375), .A2(new_n1197), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1256), .A2(new_n1213), .A3(new_n1212), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1212), .B1(new_n1256), .B2(new_n1213), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1253), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1259), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1261), .A2(new_n1257), .A3(new_n1254), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1260), .A2(new_n1262), .ZN(G402));
endmodule


