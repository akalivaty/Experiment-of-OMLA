

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U546 ( .A1(G651), .A2(n623), .ZN(n646) );
  XNOR2_X1 U547 ( .A(n713), .B(n712), .ZN(n727) );
  NOR2_X1 U548 ( .A1(n527), .A2(n526), .ZN(G164) );
  NOR2_X1 U549 ( .A1(n520), .A2(n519), .ZN(G160) );
  AND2_X1 U550 ( .A1(n794), .A2(n793), .ZN(n509) );
  AND2_X1 U551 ( .A1(n804), .A2(n791), .ZN(n510) );
  INV_X1 U552 ( .A(n717), .ZN(n694) );
  INV_X1 U553 ( .A(KEYINPUT28), .ZN(n701) );
  XNOR2_X1 U554 ( .A(KEYINPUT31), .B(KEYINPUT95), .ZN(n712) );
  OR2_X1 U555 ( .A1(n729), .A2(n731), .ZN(n714) );
  AND2_X1 U556 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U557 ( .A1(n775), .A2(n670), .ZN(n717) );
  NOR2_X1 U558 ( .A1(n792), .A2(n510), .ZN(n793) );
  AND2_X1 U559 ( .A1(n516), .A2(G2104), .ZN(n881) );
  XNOR2_X1 U560 ( .A(KEYINPUT71), .B(n542), .ZN(G171) );
  XNOR2_X1 U561 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n512) );
  NOR2_X1 U562 ( .A1(G2105), .A2(G2104), .ZN(n511) );
  XNOR2_X2 U563 ( .A(n512), .B(n511), .ZN(n880) );
  NAND2_X1 U564 ( .A1(n880), .A2(G137), .ZN(n515) );
  INV_X1 U565 ( .A(G2105), .ZN(n516) );
  NAND2_X1 U566 ( .A1(G101), .A2(n881), .ZN(n513) );
  XOR2_X1 U567 ( .A(KEYINPUT23), .B(n513), .Z(n514) );
  NAND2_X1 U568 ( .A1(n515), .A2(n514), .ZN(n520) );
  NOR2_X1 U569 ( .A1(G2104), .A2(n516), .ZN(n876) );
  NAND2_X1 U570 ( .A1(G125), .A2(n876), .ZN(n518) );
  AND2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n877) );
  NAND2_X1 U572 ( .A1(G113), .A2(n877), .ZN(n517) );
  NAND2_X1 U573 ( .A1(n518), .A2(n517), .ZN(n519) );
  NAND2_X1 U574 ( .A1(G138), .A2(n880), .ZN(n522) );
  NAND2_X1 U575 ( .A1(G102), .A2(n881), .ZN(n521) );
  NAND2_X1 U576 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U577 ( .A(n523), .B(KEYINPUT90), .ZN(n527) );
  NAND2_X1 U578 ( .A1(G126), .A2(n876), .ZN(n525) );
  NAND2_X1 U579 ( .A1(G114), .A2(n877), .ZN(n524) );
  NAND2_X1 U580 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X2 U581 ( .A1(G651), .A2(G543), .ZN(n638) );
  NAND2_X1 U582 ( .A1(n638), .A2(G90), .ZN(n528) );
  XOR2_X1 U583 ( .A(KEYINPUT69), .B(n528), .Z(n530) );
  XOR2_X1 U584 ( .A(G543), .B(KEYINPUT0), .Z(n623) );
  INV_X1 U585 ( .A(G651), .ZN(n533) );
  NOR2_X1 U586 ( .A1(n623), .A2(n533), .ZN(n642) );
  NAND2_X1 U587 ( .A1(n642), .A2(G77), .ZN(n529) );
  NAND2_X1 U588 ( .A1(n530), .A2(n529), .ZN(n532) );
  XNOR2_X1 U589 ( .A(KEYINPUT70), .B(KEYINPUT9), .ZN(n531) );
  XNOR2_X1 U590 ( .A(n532), .B(n531), .ZN(n541) );
  NOR2_X1 U591 ( .A1(G543), .A2(n533), .ZN(n534) );
  XOR2_X1 U592 ( .A(KEYINPUT66), .B(n534), .Z(n535) );
  XNOR2_X2 U593 ( .A(KEYINPUT1), .B(n535), .ZN(n639) );
  NAND2_X1 U594 ( .A1(G64), .A2(n639), .ZN(n536) );
  XOR2_X1 U595 ( .A(KEYINPUT67), .B(n536), .Z(n538) );
  NAND2_X1 U596 ( .A1(n646), .A2(G52), .ZN(n537) );
  NAND2_X1 U597 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U598 ( .A(KEYINPUT68), .B(n539), .Z(n540) );
  NAND2_X1 U599 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U600 ( .A1(G85), .A2(n638), .ZN(n544) );
  NAND2_X1 U601 ( .A1(G60), .A2(n639), .ZN(n543) );
  NAND2_X1 U602 ( .A1(n544), .A2(n543), .ZN(n548) );
  NAND2_X1 U603 ( .A1(G72), .A2(n642), .ZN(n546) );
  NAND2_X1 U604 ( .A1(G47), .A2(n646), .ZN(n545) );
  NAND2_X1 U605 ( .A1(n546), .A2(n545), .ZN(n547) );
  OR2_X1 U606 ( .A1(n548), .A2(n547), .ZN(G290) );
  AND2_X1 U607 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U608 ( .A(G132), .ZN(G219) );
  INV_X1 U609 ( .A(G82), .ZN(G220) );
  XNOR2_X1 U610 ( .A(KEYINPUT80), .B(KEYINPUT7), .ZN(n560) );
  NAND2_X1 U611 ( .A1(n638), .A2(G89), .ZN(n549) );
  XNOR2_X1 U612 ( .A(n549), .B(KEYINPUT4), .ZN(n551) );
  NAND2_X1 U613 ( .A1(G76), .A2(n642), .ZN(n550) );
  NAND2_X1 U614 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U615 ( .A(KEYINPUT5), .B(n552), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n646), .A2(G51), .ZN(n553) );
  XOR2_X1 U617 ( .A(KEYINPUT79), .B(n553), .Z(n555) );
  NAND2_X1 U618 ( .A1(G63), .A2(n639), .ZN(n554) );
  NAND2_X1 U619 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U620 ( .A(KEYINPUT6), .B(n556), .Z(n557) );
  NAND2_X1 U621 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U622 ( .A(n560), .B(n559), .ZN(G168) );
  XOR2_X1 U623 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U624 ( .A1(G7), .A2(G661), .ZN(n561) );
  XNOR2_X1 U625 ( .A(n561), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U626 ( .A(G223), .ZN(n819) );
  NAND2_X1 U627 ( .A1(n819), .A2(G567), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(KEYINPUT11), .ZN(n563) );
  XNOR2_X1 U629 ( .A(KEYINPUT73), .B(n563), .ZN(G234) );
  NAND2_X1 U630 ( .A1(n638), .A2(G81), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(KEYINPUT12), .ZN(n566) );
  NAND2_X1 U632 ( .A1(G68), .A2(n642), .ZN(n565) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(KEYINPUT13), .B(n567), .ZN(n574) );
  XOR2_X1 U635 ( .A(KEYINPUT74), .B(KEYINPUT14), .Z(n569) );
  NAND2_X1 U636 ( .A1(G56), .A2(n639), .ZN(n568) );
  XNOR2_X1 U637 ( .A(n569), .B(n568), .ZN(n572) );
  NAND2_X1 U638 ( .A1(G43), .A2(n646), .ZN(n570) );
  XNOR2_X1 U639 ( .A(KEYINPUT75), .B(n570), .ZN(n571) );
  NOR2_X1 U640 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n908) );
  INV_X1 U642 ( .A(G860), .ZN(n595) );
  OR2_X1 U643 ( .A1(n908), .A2(n595), .ZN(G153) );
  XOR2_X1 U644 ( .A(G171), .B(KEYINPUT76), .Z(G301) );
  NAND2_X1 U645 ( .A1(G868), .A2(G301), .ZN(n575) );
  XOR2_X1 U646 ( .A(KEYINPUT77), .B(n575), .Z(n585) );
  NAND2_X1 U647 ( .A1(G79), .A2(n642), .ZN(n577) );
  NAND2_X1 U648 ( .A1(G66), .A2(n639), .ZN(n576) );
  AND2_X1 U649 ( .A1(n577), .A2(n576), .ZN(n582) );
  NAND2_X1 U650 ( .A1(n638), .A2(G92), .ZN(n578) );
  XOR2_X1 U651 ( .A(KEYINPUT78), .B(n578), .Z(n580) );
  AND2_X1 U652 ( .A1(n646), .A2(G54), .ZN(n579) );
  NOR2_X1 U653 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U654 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X2 U655 ( .A(KEYINPUT15), .B(n583), .Z(n913) );
  INV_X1 U656 ( .A(G868), .ZN(n592) );
  NAND2_X1 U657 ( .A1(n913), .A2(n592), .ZN(n584) );
  NAND2_X1 U658 ( .A1(n585), .A2(n584), .ZN(G284) );
  NAND2_X1 U659 ( .A1(G91), .A2(n638), .ZN(n587) );
  NAND2_X1 U660 ( .A1(G78), .A2(n642), .ZN(n586) );
  NAND2_X1 U661 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U662 ( .A1(n646), .A2(G53), .ZN(n589) );
  NAND2_X1 U663 ( .A1(G65), .A2(n639), .ZN(n588) );
  NAND2_X1 U664 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U665 ( .A1(n591), .A2(n590), .ZN(n907) );
  INV_X1 U666 ( .A(n907), .ZN(G299) );
  NAND2_X1 U667 ( .A1(G868), .A2(G286), .ZN(n594) );
  NAND2_X1 U668 ( .A1(G299), .A2(n592), .ZN(n593) );
  NAND2_X1 U669 ( .A1(n594), .A2(n593), .ZN(G297) );
  NAND2_X1 U670 ( .A1(n595), .A2(G559), .ZN(n596) );
  INV_X1 U671 ( .A(n913), .ZN(n619) );
  NAND2_X1 U672 ( .A1(n596), .A2(n619), .ZN(n597) );
  XNOR2_X1 U673 ( .A(n597), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U674 ( .A1(G868), .A2(n908), .ZN(n600) );
  NAND2_X1 U675 ( .A1(G868), .A2(n619), .ZN(n598) );
  NOR2_X1 U676 ( .A1(G559), .A2(n598), .ZN(n599) );
  NOR2_X1 U677 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U678 ( .A(KEYINPUT81), .B(n601), .Z(G282) );
  XOR2_X1 U679 ( .A(G2100), .B(KEYINPUT82), .Z(n610) );
  NAND2_X1 U680 ( .A1(G123), .A2(n876), .ZN(n602) );
  XNOR2_X1 U681 ( .A(n602), .B(KEYINPUT18), .ZN(n604) );
  NAND2_X1 U682 ( .A1(n881), .A2(G99), .ZN(n603) );
  NAND2_X1 U683 ( .A1(n604), .A2(n603), .ZN(n608) );
  NAND2_X1 U684 ( .A1(G135), .A2(n880), .ZN(n606) );
  NAND2_X1 U685 ( .A1(G111), .A2(n877), .ZN(n605) );
  NAND2_X1 U686 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U687 ( .A1(n608), .A2(n607), .ZN(n989) );
  XNOR2_X1 U688 ( .A(G2096), .B(n989), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n609), .ZN(G156) );
  NAND2_X1 U690 ( .A1(n646), .A2(G55), .ZN(n612) );
  NAND2_X1 U691 ( .A1(G67), .A2(n639), .ZN(n611) );
  NAND2_X1 U692 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U693 ( .A(KEYINPUT85), .B(n613), .ZN(n618) );
  NAND2_X1 U694 ( .A1(G93), .A2(n638), .ZN(n615) );
  NAND2_X1 U695 ( .A1(G80), .A2(n642), .ZN(n614) );
  NAND2_X1 U696 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U697 ( .A(KEYINPUT84), .B(n616), .Z(n617) );
  NAND2_X1 U698 ( .A1(n618), .A2(n617), .ZN(n892) );
  NAND2_X1 U699 ( .A1(G559), .A2(n619), .ZN(n620) );
  XOR2_X1 U700 ( .A(KEYINPUT83), .B(n620), .Z(n655) );
  XNOR2_X1 U701 ( .A(n908), .B(n655), .ZN(n621) );
  NOR2_X1 U702 ( .A1(G860), .A2(n621), .ZN(n622) );
  XOR2_X1 U703 ( .A(n892), .B(n622), .Z(G145) );
  NAND2_X1 U704 ( .A1(G87), .A2(n623), .ZN(n624) );
  XNOR2_X1 U705 ( .A(n624), .B(KEYINPUT86), .ZN(n629) );
  NAND2_X1 U706 ( .A1(G49), .A2(n646), .ZN(n626) );
  NAND2_X1 U707 ( .A1(G74), .A2(G651), .ZN(n625) );
  NAND2_X1 U708 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U709 ( .A1(n639), .A2(n627), .ZN(n628) );
  NAND2_X1 U710 ( .A1(n629), .A2(n628), .ZN(G288) );
  NAND2_X1 U711 ( .A1(G88), .A2(n638), .ZN(n630) );
  XNOR2_X1 U712 ( .A(n630), .B(KEYINPUT88), .ZN(n637) );
  NAND2_X1 U713 ( .A1(G75), .A2(n642), .ZN(n632) );
  NAND2_X1 U714 ( .A1(G62), .A2(n639), .ZN(n631) );
  NAND2_X1 U715 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U716 ( .A1(G50), .A2(n646), .ZN(n633) );
  XNOR2_X1 U717 ( .A(KEYINPUT87), .B(n633), .ZN(n634) );
  NOR2_X1 U718 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U719 ( .A1(n637), .A2(n636), .ZN(G303) );
  NAND2_X1 U720 ( .A1(G86), .A2(n638), .ZN(n641) );
  NAND2_X1 U721 ( .A1(G61), .A2(n639), .ZN(n640) );
  NAND2_X1 U722 ( .A1(n641), .A2(n640), .ZN(n645) );
  NAND2_X1 U723 ( .A1(n642), .A2(G73), .ZN(n643) );
  XOR2_X1 U724 ( .A(KEYINPUT2), .B(n643), .Z(n644) );
  NOR2_X1 U725 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U726 ( .A1(n646), .A2(G48), .ZN(n647) );
  NAND2_X1 U727 ( .A1(n648), .A2(n647), .ZN(G305) );
  XNOR2_X1 U728 ( .A(n907), .B(G288), .ZN(n651) );
  XNOR2_X1 U729 ( .A(n908), .B(G303), .ZN(n649) );
  XNOR2_X1 U730 ( .A(n649), .B(G305), .ZN(n650) );
  XNOR2_X1 U731 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U732 ( .A(KEYINPUT89), .B(n652), .ZN(n654) );
  XNOR2_X1 U733 ( .A(G290), .B(KEYINPUT19), .ZN(n653) );
  XNOR2_X1 U734 ( .A(n654), .B(n653), .ZN(n891) );
  XNOR2_X1 U735 ( .A(n891), .B(n655), .ZN(n656) );
  NAND2_X1 U736 ( .A1(n656), .A2(G868), .ZN(n657) );
  XNOR2_X1 U737 ( .A(n892), .B(n657), .ZN(G295) );
  NAND2_X1 U738 ( .A1(G2084), .A2(G2078), .ZN(n658) );
  XOR2_X1 U739 ( .A(KEYINPUT20), .B(n658), .Z(n659) );
  NAND2_X1 U740 ( .A1(G2090), .A2(n659), .ZN(n660) );
  XNOR2_X1 U741 ( .A(KEYINPUT21), .B(n660), .ZN(n661) );
  NAND2_X1 U742 ( .A1(n661), .A2(G2072), .ZN(G158) );
  XOR2_X1 U743 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  XNOR2_X1 U744 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U745 ( .A1(G108), .A2(G120), .ZN(n662) );
  NOR2_X1 U746 ( .A1(G237), .A2(n662), .ZN(n663) );
  NAND2_X1 U747 ( .A1(G69), .A2(n663), .ZN(n823) );
  NAND2_X1 U748 ( .A1(n823), .A2(G567), .ZN(n668) );
  NOR2_X1 U749 ( .A1(G220), .A2(G219), .ZN(n664) );
  XOR2_X1 U750 ( .A(KEYINPUT22), .B(n664), .Z(n665) );
  NOR2_X1 U751 ( .A1(G218), .A2(n665), .ZN(n666) );
  NAND2_X1 U752 ( .A1(G96), .A2(n666), .ZN(n824) );
  NAND2_X1 U753 ( .A1(n824), .A2(G2106), .ZN(n667) );
  NAND2_X1 U754 ( .A1(n668), .A2(n667), .ZN(n825) );
  NAND2_X1 U755 ( .A1(G661), .A2(G483), .ZN(n669) );
  NOR2_X1 U756 ( .A1(n825), .A2(n669), .ZN(n822) );
  NAND2_X1 U757 ( .A1(n822), .A2(G36), .ZN(G176) );
  NOR2_X1 U758 ( .A1(G164), .A2(G1384), .ZN(n775) );
  NAND2_X1 U759 ( .A1(G160), .A2(G40), .ZN(n774) );
  INV_X1 U760 ( .A(n774), .ZN(n670) );
  NAND2_X1 U761 ( .A1(G8), .A2(n717), .ZN(n760) );
  NOR2_X1 U762 ( .A1(G1981), .A2(G305), .ZN(n671) );
  XOR2_X1 U763 ( .A(n671), .B(KEYINPUT24), .Z(n672) );
  NOR2_X1 U764 ( .A1(n760), .A2(n672), .ZN(n754) );
  XNOR2_X1 U765 ( .A(G1981), .B(G305), .ZN(n905) );
  XNOR2_X1 U766 ( .A(G2078), .B(KEYINPUT25), .ZN(n933) );
  NOR2_X1 U767 ( .A1(n717), .A2(n933), .ZN(n674) );
  AND2_X1 U768 ( .A1(n717), .A2(G1961), .ZN(n673) );
  NOR2_X1 U769 ( .A1(n674), .A2(n673), .ZN(n709) );
  AND2_X1 U770 ( .A1(G171), .A2(n709), .ZN(n729) );
  NAND2_X1 U771 ( .A1(G1348), .A2(n717), .ZN(n676) );
  NAND2_X1 U772 ( .A1(G2067), .A2(n694), .ZN(n675) );
  NAND2_X1 U773 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U774 ( .A1(n913), .A2(n677), .ZN(n693) );
  AND2_X1 U775 ( .A1(G1348), .A2(n913), .ZN(n680) );
  XNOR2_X1 U776 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n685) );
  INV_X1 U777 ( .A(G1341), .ZN(n678) );
  NAND2_X1 U778 ( .A1(n685), .A2(n678), .ZN(n679) );
  NOR2_X1 U779 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U780 ( .A1(n694), .A2(n681), .ZN(n691) );
  NAND2_X1 U781 ( .A1(n913), .A2(G2067), .ZN(n683) );
  NAND2_X1 U782 ( .A1(G1996), .A2(n685), .ZN(n682) );
  NAND2_X1 U783 ( .A1(n683), .A2(n682), .ZN(n684) );
  AND2_X1 U784 ( .A1(n684), .A2(n694), .ZN(n689) );
  OR2_X1 U785 ( .A1(G1996), .A2(n685), .ZN(n687) );
  INV_X1 U786 ( .A(n908), .ZN(n686) );
  NAND2_X1 U787 ( .A1(n687), .A2(n686), .ZN(n688) );
  OR2_X1 U788 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U789 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U790 ( .A1(n693), .A2(n692), .ZN(n699) );
  NAND2_X1 U791 ( .A1(n694), .A2(G2072), .ZN(n695) );
  XNOR2_X1 U792 ( .A(n695), .B(KEYINPUT27), .ZN(n697) );
  AND2_X1 U793 ( .A1(G1956), .A2(n717), .ZN(n696) );
  NOR2_X1 U794 ( .A1(n697), .A2(n696), .ZN(n700) );
  NAND2_X1 U795 ( .A1(n700), .A2(n907), .ZN(n698) );
  NAND2_X1 U796 ( .A1(n699), .A2(n698), .ZN(n704) );
  NOR2_X1 U797 ( .A1(n700), .A2(n907), .ZN(n702) );
  XNOR2_X1 U798 ( .A(n702), .B(n701), .ZN(n703) );
  NAND2_X1 U799 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U800 ( .A(KEYINPUT29), .B(n705), .ZN(n731) );
  NOR2_X1 U801 ( .A1(G2084), .A2(n717), .ZN(n735) );
  NOR2_X1 U802 ( .A1(G1966), .A2(n760), .ZN(n728) );
  NOR2_X1 U803 ( .A1(n735), .A2(n728), .ZN(n706) );
  NAND2_X1 U804 ( .A1(G8), .A2(n706), .ZN(n707) );
  XNOR2_X1 U805 ( .A(n707), .B(KEYINPUT30), .ZN(n708) );
  NOR2_X1 U806 ( .A1(G168), .A2(n708), .ZN(n711) );
  NOR2_X1 U807 ( .A1(G171), .A2(n709), .ZN(n710) );
  NOR2_X1 U808 ( .A1(n711), .A2(n710), .ZN(n713) );
  NAND2_X1 U809 ( .A1(n714), .A2(n727), .ZN(n716) );
  AND2_X1 U810 ( .A1(G286), .A2(G8), .ZN(n715) );
  NAND2_X1 U811 ( .A1(n716), .A2(n715), .ZN(n724) );
  INV_X1 U812 ( .A(G8), .ZN(n722) );
  NOR2_X1 U813 ( .A1(G1971), .A2(n760), .ZN(n719) );
  NOR2_X1 U814 ( .A1(G2090), .A2(n717), .ZN(n718) );
  NOR2_X1 U815 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U816 ( .A1(n720), .A2(G303), .ZN(n721) );
  OR2_X1 U817 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U818 ( .A(n725), .B(KEYINPUT32), .ZN(n755) );
  NAND2_X1 U819 ( .A1(G1976), .A2(G288), .ZN(n922) );
  INV_X1 U820 ( .A(n760), .ZN(n747) );
  NAND2_X1 U821 ( .A1(n922), .A2(n747), .ZN(n741) );
  INV_X1 U822 ( .A(n741), .ZN(n726) );
  AND2_X1 U823 ( .A1(n755), .A2(n726), .ZN(n738) );
  OR2_X1 U824 ( .A1(n728), .A2(n727), .ZN(n733) );
  OR2_X1 U825 ( .A1(n729), .A2(n728), .ZN(n730) );
  OR2_X1 U826 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U827 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U828 ( .A(n734), .B(KEYINPUT96), .ZN(n737) );
  NAND2_X1 U829 ( .A1(n735), .A2(G8), .ZN(n736) );
  NAND2_X1 U830 ( .A1(n737), .A2(n736), .ZN(n756) );
  NAND2_X1 U831 ( .A1(n738), .A2(n756), .ZN(n743) );
  NOR2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n919) );
  NOR2_X1 U833 ( .A1(G1971), .A2(G303), .ZN(n739) );
  NOR2_X1 U834 ( .A1(n919), .A2(n739), .ZN(n740) );
  OR2_X1 U835 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U836 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U837 ( .A(n744), .B(KEYINPUT64), .ZN(n746) );
  INV_X1 U838 ( .A(KEYINPUT33), .ZN(n745) );
  NAND2_X1 U839 ( .A1(n746), .A2(n745), .ZN(n750) );
  NAND2_X1 U840 ( .A1(n919), .A2(n747), .ZN(n748) );
  NAND2_X1 U841 ( .A1(n748), .A2(KEYINPUT33), .ZN(n749) );
  NAND2_X1 U842 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U843 ( .A(n751), .B(KEYINPUT97), .ZN(n752) );
  NOR2_X1 U844 ( .A1(n905), .A2(n752), .ZN(n753) );
  NOR2_X1 U845 ( .A1(n754), .A2(n753), .ZN(n763) );
  NAND2_X1 U846 ( .A1(n756), .A2(n755), .ZN(n759) );
  NOR2_X1 U847 ( .A1(G2090), .A2(G303), .ZN(n757) );
  NAND2_X1 U848 ( .A1(G8), .A2(n757), .ZN(n758) );
  NAND2_X1 U849 ( .A1(n759), .A2(n758), .ZN(n761) );
  NAND2_X1 U850 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U851 ( .A1(n763), .A2(n762), .ZN(n794) );
  XNOR2_X1 U852 ( .A(KEYINPUT37), .B(G2067), .ZN(n802) );
  NAND2_X1 U853 ( .A1(n881), .A2(G104), .ZN(n764) );
  XOR2_X1 U854 ( .A(KEYINPUT91), .B(n764), .Z(n766) );
  NAND2_X1 U855 ( .A1(n880), .A2(G140), .ZN(n765) );
  NAND2_X1 U856 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U857 ( .A(KEYINPUT34), .B(n767), .ZN(n772) );
  NAND2_X1 U858 ( .A1(G128), .A2(n876), .ZN(n769) );
  NAND2_X1 U859 ( .A1(G116), .A2(n877), .ZN(n768) );
  NAND2_X1 U860 ( .A1(n769), .A2(n768), .ZN(n770) );
  XOR2_X1 U861 ( .A(KEYINPUT35), .B(n770), .Z(n771) );
  NOR2_X1 U862 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U863 ( .A(KEYINPUT36), .B(n773), .ZN(n865) );
  NOR2_X1 U864 ( .A1(n802), .A2(n865), .ZN(n1010) );
  NOR2_X1 U865 ( .A1(n775), .A2(n774), .ZN(n804) );
  NAND2_X1 U866 ( .A1(n1010), .A2(n804), .ZN(n776) );
  XNOR2_X1 U867 ( .A(n776), .B(KEYINPUT92), .ZN(n800) );
  INV_X1 U868 ( .A(n800), .ZN(n792) );
  NAND2_X1 U869 ( .A1(G141), .A2(n880), .ZN(n778) );
  NAND2_X1 U870 ( .A1(G129), .A2(n876), .ZN(n777) );
  NAND2_X1 U871 ( .A1(n778), .A2(n777), .ZN(n781) );
  NAND2_X1 U872 ( .A1(n881), .A2(G105), .ZN(n779) );
  XOR2_X1 U873 ( .A(KEYINPUT38), .B(n779), .Z(n780) );
  NOR2_X1 U874 ( .A1(n781), .A2(n780), .ZN(n783) );
  NAND2_X1 U875 ( .A1(n877), .A2(G117), .ZN(n782) );
  NAND2_X1 U876 ( .A1(n783), .A2(n782), .ZN(n871) );
  AND2_X1 U877 ( .A1(n871), .A2(G1996), .ZN(n990) );
  NAND2_X1 U878 ( .A1(G131), .A2(n880), .ZN(n785) );
  NAND2_X1 U879 ( .A1(G95), .A2(n881), .ZN(n784) );
  NAND2_X1 U880 ( .A1(n785), .A2(n784), .ZN(n790) );
  NAND2_X1 U881 ( .A1(G119), .A2(n876), .ZN(n787) );
  NAND2_X1 U882 ( .A1(G107), .A2(n877), .ZN(n786) );
  NAND2_X1 U883 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U884 ( .A(KEYINPUT93), .B(n788), .Z(n789) );
  OR2_X1 U885 ( .A1(n790), .A2(n789), .ZN(n864) );
  AND2_X1 U886 ( .A1(n864), .A2(G1991), .ZN(n988) );
  OR2_X1 U887 ( .A1(n990), .A2(n988), .ZN(n791) );
  XNOR2_X1 U888 ( .A(G1986), .B(G290), .ZN(n910) );
  NAND2_X1 U889 ( .A1(n910), .A2(n804), .ZN(n795) );
  NAND2_X1 U890 ( .A1(n509), .A2(n795), .ZN(n807) );
  NOR2_X1 U891 ( .A1(G1996), .A2(n871), .ZN(n992) );
  NOR2_X1 U892 ( .A1(G1991), .A2(n864), .ZN(n998) );
  NOR2_X1 U893 ( .A1(G1986), .A2(G290), .ZN(n796) );
  NOR2_X1 U894 ( .A1(n998), .A2(n796), .ZN(n797) );
  NOR2_X1 U895 ( .A1(n510), .A2(n797), .ZN(n798) );
  NOR2_X1 U896 ( .A1(n992), .A2(n798), .ZN(n799) );
  XNOR2_X1 U897 ( .A(n799), .B(KEYINPUT39), .ZN(n801) );
  NAND2_X1 U898 ( .A1(n801), .A2(n800), .ZN(n803) );
  NAND2_X1 U899 ( .A1(n802), .A2(n865), .ZN(n1007) );
  NAND2_X1 U900 ( .A1(n803), .A2(n1007), .ZN(n805) );
  NAND2_X1 U901 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U902 ( .A1(n807), .A2(n806), .ZN(n809) );
  XNOR2_X1 U903 ( .A(KEYINPUT40), .B(KEYINPUT98), .ZN(n808) );
  XNOR2_X1 U904 ( .A(n809), .B(n808), .ZN(G329) );
  XNOR2_X1 U905 ( .A(G1341), .B(G2454), .ZN(n810) );
  XNOR2_X1 U906 ( .A(n810), .B(G2430), .ZN(n811) );
  XNOR2_X1 U907 ( .A(n811), .B(G1348), .ZN(n817) );
  XOR2_X1 U908 ( .A(G2443), .B(G2427), .Z(n813) );
  XNOR2_X1 U909 ( .A(G2438), .B(G2446), .ZN(n812) );
  XNOR2_X1 U910 ( .A(n813), .B(n812), .ZN(n815) );
  XOR2_X1 U911 ( .A(G2451), .B(G2435), .Z(n814) );
  XNOR2_X1 U912 ( .A(n815), .B(n814), .ZN(n816) );
  XNOR2_X1 U913 ( .A(n817), .B(n816), .ZN(n818) );
  NAND2_X1 U914 ( .A1(n818), .A2(G14), .ZN(n897) );
  XNOR2_X1 U915 ( .A(KEYINPUT99), .B(n897), .ZN(G401) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n819), .ZN(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n820) );
  NAND2_X1 U918 ( .A1(G661), .A2(n820), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n821) );
  NAND2_X1 U920 ( .A1(n822), .A2(n821), .ZN(G188) );
  NOR2_X1 U921 ( .A1(n824), .A2(n823), .ZN(G325) );
  XOR2_X1 U922 ( .A(KEYINPUT100), .B(G325), .Z(G261) );
  INV_X1 U924 ( .A(G120), .ZN(G236) );
  INV_X1 U925 ( .A(G108), .ZN(G238) );
  INV_X1 U926 ( .A(G96), .ZN(G221) );
  INV_X1 U927 ( .A(G69), .ZN(G235) );
  INV_X1 U928 ( .A(n825), .ZN(G319) );
  XOR2_X1 U929 ( .A(KEYINPUT41), .B(G1976), .Z(n827) );
  XNOR2_X1 U930 ( .A(G1961), .B(G1971), .ZN(n826) );
  XNOR2_X1 U931 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U932 ( .A(n828), .B(KEYINPUT104), .Z(n830) );
  XNOR2_X1 U933 ( .A(G1996), .B(G1991), .ZN(n829) );
  XNOR2_X1 U934 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U935 ( .A(G1981), .B(G1956), .Z(n832) );
  XNOR2_X1 U936 ( .A(G1986), .B(G1966), .ZN(n831) );
  XNOR2_X1 U937 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U938 ( .A(n834), .B(n833), .Z(n836) );
  XNOR2_X1 U939 ( .A(KEYINPUT103), .B(G2474), .ZN(n835) );
  XNOR2_X1 U940 ( .A(n836), .B(n835), .ZN(G229) );
  XOR2_X1 U941 ( .A(KEYINPUT43), .B(KEYINPUT102), .Z(n838) );
  XNOR2_X1 U942 ( .A(KEYINPUT101), .B(G2678), .ZN(n837) );
  XNOR2_X1 U943 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U944 ( .A(KEYINPUT42), .B(G2090), .Z(n840) );
  XNOR2_X1 U945 ( .A(G2067), .B(G2072), .ZN(n839) );
  XNOR2_X1 U946 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U947 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U948 ( .A(G2100), .B(G2096), .ZN(n843) );
  XNOR2_X1 U949 ( .A(n844), .B(n843), .ZN(n846) );
  XOR2_X1 U950 ( .A(G2084), .B(G2078), .Z(n845) );
  XNOR2_X1 U951 ( .A(n846), .B(n845), .ZN(G227) );
  NAND2_X1 U952 ( .A1(G124), .A2(n876), .ZN(n847) );
  XNOR2_X1 U953 ( .A(n847), .B(KEYINPUT44), .ZN(n849) );
  NAND2_X1 U954 ( .A1(n881), .A2(G100), .ZN(n848) );
  NAND2_X1 U955 ( .A1(n849), .A2(n848), .ZN(n853) );
  NAND2_X1 U956 ( .A1(G136), .A2(n880), .ZN(n851) );
  NAND2_X1 U957 ( .A1(G112), .A2(n877), .ZN(n850) );
  NAND2_X1 U958 ( .A1(n851), .A2(n850), .ZN(n852) );
  NOR2_X1 U959 ( .A1(n853), .A2(n852), .ZN(G162) );
  NAND2_X1 U960 ( .A1(G127), .A2(n876), .ZN(n856) );
  NAND2_X1 U961 ( .A1(n877), .A2(G115), .ZN(n854) );
  XOR2_X1 U962 ( .A(KEYINPUT105), .B(n854), .Z(n855) );
  NAND2_X1 U963 ( .A1(n856), .A2(n855), .ZN(n859) );
  XNOR2_X1 U964 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n857) );
  XNOR2_X1 U965 ( .A(n857), .B(KEYINPUT47), .ZN(n858) );
  XNOR2_X1 U966 ( .A(n859), .B(n858), .ZN(n863) );
  NAND2_X1 U967 ( .A1(G139), .A2(n880), .ZN(n861) );
  NAND2_X1 U968 ( .A1(G103), .A2(n881), .ZN(n860) );
  NAND2_X1 U969 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U970 ( .A1(n863), .A2(n862), .ZN(n1001) );
  XNOR2_X1 U971 ( .A(n1001), .B(G162), .ZN(n867) );
  XOR2_X1 U972 ( .A(n865), .B(n864), .Z(n866) );
  XNOR2_X1 U973 ( .A(n867), .B(n866), .ZN(n875) );
  XOR2_X1 U974 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n869) );
  XNOR2_X1 U975 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n868) );
  XNOR2_X1 U976 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U977 ( .A(n870), .B(n989), .Z(n873) );
  XOR2_X1 U978 ( .A(G160), .B(n871), .Z(n872) );
  XNOR2_X1 U979 ( .A(n873), .B(n872), .ZN(n874) );
  XOR2_X1 U980 ( .A(n875), .B(n874), .Z(n889) );
  NAND2_X1 U981 ( .A1(G130), .A2(n876), .ZN(n879) );
  NAND2_X1 U982 ( .A1(G118), .A2(n877), .ZN(n878) );
  NAND2_X1 U983 ( .A1(n879), .A2(n878), .ZN(n886) );
  NAND2_X1 U984 ( .A1(G142), .A2(n880), .ZN(n883) );
  NAND2_X1 U985 ( .A1(G106), .A2(n881), .ZN(n882) );
  NAND2_X1 U986 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U987 ( .A(KEYINPUT45), .B(n884), .Z(n885) );
  NOR2_X1 U988 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U989 ( .A(G164), .B(n887), .ZN(n888) );
  XNOR2_X1 U990 ( .A(n889), .B(n888), .ZN(n890) );
  NOR2_X1 U991 ( .A1(G37), .A2(n890), .ZN(G395) );
  XNOR2_X1 U992 ( .A(n891), .B(n913), .ZN(n893) );
  XNOR2_X1 U993 ( .A(n893), .B(n892), .ZN(n895) );
  XOR2_X1 U994 ( .A(G286), .B(G171), .Z(n894) );
  XNOR2_X1 U995 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U996 ( .A1(G37), .A2(n896), .ZN(G397) );
  NAND2_X1 U997 ( .A1(G319), .A2(n897), .ZN(n900) );
  NOR2_X1 U998 ( .A1(G229), .A2(G227), .ZN(n898) );
  XNOR2_X1 U999 ( .A(n898), .B(KEYINPUT49), .ZN(n899) );
  NOR2_X1 U1000 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(KEYINPUT110), .B(n901), .ZN(n903) );
  NOR2_X1 U1002 ( .A1(G395), .A2(G397), .ZN(n902) );
  NAND2_X1 U1003 ( .A1(n903), .A2(n902), .ZN(G225) );
  INV_X1 U1004 ( .A(G225), .ZN(G308) );
  INV_X1 U1005 ( .A(G303), .ZN(G166) );
  XOR2_X1 U1006 ( .A(G1966), .B(G168), .Z(n904) );
  NOR2_X1 U1007 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U1008 ( .A(KEYINPUT57), .B(n906), .ZN(n929) );
  XNOR2_X1 U1009 ( .A(G171), .B(G1961), .ZN(n918) );
  XNOR2_X1 U1010 ( .A(n907), .B(G1956), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(G1341), .B(n908), .ZN(n909) );
  NOR2_X1 U1012 ( .A1(n910), .A2(n909), .ZN(n911) );
  NAND2_X1 U1013 ( .A1(n912), .A2(n911), .ZN(n916) );
  XNOR2_X1 U1014 ( .A(G1348), .B(n913), .ZN(n914) );
  XNOR2_X1 U1015 ( .A(KEYINPUT120), .B(n914), .ZN(n915) );
  NOR2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n926) );
  XOR2_X1 U1018 ( .A(n919), .B(KEYINPUT121), .Z(n921) );
  XOR2_X1 U1019 ( .A(G166), .B(G1971), .Z(n920) );
  NOR2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n923) );
  NAND2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1022 ( .A(KEYINPUT122), .B(n924), .ZN(n925) );
  NOR2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(KEYINPUT123), .B(n927), .ZN(n928) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n931) );
  XOR2_X1 U1026 ( .A(KEYINPUT56), .B(G16), .Z(n930) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n958) );
  XOR2_X1 U1028 ( .A(KEYINPUT55), .B(KEYINPUT117), .Z(n952) );
  XNOR2_X1 U1029 ( .A(G2090), .B(G35), .ZN(n946) );
  XOR2_X1 U1030 ( .A(G25), .B(G1991), .Z(n932) );
  NAND2_X1 U1031 ( .A1(n932), .A2(G28), .ZN(n943) );
  XNOR2_X1 U1032 ( .A(G27), .B(n933), .ZN(n937) );
  XNOR2_X1 U1033 ( .A(G2067), .B(G26), .ZN(n935) );
  XNOR2_X1 U1034 ( .A(G32), .B(G1996), .ZN(n934) );
  NOR2_X1 U1035 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n940) );
  XNOR2_X1 U1037 ( .A(KEYINPUT114), .B(G2072), .ZN(n938) );
  XNOR2_X1 U1038 ( .A(G33), .B(n938), .ZN(n939) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1040 ( .A(n941), .B(KEYINPUT115), .ZN(n942) );
  NOR2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1042 ( .A(KEYINPUT53), .B(n944), .ZN(n945) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n950) );
  XOR2_X1 U1044 ( .A(KEYINPUT116), .B(G34), .Z(n948) );
  XNOR2_X1 U1045 ( .A(G2084), .B(KEYINPUT54), .ZN(n947) );
  XNOR2_X1 U1046 ( .A(n948), .B(n947), .ZN(n949) );
  NAND2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1048 ( .A(n952), .B(n951), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(G29), .A2(n953), .ZN(n954) );
  XOR2_X1 U1050 ( .A(KEYINPUT118), .B(n954), .Z(n955) );
  NAND2_X1 U1051 ( .A1(G11), .A2(n955), .ZN(n956) );
  XOR2_X1 U1052 ( .A(KEYINPUT119), .B(n956), .Z(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n984) );
  XOR2_X1 U1054 ( .A(G16), .B(KEYINPUT124), .Z(n982) );
  XNOR2_X1 U1055 ( .A(G1348), .B(KEYINPUT59), .ZN(n959) );
  XNOR2_X1 U1056 ( .A(n959), .B(G4), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(G1956), .B(G20), .ZN(n961) );
  XNOR2_X1 U1058 ( .A(G6), .B(G1981), .ZN(n960) );
  NOR2_X1 U1059 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n966) );
  XOR2_X1 U1061 ( .A(KEYINPUT125), .B(G1341), .Z(n964) );
  XNOR2_X1 U1062 ( .A(G19), .B(n964), .ZN(n965) );
  NOR2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1064 ( .A(KEYINPUT60), .B(n967), .ZN(n968) );
  XNOR2_X1 U1065 ( .A(n968), .B(KEYINPUT126), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(G1966), .B(G21), .ZN(n970) );
  XNOR2_X1 U1067 ( .A(G5), .B(G1961), .ZN(n969) );
  NOR2_X1 U1068 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n979) );
  XNOR2_X1 U1070 ( .A(G1971), .B(G22), .ZN(n974) );
  XNOR2_X1 U1071 ( .A(G23), .B(G1976), .ZN(n973) );
  NOR2_X1 U1072 ( .A1(n974), .A2(n973), .ZN(n976) );
  XOR2_X1 U1073 ( .A(G1986), .B(G24), .Z(n975) );
  NAND2_X1 U1074 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1075 ( .A(KEYINPUT58), .B(n977), .ZN(n978) );
  NOR2_X1 U1076 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1077 ( .A(n980), .B(KEYINPUT61), .ZN(n981) );
  NAND2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1080 ( .A(n985), .B(KEYINPUT127), .ZN(n1016) );
  XNOR2_X1 U1081 ( .A(KEYINPUT52), .B(KEYINPUT113), .ZN(n1012) );
  XNOR2_X1 U1082 ( .A(G160), .B(G2084), .ZN(n986) );
  XNOR2_X1 U1083 ( .A(n986), .B(KEYINPUT111), .ZN(n987) );
  NOR2_X1 U1084 ( .A1(n988), .A2(n987), .ZN(n1000) );
  NOR2_X1 U1085 ( .A1(n990), .A2(n989), .ZN(n996) );
  XOR2_X1 U1086 ( .A(G2090), .B(G162), .Z(n991) );
  XNOR2_X1 U1087 ( .A(KEYINPUT112), .B(n991), .ZN(n993) );
  NOR2_X1 U1088 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1089 ( .A(KEYINPUT51), .B(n994), .Z(n995) );
  NAND2_X1 U1090 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1091 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1006) );
  XOR2_X1 U1093 ( .A(G2072), .B(n1001), .Z(n1003) );
  XOR2_X1 U1094 ( .A(G164), .B(G2078), .Z(n1002) );
  NOR2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1096 ( .A(KEYINPUT50), .B(n1004), .Z(n1005) );
  NOR2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  NAND2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(n1012), .B(n1011), .ZN(n1013) );
  OR2_X1 U1101 ( .A1(KEYINPUT55), .A2(n1013), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(G29), .A2(n1014), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1104 ( .A(KEYINPUT62), .B(n1017), .Z(G311) );
  INV_X1 U1105 ( .A(G311), .ZN(G150) );
endmodule

