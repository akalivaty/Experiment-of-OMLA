//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1243, new_n1244, new_n1245;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n202), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0003(.A(KEYINPUT65), .ZN(new_n204));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  OAI21_X1  g0005(.A(new_n204), .B1(new_n205), .B2(G13), .ZN(new_n206));
  INV_X1    g0006(.A(G13), .ZN(new_n207));
  NAND4_X1  g0007(.A1(new_n207), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(KEYINPUT66), .B(KEYINPUT0), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n210), .B(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  INV_X1    g0017(.A(G97), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI22_X1  g0019(.A1(new_n216), .A2(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI211_X1 g0020(.A(new_n215), .B(new_n220), .C1(G107), .C2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G116), .A2(G270), .ZN(new_n222));
  AND2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G50), .ZN(new_n224));
  INV_X1    g0024(.A(G226), .ZN(new_n225));
  INV_X1    g0025(.A(G77), .ZN(new_n226));
  INV_X1    g0026(.A(G244), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(G58), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n205), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT1), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  INV_X1    g0034(.A(G20), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g0036(.A1(G58), .A2(G68), .ZN(new_n237));
  INV_X1    g0037(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n238), .A2(G50), .ZN(new_n239));
  INV_X1    g0039(.A(new_n239), .ZN(new_n240));
  AOI211_X1 g0040(.A(new_n212), .B(new_n233), .C1(new_n236), .C2(new_n240), .ZN(G361));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G264), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n243), .B(G270), .Z(new_n244));
  XNOR2_X1  g0044(.A(G238), .B(G244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G226), .B(G232), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n244), .B(new_n249), .ZN(G358));
  XOR2_X1   g0050(.A(G68), .B(G77), .Z(new_n251));
  XNOR2_X1  g0051(.A(G50), .B(G58), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(G107), .B(G116), .Z(new_n254));
  XNOR2_X1  g0054(.A(G87), .B(G97), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n253), .B(new_n256), .ZN(G351));
  OAI21_X1  g0057(.A(G20), .B1(new_n238), .B2(G50), .ZN(new_n258));
  INV_X1    g0058(.A(G150), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT8), .B(G58), .ZN(new_n265));
  OAI221_X1 g0065(.A(new_n258), .B1(new_n259), .B2(new_n261), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(new_n234), .ZN(new_n268));
  INV_X1    g0068(.A(G1), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G13), .A3(G20), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n266), .A2(new_n268), .B1(new_n224), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n268), .B1(new_n269), .B2(G20), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n272), .B1(new_n224), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n275), .B(KEYINPUT9), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT3), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n262), .ZN(new_n278));
  NAND2_X1  g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G222), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G223), .A2(G1698), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n280), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G1), .A3(G13), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n284), .B(new_n287), .C1(G77), .C2(new_n280), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n269), .B1(G41), .B2(G45), .ZN(new_n289));
  INV_X1    g0089(.A(G274), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n286), .A2(new_n289), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n288), .B(new_n292), .C1(new_n225), .C2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(G200), .B2(new_n294), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n276), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(KEYINPUT10), .B1(new_n297), .B2(KEYINPUT69), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n299), .ZN(new_n301));
  INV_X1    g0101(.A(G169), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n294), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n275), .B(new_n303), .C1(G179), .C2(new_n294), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n300), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT13), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n280), .A2(G226), .A3(new_n281), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n280), .A2(G232), .A3(G1698), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT70), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT70), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n280), .A2(new_n311), .A3(G232), .A4(G1698), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n308), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G33), .A2(G97), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n291), .B1(new_n315), .B2(new_n287), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n293), .A2(new_n214), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n306), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n286), .B1(new_n313), .B2(new_n314), .ZN(new_n320));
  NOR4_X1   g0120(.A1(new_n320), .A2(KEYINPUT13), .A3(new_n317), .A4(new_n291), .ZN(new_n321));
  OAI21_X1  g0121(.A(G200), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n260), .A2(G50), .B1(G20), .B2(new_n213), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(new_n264), .B2(new_n226), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n268), .ZN(new_n325));
  XOR2_X1   g0125(.A(KEYINPUT71), .B(KEYINPUT11), .Z(new_n326));
  XNOR2_X1  g0126(.A(new_n325), .B(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n274), .A2(new_n213), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n271), .A2(new_n213), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT12), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n329), .B(new_n330), .ZN(new_n331));
  NOR3_X1   g0131(.A1(new_n327), .A2(new_n328), .A3(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n314), .ZN(new_n333));
  AOI211_X1 g0133(.A(new_n333), .B(new_n308), .C1(new_n312), .C2(new_n310), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n318), .B(new_n292), .C1(new_n334), .C2(new_n286), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT13), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n316), .A2(new_n306), .A3(new_n318), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(new_n337), .A3(G190), .ZN(new_n338));
  AND3_X1   g0138(.A1(new_n322), .A2(new_n332), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(G169), .B1(new_n319), .B2(new_n321), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT14), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n336), .A2(new_n337), .A3(G179), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT14), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n343), .B(G169), .C1(new_n319), .C2(new_n321), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n341), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n332), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n339), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AND2_X1   g0147(.A1(KEYINPUT3), .A2(G33), .ZN(new_n348));
  NOR2_X1   g0148(.A1(KEYINPUT3), .A2(G33), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT7), .B1(new_n350), .B2(new_n235), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT7), .ZN(new_n352));
  NOR4_X1   g0152(.A1(new_n348), .A2(new_n349), .A3(new_n352), .A4(G20), .ZN(new_n353));
  OAI21_X1  g0153(.A(G68), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n229), .A2(new_n213), .ZN(new_n355));
  OAI21_X1  g0155(.A(G20), .B1(new_n355), .B2(new_n237), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n260), .A2(G159), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n354), .A2(KEYINPUT16), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT72), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n354), .A2(new_n359), .ZN(new_n362));
  XOR2_X1   g0162(.A(KEYINPUT73), .B(KEYINPUT16), .Z(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT72), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n354), .A2(new_n365), .A3(KEYINPUT16), .A4(new_n359), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n361), .A2(new_n268), .A3(new_n364), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n265), .A2(new_n270), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n273), .B2(new_n265), .ZN(new_n369));
  OR2_X1    g0169(.A1(G223), .A2(G1698), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n225), .A2(G1698), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n370), .B(new_n371), .C1(new_n348), .C2(new_n349), .ZN(new_n372));
  NAND2_X1  g0172(.A1(G33), .A2(G87), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n286), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n286), .A2(G232), .A3(new_n289), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NOR3_X1   g0176(.A1(new_n374), .A2(new_n291), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n295), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(G200), .B2(new_n377), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n367), .A2(new_n369), .A3(new_n379), .ZN(new_n380));
  XNOR2_X1  g0180(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT75), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n384), .A2(KEYINPUT17), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n367), .A2(new_n369), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n372), .A2(new_n373), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n291), .B1(new_n389), .B2(new_n287), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n302), .B1(new_n390), .B2(new_n375), .ZN(new_n391));
  INV_X1    g0191(.A(G179), .ZN(new_n392));
  NOR4_X1   g0192(.A1(new_n374), .A2(new_n376), .A3(new_n392), .A4(new_n291), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT74), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n390), .A2(G179), .A3(new_n375), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT74), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n395), .B(new_n396), .C1(new_n377), .C2(new_n302), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n388), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT18), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n388), .A2(KEYINPUT18), .A3(new_n398), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n383), .A2(new_n387), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G20), .A2(G77), .ZN(new_n404));
  XNOR2_X1  g0204(.A(KEYINPUT15), .B(G87), .ZN(new_n405));
  OAI221_X1 g0205(.A(new_n404), .B1(new_n265), .B2(new_n261), .C1(new_n264), .C2(new_n405), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n406), .A2(new_n268), .B1(new_n226), .B2(new_n271), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n273), .A2(G77), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G238), .A2(G1698), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n280), .B(new_n411), .C1(new_n230), .C2(G1698), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n412), .B(new_n287), .C1(G107), .C2(new_n280), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n413), .B(new_n292), .C1(new_n227), .C2(new_n293), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G200), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n410), .B(new_n415), .C1(new_n295), .C2(new_n414), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n302), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n417), .B(new_n409), .C1(G179), .C2(new_n414), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  XOR2_X1   g0219(.A(new_n419), .B(KEYINPUT68), .Z(new_n420));
  NAND4_X1  g0220(.A1(new_n305), .A2(new_n347), .A3(new_n403), .A4(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(G41), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n269), .B(G45), .C1(new_n422), .C2(KEYINPUT5), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT5), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(G41), .ZN(new_n425));
  OAI211_X1 g0225(.A(G264), .B(new_n286), .C1(new_n423), .C2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n217), .A2(new_n281), .ZN(new_n428));
  OAI221_X1 g0228(.A(new_n428), .B1(G257), .B2(new_n281), .C1(new_n348), .C2(new_n349), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G33), .A2(G294), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n286), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n427), .B1(new_n431), .B2(KEYINPUT87), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT77), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n290), .B1(new_n425), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n423), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n422), .A2(KEYINPUT5), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT77), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n434), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n432), .B(new_n438), .C1(KEYINPUT87), .C2(new_n431), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n278), .A2(new_n279), .B1(new_n219), .B2(G1698), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n440), .A2(new_n428), .B1(G33), .B2(G294), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n438), .B(new_n426), .C1(new_n441), .C2(new_n286), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  OAI22_X1  g0243(.A1(new_n439), .A2(G190), .B1(new_n443), .B2(G200), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n269), .A2(G33), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n270), .A2(new_n445), .A3(new_n234), .A4(new_n267), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G107), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n270), .A2(G107), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n449), .B(KEYINPUT25), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n235), .A2(G107), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n451), .B(KEYINPUT23), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n263), .A2(G116), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n280), .A2(new_n235), .A3(G87), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT22), .ZN(new_n455));
  OR2_X1    g0255(.A1(new_n455), .A2(KEYINPUT86), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n452), .B(new_n453), .C1(new_n454), .C2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n455), .A2(KEYINPUT86), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n454), .A2(new_n459), .A3(new_n456), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n458), .A2(KEYINPUT24), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT24), .ZN(new_n462));
  INV_X1    g0262(.A(new_n460), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(new_n457), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n461), .A2(new_n268), .A3(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n444), .A2(new_n448), .A3(new_n450), .A4(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n465), .A2(new_n448), .A3(new_n450), .ZN(new_n467));
  INV_X1    g0267(.A(new_n432), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n438), .B1(new_n431), .B2(KEYINPUT87), .ZN(new_n469));
  OAI21_X1  g0269(.A(G169), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n443), .A2(KEYINPUT88), .A3(G179), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT88), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(new_n442), .B2(new_n392), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n467), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n466), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(G244), .B1(new_n348), .B2(new_n349), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT4), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n477), .A2(new_n478), .B1(G33), .B2(G283), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n280), .A2(KEYINPUT4), .A3(G244), .A4(new_n281), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n478), .B1(new_n280), .B2(G250), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n479), .B(new_n480), .C1(new_n281), .C2(new_n481), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n482), .A2(new_n287), .ZN(new_n483));
  OAI211_X1 g0283(.A(G257), .B(new_n286), .C1(new_n423), .C2(new_n425), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n438), .A2(KEYINPUT78), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT78), .B1(new_n438), .B2(new_n484), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(G169), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n438), .A2(new_n484), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT78), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n438), .A2(KEYINPUT78), .A3(new_n484), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n482), .A2(new_n287), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n493), .A2(new_n494), .A3(G179), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n488), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT80), .ZN(new_n497));
  OAI21_X1  g0297(.A(G107), .B1(new_n351), .B2(new_n353), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT76), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(G107), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n501), .A2(KEYINPUT6), .A3(G97), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n218), .A2(new_n501), .ZN(new_n503));
  NOR2_X1   g0303(.A1(G97), .A2(G107), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n502), .B1(new_n505), .B2(KEYINPUT6), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n506), .A2(G20), .B1(G77), .B2(new_n260), .ZN(new_n507));
  OAI211_X1 g0307(.A(KEYINPUT76), .B(G107), .C1(new_n351), .C2(new_n353), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n500), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n268), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n271), .A2(new_n218), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n446), .B2(new_n218), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n497), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  AOI211_X1 g0314(.A(KEYINPUT80), .B(new_n512), .C1(new_n509), .C2(new_n268), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n496), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n512), .B1(new_n509), .B2(new_n268), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n491), .A2(new_n492), .B1(new_n482), .B2(new_n287), .ZN(new_n518));
  NAND2_X1  g0318(.A1(KEYINPUT79), .A2(G200), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n518), .A2(new_n295), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT79), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n518), .B1(new_n521), .B2(G200), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n517), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n235), .B(G68), .C1(new_n348), .C2(new_n349), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT81), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n280), .A2(KEYINPUT81), .A3(new_n235), .A4(G68), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT19), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n235), .B1(new_n314), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n504), .A2(new_n216), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n235), .A2(G33), .A3(G97), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n529), .A2(new_n530), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n526), .A2(new_n527), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n268), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n405), .A2(new_n271), .ZN(new_n535));
  INV_X1    g0335(.A(new_n405), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n447), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n534), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n227), .A2(G1698), .ZN(new_n539));
  OAI221_X1 g0339(.A(new_n539), .B1(G238), .B2(G1698), .C1(new_n348), .C2(new_n349), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G33), .A2(G116), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n286), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(G45), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n217), .B1(new_n543), .B2(G1), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n269), .A2(new_n290), .A3(G45), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n286), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n392), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n302), .B1(new_n542), .B2(new_n546), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n538), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n547), .A2(G190), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n533), .A2(new_n268), .B1(new_n271), .B2(new_n405), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n447), .A2(G87), .ZN(new_n553));
  OAI21_X1  g0353(.A(G200), .B1(new_n542), .B2(new_n546), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n551), .A2(new_n552), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n516), .A2(new_n523), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(G116), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n267), .A2(new_n234), .B1(G20), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(G20), .B1(G33), .B2(G283), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n262), .A2(G97), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n561), .A2(new_n562), .A3(KEYINPUT83), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT83), .B1(new_n561), .B2(new_n562), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n560), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT20), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(KEYINPUT20), .B(new_n560), .C1(new_n563), .C2(new_n564), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n281), .A2(G257), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G264), .A2(G1698), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n570), .B(new_n571), .C1(new_n348), .C2(new_n349), .ZN(new_n572));
  INV_X1    g0372(.A(G303), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n278), .A2(new_n573), .A3(new_n279), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n287), .A3(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(G270), .B(new_n286), .C1(new_n423), .C2(new_n425), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n438), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G200), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT82), .B1(new_n447), .B2(G116), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT82), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n446), .A2(new_n580), .A3(new_n559), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n271), .A2(new_n559), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n569), .A2(new_n578), .A3(new_n582), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT85), .ZN(new_n585));
  OR2_X1    g0385(.A1(new_n577), .A2(new_n295), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n567), .A2(new_n568), .B1(new_n559), .B2(new_n271), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT85), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n587), .A2(new_n588), .A3(new_n582), .A4(new_n578), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n585), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT84), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n577), .A2(G169), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(new_n587), .B2(new_n582), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n591), .B1(new_n593), .B2(KEYINPUT21), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n569), .A2(new_n582), .A3(new_n583), .ZN(new_n595));
  INV_X1    g0395(.A(new_n592), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT21), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(KEYINPUT84), .A3(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n592), .A2(new_n598), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n577), .A2(new_n392), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n595), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n590), .A2(new_n594), .A3(new_n599), .A4(new_n602), .ZN(new_n603));
  NOR4_X1   g0403(.A1(new_n421), .A2(new_n476), .A3(new_n558), .A4(new_n603), .ZN(G372));
  NOR2_X1   g0404(.A1(new_n391), .A2(new_n393), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT18), .B1(new_n388), .B2(new_n606), .ZN(new_n607));
  AOI211_X1 g0407(.A(new_n400), .B(new_n605), .C1(new_n367), .C2(new_n369), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n380), .A2(new_n386), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n610), .A2(new_n382), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n345), .A2(new_n346), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n611), .B1(new_n612), .B2(new_n418), .ZN(new_n613));
  INV_X1    g0413(.A(new_n339), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n609), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n300), .A2(new_n301), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n304), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT90), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n493), .A2(new_n494), .A3(G179), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n302), .B1(new_n493), .B2(new_n494), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n488), .A2(KEYINPUT90), .A3(new_n495), .ZN(new_n623));
  AOI211_X1 g0423(.A(new_n517), .B(new_n556), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT91), .B1(new_n624), .B2(KEYINPUT26), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT26), .ZN(new_n626));
  OR3_X1    g0426(.A1(new_n516), .A2(new_n626), .A3(new_n556), .ZN(new_n627));
  INV_X1    g0427(.A(new_n517), .ZN(new_n628));
  INV_X1    g0428(.A(new_n623), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT90), .B1(new_n488), .B2(new_n495), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n628), .B(new_n557), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT91), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(new_n632), .A3(new_n626), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n625), .A2(new_n627), .A3(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n516), .A2(new_n523), .A3(new_n466), .A4(new_n557), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n594), .A2(new_n599), .A3(new_n602), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n475), .ZN(new_n639));
  AOI21_X1  g0439(.A(KEYINPUT89), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n637), .B1(new_n467), .B2(new_n474), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT89), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n641), .A2(new_n635), .A3(new_n642), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n634), .B(new_n550), .C1(new_n640), .C2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n618), .B1(new_n645), .B2(new_n421), .ZN(G369));
  INV_X1    g0446(.A(KEYINPUT92), .ZN(new_n647));
  INV_X1    g0447(.A(new_n603), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n207), .A2(G20), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  OR3_X1    g0450(.A1(new_n650), .A2(KEYINPUT27), .A3(G1), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT27), .B1(new_n650), .B2(G1), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(G213), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(G343), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n595), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n647), .B1(new_n648), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n637), .A2(new_n595), .A3(new_n656), .ZN(new_n659));
  MUX2_X1   g0459(.A(new_n647), .B(new_n658), .S(new_n659), .Z(new_n660));
  INV_X1    g0460(.A(G330), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n467), .A2(new_n656), .ZN(new_n663));
  OAI22_X1  g0463(.A1(new_n476), .A2(new_n663), .B1(new_n475), .B2(new_n655), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g0465(.A(new_n655), .B(KEYINPUT93), .Z(new_n666));
  NOR2_X1   g0466(.A1(new_n475), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n638), .A2(new_n656), .ZN(new_n668));
  INV_X1    g0468(.A(new_n476), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n665), .A2(new_n670), .ZN(G399));
  AND3_X1   g0471(.A1(new_n516), .A2(new_n523), .A3(new_n557), .ZN(new_n672));
  INV_X1    g0472(.A(new_n666), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n672), .A2(new_n669), .A3(new_n648), .A4(new_n673), .ZN(new_n674));
  NOR4_X1   g0474(.A1(new_n431), .A2(new_n542), .A3(new_n427), .A4(new_n546), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n675), .A2(new_n494), .A3(new_n493), .A4(new_n601), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(KEYINPUT30), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT30), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n518), .A2(new_n678), .A3(new_n675), .A4(new_n601), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n442), .A2(new_n577), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n518), .A2(G179), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n547), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n677), .A2(new_n679), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(new_n673), .ZN(new_n684));
  XOR2_X1   g0484(.A(KEYINPUT94), .B(KEYINPUT31), .Z(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT95), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n677), .A2(new_n679), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n681), .A2(new_n682), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n656), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT31), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT95), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n684), .A2(new_n694), .A3(new_n685), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n674), .A2(new_n687), .A3(new_n693), .A4(new_n695), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n631), .A2(KEYINPUT26), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n699), .B(new_n550), .C1(new_n641), .C2(new_n635), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n516), .A2(KEYINPUT26), .A3(new_n556), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n655), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT29), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT29), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n644), .A2(new_n704), .A3(new_n673), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n698), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n269), .ZN(new_n707));
  INV_X1    g0507(.A(new_n209), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G41), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n530), .A2(G116), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(G1), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n239), .B2(new_n710), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n707), .A2(new_n714), .ZN(G364));
  NOR2_X1   g0515(.A1(G179), .A2(G200), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n235), .B1(new_n716), .B2(G190), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(KEYINPUT99), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n717), .A2(KEYINPUT99), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G200), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n235), .A2(new_n392), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n295), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OAI22_X1  g0526(.A1(new_n721), .A2(new_n218), .B1(new_n726), .B2(new_n224), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n235), .A2(G190), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n729), .A2(KEYINPUT96), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(KEYINPUT96), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n722), .A2(G179), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G107), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n235), .A2(new_n295), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n732), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n735), .B(new_n280), .C1(new_n216), .C2(new_n737), .ZN(new_n738));
  XOR2_X1   g0538(.A(new_n738), .B(KEYINPUT98), .Z(new_n739));
  NOR2_X1   g0539(.A1(new_n724), .A2(G190), .ZN(new_n740));
  AOI211_X1 g0540(.A(new_n727), .B(new_n739), .C1(G68), .C2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n392), .A2(G200), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n728), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G77), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n730), .A2(new_n731), .A3(new_n716), .ZN(new_n746));
  XNOR2_X1  g0546(.A(KEYINPUT97), .B(G159), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT32), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n736), .A2(new_n742), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G58), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n741), .A2(new_n745), .A3(new_n750), .A4(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(G294), .ZN(new_n755));
  INV_X1    g0555(.A(G311), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n721), .A2(new_n755), .B1(new_n756), .B2(new_n743), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(G326), .B2(new_n725), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n758), .B(KEYINPUT100), .Z(new_n759));
  INV_X1    g0559(.A(new_n746), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n759), .B1(G329), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n752), .A2(G322), .ZN(new_n762));
  INV_X1    g0562(.A(G317), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(KEYINPUT33), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n763), .A2(KEYINPUT33), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n740), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n734), .A2(G283), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n761), .A2(new_n762), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n350), .B1(new_n737), .B2(new_n573), .ZN(new_n769));
  XOR2_X1   g0569(.A(new_n769), .B(KEYINPUT101), .Z(new_n770));
  OAI21_X1  g0570(.A(new_n754), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n234), .B1(G20), .B2(new_n302), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G13), .A2(G33), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G20), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n660), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(G355), .A2(new_n209), .A3(new_n280), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n253), .A2(new_n543), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n708), .A2(new_n280), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(G45), .B2(new_n239), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n778), .B1(G116), .B2(new_n209), .C1(new_n779), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n776), .A2(new_n772), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n269), .B1(new_n649), .B2(G45), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n709), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n773), .A2(new_n777), .A3(new_n784), .A4(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n662), .ZN(new_n789));
  INV_X1    g0589(.A(new_n787), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n660), .A2(new_n661), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n788), .A2(new_n792), .ZN(G396));
  OAI21_X1  g0593(.A(new_n416), .B1(new_n410), .B2(new_n655), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n418), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n418), .A2(new_n656), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(new_n645), .B2(new_n666), .ZN(new_n799));
  INV_X1    g0599(.A(new_n798), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n644), .A2(new_n673), .A3(new_n800), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(new_n698), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n790), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n721), .A2(new_n218), .B1(new_n755), .B2(new_n751), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT102), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n734), .A2(G87), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n808), .B1(new_n559), .B2(new_n743), .C1(new_n756), .C2(new_n746), .ZN(new_n809));
  INV_X1    g0609(.A(new_n740), .ZN(new_n810));
  INV_X1    g0610(.A(G283), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n726), .A2(new_n573), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n350), .B1(new_n737), .B2(new_n501), .ZN(new_n814));
  NOR4_X1   g0614(.A1(new_n809), .A2(new_n812), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n740), .A2(G150), .B1(G143), .B2(new_n752), .ZN(new_n816));
  INV_X1    g0616(.A(G137), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n816), .B1(new_n817), .B2(new_n726), .C1(new_n743), .C2(new_n748), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT34), .ZN(new_n819));
  INV_X1    g0619(.A(new_n737), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n818), .A2(new_n819), .B1(G50), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n213), .B2(new_n733), .ZN(new_n822));
  INV_X1    g0622(.A(G132), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n746), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n721), .A2(new_n229), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n280), .B1(new_n818), .B2(new_n819), .ZN(new_n826));
  NOR4_X1   g0626(.A1(new_n822), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n772), .B1(new_n815), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n828), .A2(new_n787), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n772), .A2(new_n774), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n829), .B1(G77), .B2(new_n831), .C1(new_n775), .C2(new_n800), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n804), .A2(new_n832), .ZN(G384));
  NAND2_X1  g0633(.A1(new_n346), .A2(new_n656), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT104), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n347), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n345), .A2(new_n346), .A3(new_n656), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n798), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n690), .A2(KEYINPUT31), .A3(new_n656), .ZN(new_n842));
  INV_X1    g0642(.A(new_n685), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n683), .B2(new_n655), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n674), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT38), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n388), .A2(new_n654), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n383), .A2(new_n387), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n401), .A2(new_n402), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT37), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n394), .A2(new_n397), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n854), .A2(new_n653), .B1(new_n367), .B2(new_n369), .ZN(new_n855));
  INV_X1    g0655(.A(new_n380), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n853), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n367), .A2(new_n369), .B1(new_n605), .B2(new_n653), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n859), .A2(KEYINPUT37), .A3(new_n380), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n848), .B1(new_n852), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n388), .B1(new_n398), .B2(new_n654), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT37), .B1(new_n863), .B2(new_n380), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n380), .A2(KEYINPUT37), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n865), .A2(new_n858), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(KEYINPUT38), .B(new_n867), .C1(new_n403), .C2(new_n849), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n862), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n847), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n849), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n611), .B2(new_n609), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT106), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n857), .A2(new_n874), .A3(new_n860), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT106), .B1(new_n864), .B2(new_n866), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n873), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n848), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n868), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT108), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n878), .A2(KEYINPUT108), .A3(new_n868), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n841), .A2(KEYINPUT40), .A3(new_n846), .ZN(new_n884));
  OAI22_X1  g0684(.A1(new_n871), .A2(KEYINPUT40), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n846), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n421), .A2(new_n886), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n885), .B(new_n887), .Z(new_n888));
  NOR2_X1   g0688(.A1(new_n888), .A2(new_n661), .ZN(new_n889));
  INV_X1    g0689(.A(new_n840), .ZN(new_n890));
  AOI211_X1 g0690(.A(new_n837), .B(new_n339), .C1(new_n345), .C2(new_n346), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n890), .B1(new_n891), .B2(new_n836), .ZN(new_n892));
  AOI211_X1 g0692(.A(new_n870), .B(new_n892), .C1(new_n801), .C2(new_n797), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n609), .B2(new_n653), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT39), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n878), .A2(new_n895), .A3(new_n868), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT107), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n878), .A2(KEYINPUT107), .A3(new_n895), .A4(new_n868), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT105), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n869), .B2(KEYINPUT39), .ZN(new_n901));
  AOI211_X1 g0701(.A(KEYINPUT105), .B(new_n895), .C1(new_n862), .C2(new_n868), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n898), .B(new_n899), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n612), .A2(new_n656), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n894), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n421), .B1(new_n705), .B2(new_n703), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n907), .A2(new_n617), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n906), .B(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n889), .B1(new_n909), .B2(KEYINPUT109), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n909), .B(KEYINPUT109), .Z(new_n911));
  OAI221_X1 g0711(.A(new_n910), .B1(new_n269), .B2(new_n649), .C1(new_n911), .C2(new_n889), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n559), .B1(new_n506), .B2(KEYINPUT35), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n913), .B(new_n236), .C1(KEYINPUT35), .C2(new_n506), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT36), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT103), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n213), .B2(G50), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n224), .A2(KEYINPUT103), .A3(G68), .ZN(new_n918));
  OAI21_X1  g0718(.A(G77), .B1(new_n229), .B2(new_n213), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n917), .B(new_n918), .C1(new_n239), .C2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n920), .A2(G1), .A3(new_n207), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n912), .A2(new_n915), .A3(new_n921), .ZN(G367));
  INV_X1    g0722(.A(new_n721), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(G68), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n725), .A2(G143), .B1(G150), .B2(new_n752), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI221_X1 g0726(.A(new_n280), .B1(new_n224), .B2(new_n743), .C1(new_n926), .C2(KEYINPUT110), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(KEYINPUT110), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n733), .A2(new_n226), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n747), .B2(new_n740), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n928), .B(new_n930), .C1(new_n229), .C2(new_n737), .ZN(new_n931));
  XOR2_X1   g0731(.A(KEYINPUT111), .B(G137), .Z(new_n932));
  AOI211_X1 g0732(.A(new_n927), .B(new_n931), .C1(new_n760), .C2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n744), .A2(G283), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n737), .A2(new_n559), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n760), .A2(G317), .B1(new_n935), .B2(KEYINPUT46), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n734), .A2(G97), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n350), .B1(new_n810), .B2(new_n755), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(G311), .B2(new_n725), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n940), .B1(KEYINPUT46), .B2(new_n935), .C1(new_n501), .C2(new_n721), .ZN(new_n941));
  AOI211_X1 g0741(.A(new_n938), .B(new_n941), .C1(G303), .C2(new_n752), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n933), .B1(new_n934), .B2(new_n942), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT47), .Z(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n772), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n552), .A2(new_n553), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n656), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n557), .A2(new_n947), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n947), .A2(new_n550), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n948), .A2(new_n776), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n780), .ZN(new_n951));
  OAI221_X1 g0751(.A(new_n783), .B1(new_n209), .B2(new_n405), .C1(new_n244), .C2(new_n951), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n945), .A2(new_n787), .A3(new_n950), .A4(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT112), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n709), .B(KEYINPUT41), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n516), .B(new_n523), .C1(new_n673), .C2(new_n517), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n628), .B(new_n666), .C1(new_n629), .C2(new_n630), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n670), .A2(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT44), .Z(new_n960));
  NAND2_X1  g0760(.A1(new_n670), .A2(new_n958), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT45), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(new_n665), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n668), .A2(new_n669), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n664), .B2(new_n668), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n662), .B(new_n966), .Z(new_n967));
  OR2_X1    g0767(.A1(new_n967), .A2(new_n706), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n964), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n955), .B1(new_n969), .B2(new_n706), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n970), .A2(new_n785), .ZN(new_n971));
  INV_X1    g0771(.A(new_n958), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n972), .A2(new_n965), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT42), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n516), .B1(new_n972), .B2(new_n475), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n673), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n948), .A2(new_n949), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n974), .A2(new_n976), .B1(KEYINPUT43), .B2(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n977), .A2(KEYINPUT43), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n978), .B(new_n979), .Z(new_n980));
  NOR2_X1   g0780(.A1(new_n665), .A2(new_n972), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n980), .B(new_n981), .Z(new_n982));
  OAI21_X1  g0782(.A(new_n954), .B1(new_n971), .B2(new_n982), .ZN(G387));
  NOR2_X1   g0783(.A1(new_n967), .A2(new_n785), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT113), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n967), .A2(new_n706), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n968), .A2(new_n709), .A3(new_n986), .ZN(new_n987));
  NOR3_X1   g0787(.A1(new_n664), .A2(G20), .A3(new_n775), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n820), .A2(G77), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n989), .B1(new_n213), .B2(new_n743), .C1(new_n810), .C2(new_n265), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n350), .B(new_n990), .C1(G50), .C2(new_n752), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n725), .A2(KEYINPUT115), .A3(G159), .ZN(new_n992));
  AOI21_X1  g0792(.A(KEYINPUT115), .B1(new_n725), .B2(G159), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n721), .A2(new_n405), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n993), .B(new_n994), .C1(G150), .C2(new_n760), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n991), .A2(new_n937), .A3(new_n992), .A4(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n740), .A2(G311), .B1(new_n725), .B2(G322), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT116), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n573), .B2(new_n743), .C1(new_n763), .C2(new_n751), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT48), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n811), .B2(new_n721), .C1(new_n755), .C2(new_n737), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT49), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n734), .A2(G116), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n760), .A2(G326), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1003), .A2(new_n350), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n996), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n772), .ZN(new_n1009));
  NOR3_X1   g0809(.A1(new_n265), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n711), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(G68), .A2(G77), .ZN(new_n1013));
  OAI21_X1  g0813(.A(KEYINPUT50), .B1(new_n265), .B2(G50), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1012), .A2(new_n543), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n780), .B(new_n1015), .C1(new_n249), .C2(new_n543), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1011), .A2(new_n209), .A3(new_n280), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(G107), .C2(new_n209), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT114), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n783), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1009), .A2(new_n787), .A3(new_n1020), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n985), .B(new_n987), .C1(new_n988), .C2(new_n1021), .ZN(G393));
  OAI21_X1  g0822(.A(new_n783), .B1(new_n951), .B2(new_n256), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G97), .B2(new_n708), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n721), .A2(new_n226), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n350), .B1(new_n820), .B2(G68), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n807), .B(new_n1026), .C1(new_n224), .C2(new_n810), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1025), .B(new_n1027), .C1(G143), .C2(new_n760), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n265), .B2(new_n743), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n725), .A2(G150), .B1(G159), .B2(new_n752), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT117), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT51), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n743), .A2(new_n755), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n760), .A2(G322), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n735), .B(new_n1034), .C1(new_n559), .C2(new_n721), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n725), .A2(G317), .B1(G311), .B2(new_n752), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT52), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n350), .B1(new_n810), .B2(new_n573), .ZN(new_n1038));
  NOR3_X1   g0838(.A1(new_n1035), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n811), .B2(new_n737), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n1029), .A2(new_n1032), .B1(new_n1033), .B2(new_n1040), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n790), .B(new_n1024), .C1(new_n1041), .C2(new_n772), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1042), .A2(KEYINPUT118), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(KEYINPUT118), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n972), .A2(new_n776), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n710), .B1(new_n964), .B2(new_n968), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1046), .B1(new_n785), .B2(new_n964), .C1(new_n1048), .C2(new_n969), .ZN(G390));
  OAI211_X1 g0849(.A(new_n655), .B(new_n795), .C1(new_n700), .C2(new_n701), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n797), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n839), .A2(new_n840), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n904), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1053), .A2(new_n881), .A3(new_n882), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n801), .A2(new_n797), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n904), .B1(new_n1055), .B2(new_n1052), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1054), .B1(new_n1056), .B2(new_n903), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT119), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1052), .A2(G330), .A3(new_n800), .A4(new_n846), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  AND3_X1   g0860(.A1(new_n1057), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1058), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n697), .A2(new_n841), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1054), .B(new_n1064), .C1(new_n1056), .C2(new_n903), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1063), .A2(new_n786), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n772), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n810), .A2(new_n501), .B1(new_n218), .B2(new_n743), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1068), .A2(KEYINPUT124), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n746), .A2(new_n755), .ZN(new_n1070));
  OR3_X1    g0870(.A1(new_n1069), .A2(new_n1025), .A3(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1068), .A2(KEYINPUT124), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n350), .B1(new_n216), .B2(new_n737), .C1(new_n733), .C2(new_n213), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1074), .B1(new_n559), .B2(new_n751), .C1(new_n811), .C2(new_n726), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n932), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n280), .B1(new_n810), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(G159), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n721), .A2(new_n1078), .B1(new_n733), .B2(new_n224), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1077), .B(new_n1079), .C1(G125), .C2(new_n760), .ZN(new_n1080));
  XOR2_X1   g0880(.A(KEYINPUT54), .B(G143), .Z(new_n1081));
  NAND2_X1  g0881(.A1(new_n744), .A2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n737), .A2(new_n259), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT53), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n725), .A2(G128), .B1(G132), .B2(new_n752), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1080), .A2(new_n1082), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1067), .B1(new_n1075), .B2(new_n1086), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n790), .B(new_n1087), .C1(new_n265), .C2(new_n830), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n903), .B2(new_n775), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1066), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT123), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(KEYINPUT119), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1057), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n1065), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT120), .ZN(new_n1096));
  NOR4_X1   g0896(.A1(new_n558), .A2(new_n476), .A3(new_n603), .A4(new_n666), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n842), .A2(new_n844), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1096), .B(G330), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n800), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1096), .B1(new_n846), .B2(G330), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n892), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT121), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1051), .B1(new_n697), .B2(new_n841), .ZN(new_n1105));
  OAI211_X1 g0905(.A(KEYINPUT121), .B(new_n892), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1052), .B1(new_n697), .B2(new_n800), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1055), .B1(new_n1060), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n421), .A2(new_n886), .A3(new_n661), .ZN(new_n1111));
  NOR3_X1   g0911(.A1(new_n907), .A2(new_n1111), .A3(new_n617), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n1110), .A2(KEYINPUT122), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(KEYINPUT122), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1091), .B1(new_n1095), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT122), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1110), .A2(KEYINPUT122), .A3(new_n1112), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1063), .A2(new_n1121), .A3(KEYINPUT123), .A4(new_n1065), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1116), .A2(new_n1122), .B1(new_n1095), .B2(new_n1115), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1090), .B1(new_n1123), .B2(new_n709), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(G378));
  NAND2_X1  g0925(.A1(new_n1116), .A2(new_n1122), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n1112), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n305), .B(new_n1128), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n275), .A2(new_n654), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1129), .B(new_n1130), .ZN(new_n1131));
  OR3_X1    g0931(.A1(new_n885), .A2(new_n661), .A3(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1131), .B1(new_n885), .B2(new_n661), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n906), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1132), .A2(new_n905), .A3(new_n894), .A4(new_n1133), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1127), .A2(KEYINPUT57), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT57), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1112), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n1116), .B2(new_n1122), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1140), .B1(new_n1142), .B2(new_n1137), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1139), .A2(new_n709), .A3(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1135), .A2(new_n786), .A3(new_n1136), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n787), .B1(G50), .B2(new_n831), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n751), .A2(new_n501), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n923), .A2(G68), .B1(new_n536), .B2(new_n744), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n1148), .B1(new_n229), .B2(new_n733), .C1(new_n218), .C2(new_n810), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1147), .B(new_n1149), .C1(G116), .C2(new_n725), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n760), .A2(G283), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n280), .A2(G41), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1150), .A2(new_n989), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT58), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n224), .B1(new_n348), .B2(G41), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n923), .A2(G150), .B1(G137), .B2(new_n744), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n820), .A2(new_n1081), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n740), .A2(G132), .B1(G128), .B2(new_n752), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(G125), .B2(new_n725), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT59), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(G33), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1163));
  AOI21_X1  g0963(.A(G41), .B1(new_n760), .B2(G124), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1163), .B(new_n1164), .C1(new_n748), .C2(new_n733), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1154), .B(new_n1155), .C1(new_n1162), .C2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1146), .B1(new_n1166), .B2(new_n772), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n1131), .B2(new_n775), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT125), .Z(new_n1169));
  AND2_X1   g0969(.A1(new_n1145), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1144), .A2(new_n1170), .ZN(G375));
  NAND3_X1  g0971(.A1(new_n1141), .A2(new_n1109), .A3(new_n1107), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1119), .A2(new_n1120), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n955), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n892), .A2(new_n774), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n929), .B(new_n994), .C1(G294), .C2(new_n725), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n751), .A2(new_n811), .B1(new_n743), .B2(new_n501), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n280), .B(new_n1177), .C1(new_n760), .C2(G303), .ZN(new_n1178));
  AND2_X1   g0978(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n218), .B2(new_n737), .C1(new_n559), .C2(new_n810), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n280), .B1(new_n726), .B2(new_n823), .C1(new_n733), .C2(new_n229), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G50), .B2(new_n923), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n744), .A2(G150), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n740), .A2(new_n1081), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n1076), .A2(new_n751), .B1(new_n1078), .B2(new_n737), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n760), .B2(G128), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .A4(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1067), .B1(new_n1180), .B2(new_n1187), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n790), .B(new_n1188), .C1(new_n213), .C2(new_n830), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1110), .A2(new_n786), .B1(new_n1175), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1174), .A2(new_n1190), .ZN(G381));
  NAND3_X1  g0991(.A1(new_n1144), .A2(new_n1124), .A3(new_n1170), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(G384), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(G381), .A2(G396), .A3(G393), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(G387), .A2(G390), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .A4(new_n1196), .ZN(G407));
  OAI211_X1 g0997(.A(G407), .B(G213), .C1(G343), .C2(new_n1192), .ZN(G409));
  XNOR2_X1  g0998(.A(G387), .B(G390), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(G393), .B(G396), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1199), .B(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(G375), .A2(G378), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1127), .A2(new_n955), .A3(new_n1138), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1145), .A2(KEYINPUT126), .A3(new_n1168), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1145), .A2(new_n1168), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT126), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1204), .A2(new_n1124), .A3(new_n1205), .A4(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(G343), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(G213), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT60), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1172), .A2(new_n1213), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n709), .B(new_n1214), .C1(new_n1173), .C2(new_n1213), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1215), .A2(G384), .A3(new_n1190), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(G384), .B1(new_n1215), .B2(new_n1190), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1203), .A2(new_n1212), .A3(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1202), .B1(new_n1221), .B2(KEYINPUT63), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1218), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1210), .A2(G213), .A3(G2897), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1223), .A2(new_n1216), .A3(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1224), .B1(new_n1223), .B2(new_n1216), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1124), .B1(new_n1144), .B2(new_n1170), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1227), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(KEYINPUT63), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT61), .B1(new_n1231), .B2(new_n1220), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1222), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1220), .A2(KEYINPUT62), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT62), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1203), .A2(new_n1212), .A3(new_n1235), .A4(new_n1219), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT61), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1230), .A2(KEYINPUT127), .A3(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT127), .B1(new_n1230), .B2(new_n1238), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1237), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1233), .B1(new_n1241), .B2(new_n1201), .ZN(G405));
  NAND3_X1  g1042(.A1(new_n1202), .A2(new_n1192), .A3(new_n1203), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1201), .B1(new_n1193), .B2(new_n1228), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(new_n1219), .ZN(G402));
endmodule


