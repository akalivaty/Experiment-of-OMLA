//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n819, new_n821,
    new_n822, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942;
  INV_X1    g000(.A(G36gat), .ZN(new_n202));
  AND2_X1   g001(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n206), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n210));
  XNOR2_X1  g009(.A(G43gat), .B(G50gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n210), .A2(new_n211), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT17), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT93), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT93), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n212), .A2(new_n213), .A3(new_n217), .A4(KEYINPUT17), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G15gat), .B(G22gat), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n220), .A2(G1gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT92), .ZN(new_n222));
  AOI21_X1  g021(.A(G8gat), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n220), .B1(new_n224), .B2(G1gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n223), .A2(new_n226), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n214), .A2(new_n215), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n219), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n214), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n227), .A2(new_n228), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n230), .A2(new_n231), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT18), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n234), .B1(new_n219), .B2(new_n229), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(KEYINPUT18), .A3(new_n231), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n233), .B(new_n232), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n231), .B(KEYINPUT13), .Z(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n238), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G113gat), .B(G141gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(G197gat), .ZN(new_n246));
  XOR2_X1   g045(.A(KEYINPUT11), .B(G169gat), .Z(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT12), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n244), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n238), .A2(new_n249), .A3(new_n240), .A4(new_n243), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(KEYINPUT94), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT94), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n244), .A2(new_n254), .A3(new_n250), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G15gat), .B(G43gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(G71gat), .B(G99gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n261));
  OAI221_X1 g060(.A(new_n260), .B1(G183gat), .B2(G190gat), .C1(new_n261), .C2(KEYINPUT65), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n262), .B1(KEYINPUT65), .B2(new_n261), .ZN(new_n263));
  INV_X1    g062(.A(G169gat), .ZN(new_n264));
  INV_X1    g063(.A(G176gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT23), .ZN(new_n267));
  NAND2_X1  g066(.A1(G169gat), .A2(G176gat), .ZN(new_n268));
  OR2_X1    g067(.A1(new_n268), .A2(KEYINPUT66), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(KEYINPUT66), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n263), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n260), .B1(G183gat), .B2(G190gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n274), .A2(new_n261), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n267), .A2(KEYINPUT25), .A3(new_n271), .ZN(new_n276));
  OAI22_X1  g075(.A1(new_n273), .A2(KEYINPUT25), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G183gat), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT67), .B1(new_n278), .B2(KEYINPUT27), .ZN(new_n279));
  AOI21_X1  g078(.A(G190gat), .B1(new_n278), .B2(KEYINPUT27), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT27), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(new_n282), .A3(G183gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n279), .A2(new_n280), .A3(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT28), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n287), .B1(new_n282), .B2(G183gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(new_n280), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT69), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT69), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n286), .A2(new_n292), .A3(new_n289), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n264), .A2(new_n265), .A3(KEYINPUT70), .ZN(new_n295));
  AOI22_X1  g094(.A1(new_n269), .A2(new_n270), .B1(KEYINPUT26), .B2(new_n295), .ZN(new_n296));
  OR2_X1    g095(.A1(new_n295), .A2(KEYINPUT26), .ZN(new_n297));
  AOI22_X1  g096(.A1(new_n296), .A2(new_n297), .B1(G183gat), .B2(G190gat), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT71), .B1(new_n294), .B2(new_n298), .ZN(new_n299));
  AOI221_X4 g098(.A(KEYINPUT69), .B1(new_n280), .B2(new_n288), .C1(new_n284), .C2(new_n285), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n292), .B1(new_n286), .B2(new_n289), .ZN(new_n301));
  OAI211_X1 g100(.A(KEYINPUT71), .B(new_n298), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n277), .B1(new_n299), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT73), .ZN(new_n305));
  INV_X1    g104(.A(G113gat), .ZN(new_n306));
  INV_X1    g105(.A(G120gat), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT1), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(new_n306), .B2(new_n307), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n310));
  INV_X1    g109(.A(G127gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n310), .B1(new_n311), .B2(G134gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G127gat), .B(G134gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n313), .B(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n304), .A2(new_n305), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G227gat), .A2(G233gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n318), .B(KEYINPUT64), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT71), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(new_n302), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n313), .B(new_n314), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT73), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n316), .A2(new_n305), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n323), .A2(new_n277), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n317), .A2(new_n319), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT33), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n259), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(KEYINPUT74), .A3(KEYINPUT32), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n328), .A2(KEYINPUT32), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OR2_X1    g134(.A1(new_n259), .A2(new_n329), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n328), .A2(KEYINPUT32), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n328), .A2(KEYINPUT75), .A3(KEYINPUT32), .A4(new_n336), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n332), .A2(new_n335), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n317), .A2(new_n327), .ZN(new_n342));
  INV_X1    g141(.A(new_n319), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n344), .A2(KEYINPUT34), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(KEYINPUT34), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT76), .B1(new_n341), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G78gat), .B(G106gat), .ZN(new_n349));
  INV_X1    g148(.A(G50gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(G228gat), .A2(G233gat), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G155gat), .ZN(new_n354));
  INV_X1    g153(.A(G162gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n354), .A2(new_n355), .A3(KEYINPUT79), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n357), .B1(G155gat), .B2(G162gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n356), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(G148gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(G141gat), .ZN(new_n362));
  INV_X1    g161(.A(G141gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(G148gat), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT2), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  OR2_X1    g164(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n354), .A2(new_n355), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n359), .B1(new_n367), .B2(KEYINPUT2), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n362), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n364), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n362), .A2(new_n369), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n368), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n366), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT29), .ZN(new_n376));
  XOR2_X1   g175(.A(G211gat), .B(G218gat), .Z(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT77), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT22), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n379), .A2(new_n380), .B1(G211gat), .B2(G218gat), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n381), .B1(new_n379), .B2(new_n380), .ZN(new_n382));
  XNOR2_X1  g181(.A(G197gat), .B(G204gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n378), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n378), .B1(new_n382), .B2(new_n383), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n376), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n375), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n382), .A2(new_n383), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n377), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n384), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n366), .A2(new_n373), .A3(new_n388), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n392), .B1(new_n376), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n353), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n366), .A2(new_n373), .A3(KEYINPUT81), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT81), .B1(new_n366), .B2(new_n373), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT29), .B1(new_n391), .B2(new_n384), .ZN(new_n399));
  OAI22_X1  g198(.A1(new_n397), .A2(new_n398), .B1(new_n399), .B2(KEYINPUT3), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n393), .A2(new_n376), .ZN(new_n401));
  INV_X1    g200(.A(new_n392), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n400), .A2(new_n403), .A3(new_n352), .ZN(new_n404));
  INV_X1    g203(.A(G22gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n395), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT87), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n405), .B1(new_n395), .B2(new_n404), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n351), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT86), .B(KEYINPUT31), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n404), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(G22gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n351), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n413), .A2(new_n407), .A3(new_n414), .A4(new_n406), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n410), .A2(new_n411), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n411), .B1(new_n410), .B2(new_n415), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(new_n341), .B2(new_n347), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n335), .A2(new_n331), .A3(new_n330), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n339), .A2(new_n340), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n347), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT76), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n348), .A2(new_n419), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT91), .ZN(new_n427));
  INV_X1    g226(.A(G226gat), .ZN(new_n428));
  INV_X1    g227(.A(G233gat), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n304), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  AND2_X1   g229(.A1(new_n277), .A2(new_n320), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n376), .B1(new_n428), .B2(new_n429), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n392), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n431), .A2(G226gat), .A3(G233gat), .ZN(new_n435));
  INV_X1    g234(.A(new_n304), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n435), .B(new_n402), .C1(new_n436), .C2(new_n432), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(G8gat), .B(G36gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(G64gat), .B(G92gat), .ZN(new_n440));
  XOR2_X1   g239(.A(new_n439), .B(new_n440), .Z(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n434), .A2(KEYINPUT30), .A3(new_n437), .A4(new_n441), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n434), .A2(new_n437), .A3(new_n441), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT78), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT30), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n434), .A2(KEYINPUT78), .A3(new_n437), .A4(new_n441), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n445), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n316), .A2(new_n375), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n453), .A2(KEYINPUT4), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT81), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n374), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n456), .A2(new_n316), .A3(new_n396), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT4), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n454), .B1(new_n458), .B2(KEYINPUT82), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT82), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n457), .A2(new_n460), .A3(KEYINPUT4), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n374), .A2(KEYINPUT3), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n463), .A2(new_n324), .A3(new_n393), .ZN(new_n464));
  NAND2_X1  g263(.A1(G225gat), .A2(G233gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n462), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT5), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n324), .A2(new_n374), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n465), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT83), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT83), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n471), .A2(new_n475), .A3(new_n472), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n469), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n468), .A2(KEYINPUT84), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT84), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n466), .B1(new_n459), .B2(new_n461), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n475), .B1(new_n471), .B2(new_n472), .ZN(new_n481));
  AOI211_X1 g280(.A(KEYINPUT83), .B(new_n465), .C1(new_n453), .C2(new_n470), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT5), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n479), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n466), .A2(KEYINPUT5), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n453), .A2(KEYINPUT4), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(KEYINPUT4), .B2(new_n457), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G1gat), .B(G29gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(KEYINPUT0), .ZN(new_n492));
  XNOR2_X1  g291(.A(G57gat), .B(G85gat), .ZN(new_n493));
  XOR2_X1   g292(.A(new_n492), .B(new_n493), .Z(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT85), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n478), .A2(new_n484), .B1(new_n488), .B2(new_n486), .ZN(new_n498));
  OR3_X1    g297(.A1(new_n498), .A2(KEYINPUT85), .A3(new_n494), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT6), .B1(new_n498), .B2(new_n494), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n498), .A2(new_n494), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT6), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n452), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT91), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n348), .A2(new_n419), .A3(new_n505), .A4(new_n425), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n427), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT35), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n500), .A2(new_n496), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT90), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n510), .A3(new_n503), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n502), .A2(KEYINPUT90), .A3(KEYINPUT6), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n452), .A2(KEYINPUT35), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n422), .A2(new_n423), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n419), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n508), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n418), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n465), .B1(new_n488), .B2(new_n464), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n522), .B(KEYINPUT39), .C1(new_n472), .C2(new_n471), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n523), .B(new_n494), .C1(KEYINPUT39), .C2(new_n522), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(KEYINPUT40), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n525), .A2(new_n496), .A3(new_n452), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n448), .A2(new_n450), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n438), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT37), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT89), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n531), .A2(new_n441), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT38), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n529), .A2(KEYINPUT89), .A3(new_n530), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n402), .B1(new_n430), .B2(new_n433), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n435), .B(new_n392), .C1(new_n436), .C2(new_n432), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n535), .A2(KEYINPUT37), .A3(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT88), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n532), .A2(new_n533), .A3(new_n534), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n438), .A2(KEYINPUT37), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n532), .A2(new_n534), .A3(new_n540), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n528), .B(new_n539), .C1(new_n541), .C2(new_n533), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n511), .A2(new_n512), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n520), .B(new_n526), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n341), .A2(new_n347), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n515), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT36), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n348), .A2(KEYINPUT36), .A3(new_n545), .A4(new_n425), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n504), .A2(new_n520), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n544), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n256), .B1(new_n519), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G57gat), .B(G64gat), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G71gat), .B(G78gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(KEYINPUT95), .B(KEYINPUT21), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G231gat), .A2(G233gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G127gat), .B(G155gat), .Z(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT20), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n563), .B(new_n565), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n227), .A2(new_n228), .B1(KEYINPUT21), .B2(new_n558), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT97), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n566), .B(new_n568), .Z(new_n569));
  XNOR2_X1  g368(.A(G183gat), .B(G211gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n570), .B(new_n571), .Z(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n569), .B(new_n573), .ZN(new_n574));
  AND2_X1   g373(.A1(G232gat), .A2(G233gat), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(KEYINPUT41), .ZN(new_n576));
  XNOR2_X1  g375(.A(G134gat), .B(G162gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(G99gat), .B(G106gat), .Z(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G85gat), .A2(G92gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT98), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT7), .ZN(new_n584));
  NAND2_X1  g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  INV_X1    g384(.A(G85gat), .ZN(new_n586));
  INV_X1    g385(.A(G92gat), .ZN(new_n587));
  AOI22_X1  g386(.A1(KEYINPUT8), .A2(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT99), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n581), .B1(new_n584), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n584), .A2(new_n581), .A3(new_n589), .ZN(new_n592));
  AOI22_X1  g391(.A1(new_n591), .A2(new_n592), .B1(new_n214), .B2(new_n215), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n219), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G190gat), .B(G218gat), .Z(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n592), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n597), .A2(new_n590), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n598), .A2(new_n214), .B1(KEYINPUT41), .B2(new_n575), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n594), .A2(new_n596), .A3(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n596), .B1(new_n594), .B2(new_n599), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n579), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n594), .A2(new_n599), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n595), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n605), .A2(new_n578), .A3(new_n600), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n574), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n559), .B1(new_n597), .B2(new_n590), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n591), .A2(new_n558), .A3(new_n592), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT10), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n598), .A2(KEYINPUT10), .A3(new_n558), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G230gat), .A2(G233gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n609), .A2(new_n610), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n617), .A2(G230gat), .A3(G233gat), .ZN(new_n618));
  XOR2_X1   g417(.A(G120gat), .B(G148gat), .Z(new_n619));
  XNOR2_X1  g418(.A(G176gat), .B(G204gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n616), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n615), .B(KEYINPUT100), .Z(new_n623));
  AOI21_X1  g422(.A(new_n623), .B1(new_n612), .B2(new_n613), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n621), .B1(new_n625), .B2(new_n618), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n608), .A2(new_n627), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n501), .A2(KEYINPUT101), .A3(new_n503), .ZN(new_n629));
  AOI21_X1  g428(.A(KEYINPUT101), .B1(new_n501), .B2(new_n503), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n553), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g432(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n634));
  NAND3_X1  g433(.A1(new_n553), .A2(new_n452), .A3(new_n628), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT16), .B(G8gat), .Z(new_n636));
  XOR2_X1   g435(.A(new_n636), .B(KEYINPUT103), .Z(new_n637));
  OAI21_X1  g436(.A(new_n634), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n635), .A2(G8gat), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n636), .A2(KEYINPUT42), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n638), .B(new_n639), .C1(new_n635), .C2(new_n640), .ZN(G1325gat));
  NAND2_X1  g440(.A1(new_n553), .A2(new_n628), .ZN(new_n642));
  OAI21_X1  g441(.A(G15gat), .B1(new_n642), .B2(new_n550), .ZN(new_n643));
  INV_X1    g442(.A(new_n628), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n644), .A2(new_n546), .A3(G15gat), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n553), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n643), .A2(new_n646), .ZN(G1326gat));
  NOR2_X1   g446(.A1(new_n642), .A2(new_n520), .ZN(new_n648));
  XOR2_X1   g447(.A(KEYINPUT43), .B(G22gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(G1327gat));
  NAND2_X1  g449(.A1(new_n519), .A2(new_n552), .ZN(new_n651));
  INV_X1    g450(.A(new_n607), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(KEYINPUT44), .ZN(new_n654));
  AOI21_X1  g453(.A(KEYINPUT105), .B1(new_n508), .B2(new_n518), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT105), .ZN(new_n656));
  AOI211_X1 g455(.A(new_n656), .B(new_n517), .C1(new_n507), .C2(KEYINPUT35), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n552), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  AND3_X1   g457(.A1(new_n603), .A2(new_n606), .A3(KEYINPUT106), .ZN(new_n659));
  AOI21_X1  g458(.A(KEYINPUT106), .B1(new_n603), .B2(new_n606), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(KEYINPUT44), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n658), .A2(KEYINPUT107), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(KEYINPUT107), .B1(new_n658), .B2(new_n662), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n654), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n574), .A2(new_n256), .A3(new_n627), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n666), .B(KEYINPUT104), .Z(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n631), .ZN(new_n669));
  OAI21_X1  g468(.A(G29gat), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n651), .A2(new_n652), .A3(new_n666), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n671), .A2(G29gat), .A3(new_n669), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n672), .B(KEYINPUT45), .Z(new_n673));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n673), .ZN(G1328gat));
  INV_X1    g473(.A(new_n452), .ZN(new_n675));
  OAI21_X1  g474(.A(G36gat), .B1(new_n668), .B2(new_n675), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n671), .A2(G36gat), .A3(new_n675), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT46), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(G1329gat));
  INV_X1    g478(.A(new_n546), .ZN(new_n680));
  INV_X1    g479(.A(G43gat), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n671), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n683), .B(KEYINPUT108), .Z(new_n684));
  INV_X1    g483(.A(new_n550), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n665), .A2(new_n685), .A3(new_n667), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n684), .B1(G43gat), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n667), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT107), .ZN(new_n689));
  INV_X1    g488(.A(new_n552), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n519), .A2(new_n656), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n508), .A2(KEYINPUT105), .A3(new_n518), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n662), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n689), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n658), .A2(KEYINPUT107), .A3(new_n662), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n688), .B1(new_n697), .B2(new_n654), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n681), .B1(new_n698), .B2(new_n685), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT47), .B1(new_n671), .B2(new_n682), .ZN(new_n700));
  OAI22_X1  g499(.A1(new_n687), .A2(KEYINPUT47), .B1(new_n699), .B2(new_n700), .ZN(G1330gat));
  INV_X1    g500(.A(KEYINPUT48), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n350), .B1(new_n698), .B2(new_n418), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n671), .A2(G50gat), .A3(new_n520), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(G50gat), .B1(new_n668), .B2(new_n520), .ZN(new_n706));
  INV_X1    g505(.A(new_n704), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n706), .A2(KEYINPUT48), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n708), .ZN(G1331gat));
  INV_X1    g508(.A(new_n256), .ZN(new_n710));
  INV_X1    g509(.A(new_n627), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n608), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n658), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n631), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g515(.A(new_n452), .B(KEYINPUT109), .ZN(new_n717));
  AOI211_X1 g516(.A(new_n717), .B(new_n713), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n718));
  NOR2_X1   g517(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT110), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT111), .Z(new_n721));
  XNOR2_X1  g520(.A(new_n718), .B(new_n721), .ZN(G1333gat));
  OAI21_X1  g521(.A(G71gat), .B1(new_n713), .B2(new_n550), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n546), .A2(G71gat), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n723), .B1(new_n713), .B2(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(G1334gat));
  NAND2_X1  g526(.A1(new_n714), .A2(new_n418), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g528(.A1(new_n574), .A2(new_n710), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(new_n711), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n665), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G85gat), .B1(new_n733), .B2(new_n669), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT51), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n731), .A2(new_n607), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n735), .B1(new_n693), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n658), .A2(KEYINPUT51), .A3(new_n736), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n631), .A2(new_n586), .A3(new_n627), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n734), .B1(new_n741), .B2(new_n742), .ZN(G1336gat));
  INV_X1    g542(.A(new_n717), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n744), .A2(new_n587), .A3(new_n627), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT114), .B1(new_n740), .B2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT114), .ZN(new_n748));
  AOI211_X1 g547(.A(new_n748), .B(new_n745), .C1(new_n738), .C2(new_n739), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n665), .A2(new_n744), .A3(new_n732), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G92gat), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n745), .B1(new_n738), .B2(new_n739), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT113), .ZN(new_n756));
  OAI21_X1  g555(.A(KEYINPUT52), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  AOI211_X1 g556(.A(KEYINPUT113), .B(new_n745), .C1(new_n738), .C2(new_n739), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(G92gat), .B1(new_n733), .B2(new_n675), .ZN(new_n760));
  AOI22_X1  g559(.A1(new_n753), .A2(new_n754), .B1(new_n759), .B2(new_n760), .ZN(G1337gat));
  OAI21_X1  g560(.A(G99gat), .B1(new_n733), .B2(new_n550), .ZN(new_n762));
  OR3_X1    g561(.A1(new_n546), .A2(G99gat), .A3(new_n711), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n741), .B2(new_n763), .ZN(G1338gat));
  INV_X1    g563(.A(G106gat), .ZN(new_n765));
  INV_X1    g564(.A(new_n732), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n766), .B1(new_n697), .B2(new_n654), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n765), .B1(new_n767), .B2(new_n418), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n520), .A2(new_n711), .A3(G106gat), .ZN(new_n769));
  INV_X1    g568(.A(new_n739), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT51), .B1(new_n658), .B2(new_n736), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT115), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT115), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n740), .A2(new_n774), .A3(new_n769), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT53), .B1(new_n768), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(G106gat), .B1(new_n733), .B2(new_n520), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n778), .A2(new_n779), .A3(new_n772), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n777), .A2(new_n780), .ZN(G1339gat));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n612), .A2(new_n613), .A3(new_n623), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n616), .A2(KEYINPUT54), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n621), .B1(new_n624), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT55), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(new_n622), .ZN(new_n788));
  OAI22_X1  g587(.A1(new_n239), .A2(new_n231), .B1(new_n241), .B2(new_n242), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n248), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n252), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n784), .A2(KEYINPUT55), .A3(new_n786), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n788), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n793), .A2(new_n661), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n253), .A2(new_n788), .A3(new_n255), .A4(new_n792), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n791), .A2(new_n627), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OR2_X1    g597(.A1(new_n659), .A2(new_n660), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n782), .B(new_n795), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n574), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n799), .B1(new_n796), .B2(new_n797), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT116), .B1(new_n802), .B2(new_n794), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n800), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n628), .A2(new_n256), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n804), .A2(KEYINPUT117), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT117), .B1(new_n804), .B2(new_n805), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n516), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n669), .A2(new_n744), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n811), .A2(new_n306), .A3(new_n256), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n427), .A2(new_n506), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n808), .A2(new_n813), .A3(new_n631), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(new_n744), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n710), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n812), .B1(new_n816), .B2(new_n306), .ZN(G1340gat));
  NOR3_X1   g616(.A1(new_n811), .A2(new_n307), .A3(new_n711), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n815), .A2(new_n627), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n818), .B1(new_n819), .B2(new_n307), .ZN(G1341gat));
  NAND3_X1  g619(.A1(new_n815), .A2(new_n311), .A3(new_n574), .ZN(new_n821));
  OAI21_X1  g620(.A(G127gat), .B1(new_n811), .B2(new_n801), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(G1342gat));
  NOR4_X1   g622(.A1(new_n814), .A2(G134gat), .A3(new_n452), .A4(new_n607), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(KEYINPUT56), .ZN(new_n825));
  OAI21_X1  g624(.A(G134gat), .B1(new_n811), .B2(new_n607), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT118), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(G1343gat));
  INV_X1    g627(.A(KEYINPUT58), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n798), .A2(new_n652), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n801), .B1(new_n830), .B2(new_n794), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n805), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n520), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n806), .A2(new_n807), .A3(new_n520), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n836), .B2(KEYINPUT57), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n810), .A2(new_n550), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n837), .A2(new_n710), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(G141gat), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n829), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n804), .A2(new_n805), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n804), .A2(KEYINPUT117), .A3(new_n805), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n418), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n833), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n838), .B1(new_n849), .B2(new_n835), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n363), .B1(new_n850), .B2(new_n710), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n808), .A2(new_n631), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n685), .A2(new_n520), .ZN(new_n853));
  XOR2_X1   g652(.A(new_n853), .B(KEYINPUT119), .Z(new_n854));
  NOR2_X1   g653(.A1(new_n256), .A2(G141gat), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NOR4_X1   g655(.A1(new_n852), .A2(new_n854), .A3(new_n744), .A4(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT121), .B1(new_n851), .B2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n859));
  INV_X1    g658(.A(new_n857), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n841), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n843), .A2(new_n858), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n843), .B1(new_n858), .B2(new_n861), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n862), .A2(new_n863), .ZN(G1344gat));
  NOR3_X1   g663(.A1(new_n852), .A2(new_n854), .A3(new_n744), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n865), .A2(new_n627), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n361), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n850), .A2(new_n867), .A3(new_n627), .ZN(new_n869));
  INV_X1    g668(.A(new_n793), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n830), .B1(new_n652), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n805), .B1(new_n871), .B2(new_n574), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT57), .B1(new_n872), .B2(new_n418), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n873), .B1(new_n808), .B2(new_n834), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n839), .A2(new_n627), .ZN(new_n875));
  OAI211_X1 g674(.A(KEYINPUT59), .B(G148gat), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n868), .A2(new_n869), .A3(new_n876), .ZN(G1345gat));
  NAND3_X1  g676(.A1(new_n865), .A2(new_n354), .A3(new_n574), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n837), .A2(new_n839), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(new_n801), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n878), .B1(new_n880), .B2(new_n354), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n881), .B(KEYINPUT122), .Z(G1346gat));
  OAI21_X1  g681(.A(G162gat), .B1(new_n879), .B2(new_n661), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n852), .A2(new_n854), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n884), .A2(new_n355), .A3(new_n675), .A4(new_n652), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(G1347gat));
  NOR2_X1   g685(.A1(new_n631), .A2(new_n675), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n808), .A2(new_n809), .A3(new_n887), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n888), .A2(new_n264), .A3(new_n256), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n806), .A2(new_n807), .A3(new_n631), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n813), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n717), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n710), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n889), .B1(new_n893), .B2(new_n264), .ZN(G1348gat));
  OAI21_X1  g693(.A(G176gat), .B1(new_n888), .B2(new_n711), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n744), .A2(new_n265), .A3(new_n627), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n891), .B2(new_n896), .ZN(G1349gat));
  NAND2_X1  g696(.A1(new_n282), .A2(G183gat), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n278), .A2(KEYINPUT27), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n892), .A2(new_n898), .A3(new_n899), .A4(new_n574), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT60), .ZN(new_n901));
  OAI21_X1  g700(.A(G183gat), .B1(new_n888), .B2(new_n801), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n903), .A2(KEYINPUT124), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n903), .A2(KEYINPUT124), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n900), .A2(new_n902), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(KEYINPUT60), .ZN(new_n908));
  AOI211_X1 g707(.A(KEYINPUT123), .B(new_n901), .C1(new_n900), .C2(new_n902), .ZN(new_n909));
  OAI22_X1  g708(.A1(new_n904), .A2(new_n905), .B1(new_n908), .B2(new_n909), .ZN(G1350gat));
  OAI21_X1  g709(.A(G190gat), .B1(new_n888), .B2(new_n607), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT61), .ZN(new_n912));
  INV_X1    g711(.A(G190gat), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n892), .A2(new_n913), .A3(new_n799), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(G1351gat));
  NAND2_X1  g714(.A1(new_n887), .A2(new_n550), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n874), .A2(new_n916), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n710), .A2(G197gat), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n853), .A2(new_n744), .ZN(new_n920));
  XOR2_X1   g719(.A(new_n920), .B(KEYINPUT125), .Z(new_n921));
  AND2_X1   g720(.A1(new_n921), .A2(new_n890), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n922), .A2(new_n710), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n919), .B1(new_n923), .B2(G197gat), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT126), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n924), .B(new_n925), .ZN(G1352gat));
  NAND2_X1  g725(.A1(new_n917), .A2(new_n627), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(G204gat), .ZN(new_n928));
  INV_X1    g727(.A(G204gat), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n922), .A2(new_n929), .A3(new_n627), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n930), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT127), .B1(new_n930), .B2(KEYINPUT62), .ZN(new_n932));
  OAI221_X1 g731(.A(new_n928), .B1(KEYINPUT62), .B2(new_n930), .C1(new_n931), .C2(new_n932), .ZN(G1353gat));
  INV_X1    g732(.A(G211gat), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n922), .A2(new_n934), .A3(new_n574), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n917), .A2(new_n574), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n936), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT63), .B1(new_n936), .B2(G211gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(G1354gat));
  INV_X1    g738(.A(G218gat), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n922), .A2(new_n940), .A3(new_n799), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n874), .A2(new_n607), .A3(new_n916), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n942), .B2(new_n940), .ZN(G1355gat));
endmodule


