

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737;

  INV_X1 U365 ( .A(n640), .ZN(n346) );
  INV_X1 U366 ( .A(KEYINPUT89), .ZN(n343) );
  XNOR2_X1 U367 ( .A(n432), .B(n345), .ZN(n716) );
  XNOR2_X1 U368 ( .A(n358), .B(n434), .ZN(n724) );
  XNOR2_X1 U369 ( .A(n430), .B(n470), .ZN(n345) );
  INV_X1 U370 ( .A(G113), .ZN(n476) );
  XNOR2_X1 U371 ( .A(n344), .B(G113), .ZN(n362) );
  XNOR2_X1 U372 ( .A(n365), .B(G107), .ZN(n463) );
  INV_X2 U373 ( .A(G119), .ZN(n344) );
  XNOR2_X1 U374 ( .A(n464), .B(KEYINPUT4), .ZN(n440) );
  XNOR2_X1 U375 ( .A(n487), .B(n343), .ZN(n502) );
  XNOR2_X2 U376 ( .A(n455), .B(KEYINPUT0), .ZN(n487) );
  NAND2_X1 U377 ( .A1(n347), .A2(n346), .ZN(n641) );
  INV_X1 U378 ( .A(n690), .ZN(n347) );
  NOR2_X2 U379 ( .A1(n709), .A2(n589), .ZN(n690) );
  XNOR2_X1 U380 ( .A(G134), .B(G131), .ZN(n379) );
  INV_X1 U381 ( .A(G125), .ZN(n359) );
  NAND2_X1 U382 ( .A1(n360), .A2(n592), .ZN(n501) );
  INV_X1 U383 ( .A(G953), .ZN(n726) );
  NOR2_X2 U384 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X2 U385 ( .A1(n555), .A2(n454), .ZN(n455) );
  INV_X1 U386 ( .A(G116), .ZN(n365) );
  NOR2_X1 U387 ( .A1(n547), .A2(n607), .ZN(n534) );
  AND2_X2 U388 ( .A1(n361), .A2(n540), .ZN(n495) );
  OR2_X2 U389 ( .A1(n690), .A2(n689), .ZN(n691) );
  OR2_X2 U390 ( .A1(n690), .A2(n424), .ZN(n652) );
  NOR2_X1 U391 ( .A1(n692), .A2(n690), .ZN(n703) );
  INV_X1 U392 ( .A(G146), .ZN(n385) );
  XNOR2_X1 U393 ( .A(n387), .B(G110), .ZN(n372) );
  XNOR2_X1 U394 ( .A(G140), .B(G107), .ZN(n387) );
  XNOR2_X1 U395 ( .A(G104), .B(KEYINPUT77), .ZN(n371) );
  XNOR2_X1 U396 ( .A(n357), .B(KEYINPUT28), .ZN(n356) );
  NOR2_X1 U397 ( .A1(n566), .A2(n542), .ZN(n357) );
  XNOR2_X1 U398 ( .A(n543), .B(n395), .ZN(n491) );
  XNOR2_X1 U399 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U400 ( .A(n460), .B(n373), .ZN(n461) );
  XNOR2_X1 U401 ( .A(n468), .B(n467), .ZN(n469) );
  NOR2_X1 U402 ( .A1(G902), .A2(n700), .ZN(n468) );
  INV_X1 U403 ( .A(KEYINPUT47), .ZN(n350) );
  INV_X1 U404 ( .A(G902), .ZN(n443) );
  XNOR2_X1 U405 ( .A(n463), .B(n364), .ZN(n429) );
  INV_X1 U406 ( .A(KEYINPUT16), .ZN(n364) );
  XOR2_X1 U407 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n459) );
  XNOR2_X1 U408 ( .A(n473), .B(n375), .ZN(n474) );
  XNOR2_X1 U409 ( .A(G143), .B(G131), .ZN(n471) );
  AND2_X1 U410 ( .A1(n629), .A2(n587), .ZN(n363) );
  INV_X1 U411 ( .A(KEYINPUT102), .ZN(n485) );
  XNOR2_X1 U412 ( .A(n423), .B(n422), .ZN(n654) );
  XOR2_X1 U413 ( .A(KEYINPUT5), .B(G116), .Z(n419) );
  XOR2_X1 U414 ( .A(G110), .B(G119), .Z(n403) );
  XNOR2_X1 U415 ( .A(n352), .B(n351), .ZN(n358) );
  INV_X1 U416 ( .A(G140), .ZN(n351) );
  XNOR2_X1 U417 ( .A(KEYINPUT69), .B(KEYINPUT10), .ZN(n352) );
  XNOR2_X1 U418 ( .A(n372), .B(n371), .ZN(n389) );
  XNOR2_X1 U419 ( .A(n716), .B(n441), .ZN(n644) );
  XNOR2_X1 U420 ( .A(n354), .B(n353), .ZN(n557) );
  INV_X1 U421 ( .A(KEYINPUT107), .ZN(n353) );
  INV_X1 U422 ( .A(KEYINPUT33), .ZN(n367) );
  XNOR2_X1 U423 ( .A(n462), .B(n461), .ZN(n466) );
  AND2_X1 U424 ( .A1(n647), .A2(G953), .ZN(n708) );
  XNOR2_X1 U425 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n535) );
  NOR2_X1 U426 ( .A1(n594), .A2(n377), .ZN(n681) );
  AND2_X1 U427 ( .A1(n560), .A2(n675), .ZN(n674) );
  XNOR2_X1 U428 ( .A(KEYINPUT100), .B(n508), .ZN(n568) );
  AND2_X1 U429 ( .A1(n583), .A2(n363), .ZN(n348) );
  NOR2_X1 U430 ( .A1(n635), .A2(n631), .ZN(n349) );
  XNOR2_X1 U431 ( .A(n415), .B(n414), .ZN(n540) );
  INV_X1 U432 ( .A(n540), .ZN(n360) );
  NOR2_X2 U433 ( .A1(n621), .A2(n502), .ZN(n456) );
  NOR2_X1 U434 ( .A1(n634), .A2(n633), .ZN(n638) );
  OR2_X1 U435 ( .A1(n560), .A2(n350), .ZN(n558) );
  NAND2_X1 U436 ( .A1(n356), .A2(n355), .ZN(n354) );
  INV_X1 U437 ( .A(n543), .ZN(n355) );
  XNOR2_X2 U438 ( .A(n359), .B(G146), .ZN(n434) );
  AND2_X1 U439 ( .A1(n540), .A2(n526), .ZN(n593) );
  AND2_X1 U440 ( .A1(n567), .A2(n360), .ZN(n513) );
  AND2_X1 U441 ( .A1(n361), .A2(n514), .ZN(n660) );
  XNOR2_X1 U442 ( .A(n490), .B(n489), .ZN(n361) );
  XNOR2_X2 U443 ( .A(n420), .B(n362), .ZN(n430) );
  AND2_X1 U444 ( .A1(n583), .A2(n629), .ZN(n632) );
  NOR2_X2 U445 ( .A1(n366), .A2(G902), .ZN(n392) );
  XNOR2_X1 U446 ( .A(n366), .B(KEYINPUT57), .ZN(n684) );
  XNOR2_X2 U447 ( .A(n390), .B(n423), .ZN(n366) );
  XNOR2_X2 U448 ( .A(n368), .B(n367), .ZN(n621) );
  NAND2_X1 U449 ( .A1(n370), .A2(n369), .ZN(n368) );
  INV_X1 U450 ( .A(n567), .ZN(n369) );
  XNOR2_X1 U451 ( .A(n498), .B(KEYINPUT103), .ZN(n370) );
  XNOR2_X2 U452 ( .A(n571), .B(KEYINPUT19), .ZN(n555) );
  BUF_X1 U453 ( .A(n491), .Z(n594) );
  XOR2_X2 U454 ( .A(G478), .B(n469), .Z(n509) );
  XNOR2_X2 U455 ( .A(n484), .B(KEYINPUT35), .ZN(n733) );
  XNOR2_X1 U456 ( .A(KEYINPUT96), .B(KEYINPUT97), .ZN(n373) );
  AND2_X1 U457 ( .A1(G221), .A2(n457), .ZN(n374) );
  AND2_X1 U458 ( .A1(G214), .A2(n472), .ZN(n375) );
  OR2_X1 U459 ( .A1(n540), .A2(n528), .ZN(n376) );
  XOR2_X1 U460 ( .A(KEYINPUT36), .B(n572), .Z(n377) );
  OR2_X1 U461 ( .A1(n623), .A2(n622), .ZN(n378) );
  XNOR2_X1 U462 ( .A(n477), .B(n476), .ZN(n478) );
  INV_X1 U463 ( .A(KEYINPUT74), .ZN(n416) );
  INV_X1 U464 ( .A(KEYINPUT66), .ZN(n393) );
  XNOR2_X1 U465 ( .A(n421), .B(n430), .ZN(n422) );
  XNOR2_X1 U466 ( .A(n480), .B(G475), .ZN(n481) );
  XNOR2_X1 U467 ( .A(n482), .B(n481), .ZN(n507) );
  XNOR2_X1 U468 ( .A(n536), .B(n535), .ZN(n734) );
  XNOR2_X1 U469 ( .A(n627), .B(n626), .ZN(G75) );
  XOR2_X1 U470 ( .A(n379), .B(G137), .Z(n382) );
  INV_X1 U471 ( .A(n382), .ZN(n381) );
  XNOR2_X2 U472 ( .A(G143), .B(G128), .ZN(n464) );
  INV_X1 U473 ( .A(n440), .ZN(n380) );
  NAND2_X1 U474 ( .A1(n381), .A2(n380), .ZN(n384) );
  NAND2_X1 U475 ( .A1(n382), .A2(n440), .ZN(n383) );
  NAND2_X1 U476 ( .A1(n384), .A2(n383), .ZN(n723) );
  XNOR2_X1 U477 ( .A(KEYINPUT68), .B(G101), .ZN(n433) );
  XNOR2_X1 U478 ( .A(n433), .B(n385), .ZN(n386) );
  XNOR2_X2 U479 ( .A(n723), .B(n386), .ZN(n423) );
  NAND2_X1 U480 ( .A1(G227), .A2(n726), .ZN(n388) );
  XNOR2_X1 U481 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U482 ( .A(KEYINPUT70), .B(G469), .ZN(n391) );
  XNOR2_X2 U483 ( .A(n392), .B(n391), .ZN(n543) );
  INV_X1 U484 ( .A(KEYINPUT1), .ZN(n394) );
  XNOR2_X2 U485 ( .A(KEYINPUT15), .B(G902), .ZN(n635) );
  NAND2_X1 U486 ( .A1(G234), .A2(n635), .ZN(n396) );
  XNOR2_X1 U487 ( .A(KEYINPUT20), .B(n396), .ZN(n410) );
  NAND2_X1 U488 ( .A1(n410), .A2(G221), .ZN(n400) );
  XOR2_X1 U489 ( .A(KEYINPUT92), .B(KEYINPUT21), .Z(n398) );
  INV_X1 U490 ( .A(KEYINPUT91), .ZN(n397) );
  XNOR2_X1 U491 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U492 ( .A(n400), .B(n399), .ZN(n592) );
  NAND2_X1 U493 ( .A1(G234), .A2(n726), .ZN(n401) );
  XOR2_X1 U494 ( .A(KEYINPUT8), .B(n401), .Z(n457) );
  XNOR2_X1 U495 ( .A(n724), .B(n374), .ZN(n409) );
  XNOR2_X1 U496 ( .A(G128), .B(G137), .ZN(n402) );
  XNOR2_X1 U497 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U498 ( .A(KEYINPUT24), .B(KEYINPUT71), .Z(n405) );
  XNOR2_X1 U499 ( .A(KEYINPUT23), .B(KEYINPUT76), .ZN(n404) );
  XNOR2_X1 U500 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U501 ( .A(n407), .B(n406), .Z(n408) );
  XNOR2_X1 U502 ( .A(n409), .B(n408), .ZN(n704) );
  NOR2_X1 U503 ( .A1(G902), .A2(n704), .ZN(n415) );
  XOR2_X1 U504 ( .A(KEYINPUT25), .B(KEYINPUT75), .Z(n412) );
  NAND2_X1 U505 ( .A1(n410), .A2(G217), .ZN(n411) );
  XNOR2_X1 U506 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U507 ( .A(KEYINPUT90), .B(n413), .Z(n414) );
  NOR2_X2 U508 ( .A1(n491), .A2(n501), .ZN(n417) );
  XNOR2_X2 U509 ( .A(n417), .B(n416), .ZN(n498) );
  NOR2_X1 U510 ( .A1(G953), .A2(G237), .ZN(n472) );
  NAND2_X1 U511 ( .A1(n472), .A2(G210), .ZN(n418) );
  XNOR2_X1 U512 ( .A(n419), .B(n418), .ZN(n421) );
  XNOR2_X1 U513 ( .A(KEYINPUT3), .B(KEYINPUT85), .ZN(n420) );
  NAND2_X1 U514 ( .A1(n654), .A2(n443), .ZN(n425) );
  INV_X1 U515 ( .A(G472), .ZN(n424) );
  XNOR2_X2 U516 ( .A(n425), .B(n424), .ZN(n542) );
  XNOR2_X1 U517 ( .A(KEYINPUT101), .B(KEYINPUT6), .ZN(n426) );
  XNOR2_X1 U518 ( .A(n542), .B(n426), .ZN(n567) );
  INV_X1 U519 ( .A(KEYINPUT72), .ZN(n427) );
  XNOR2_X1 U520 ( .A(n427), .B(G110), .ZN(n428) );
  XNOR2_X1 U521 ( .A(n429), .B(n428), .ZN(n432) );
  XOR2_X1 U522 ( .A(G104), .B(G122), .Z(n470) );
  XNOR2_X1 U523 ( .A(n434), .B(n433), .ZN(n438) );
  XNOR2_X1 U524 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n436) );
  NAND2_X1 U525 ( .A1(n726), .A2(G224), .ZN(n435) );
  XNOR2_X1 U526 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U527 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U528 ( .A(n440), .B(n439), .ZN(n441) );
  NAND2_X1 U529 ( .A1(n644), .A2(n635), .ZN(n446) );
  INV_X1 U530 ( .A(G237), .ZN(n442) );
  NAND2_X1 U531 ( .A1(n443), .A2(n442), .ZN(n447) );
  NAND2_X1 U532 ( .A1(n447), .A2(G210), .ZN(n444) );
  XNOR2_X1 U533 ( .A(n444), .B(KEYINPUT78), .ZN(n445) );
  XNOR2_X2 U534 ( .A(n446), .B(n445), .ZN(n581) );
  NAND2_X1 U535 ( .A1(n447), .A2(G214), .ZN(n448) );
  XNOR2_X1 U536 ( .A(n448), .B(KEYINPUT86), .ZN(n579) );
  INV_X1 U537 ( .A(n579), .ZN(n610) );
  OR2_X2 U538 ( .A1(n581), .A2(n610), .ZN(n571) );
  NAND2_X1 U539 ( .A1(G234), .A2(G237), .ZN(n449) );
  XNOR2_X1 U540 ( .A(n449), .B(KEYINPUT14), .ZN(n451) );
  NAND2_X1 U541 ( .A1(G952), .A2(n451), .ZN(n450) );
  XOR2_X1 U542 ( .A(KEYINPUT87), .B(n450), .Z(n620) );
  NOR2_X1 U543 ( .A1(n620), .A2(G953), .ZN(n525) );
  INV_X1 U544 ( .A(n525), .ZN(n453) );
  NAND2_X1 U545 ( .A1(G902), .A2(n451), .ZN(n521) );
  XOR2_X1 U546 ( .A(G898), .B(KEYINPUT88), .Z(n713) );
  NAND2_X1 U547 ( .A1(G953), .A2(n713), .ZN(n717) );
  OR2_X1 U548 ( .A1(n521), .A2(n717), .ZN(n452) );
  NAND2_X1 U549 ( .A1(n453), .A2(n452), .ZN(n454) );
  XNOR2_X1 U550 ( .A(n456), .B(KEYINPUT34), .ZN(n483) );
  NAND2_X1 U551 ( .A1(G217), .A2(n457), .ZN(n462) );
  XNOR2_X1 U552 ( .A(G134), .B(G122), .ZN(n458) );
  XNOR2_X1 U553 ( .A(n459), .B(n458), .ZN(n460) );
  XOR2_X1 U554 ( .A(n464), .B(n463), .Z(n465) );
  XNOR2_X1 U555 ( .A(n466), .B(n465), .ZN(n700) );
  XNOR2_X1 U556 ( .A(KEYINPUT99), .B(KEYINPUT98), .ZN(n467) );
  XNOR2_X1 U557 ( .A(n471), .B(n470), .ZN(n473) );
  XNOR2_X1 U558 ( .A(n724), .B(n474), .ZN(n479) );
  XOR2_X1 U559 ( .A(KEYINPUT94), .B(KEYINPUT11), .Z(n475) );
  XNOR2_X1 U560 ( .A(KEYINPUT12), .B(n475), .ZN(n477) );
  XNOR2_X1 U561 ( .A(n479), .B(n478), .ZN(n693) );
  NOR2_X1 U562 ( .A1(G902), .A2(n693), .ZN(n482) );
  XNOR2_X1 U563 ( .A(KEYINPUT95), .B(KEYINPUT13), .ZN(n480) );
  NOR2_X1 U564 ( .A1(n509), .A2(n507), .ZN(n548) );
  NAND2_X1 U565 ( .A1(n483), .A2(n548), .ZN(n484) );
  NAND2_X1 U566 ( .A1(n507), .A2(n509), .ZN(n486) );
  XNOR2_X2 U567 ( .A(n486), .B(n485), .ZN(n612) );
  AND2_X1 U568 ( .A1(n612), .A2(n592), .ZN(n488) );
  INV_X1 U569 ( .A(n487), .ZN(n499) );
  NAND2_X1 U570 ( .A1(n488), .A2(n499), .ZN(n490) );
  XNOR2_X1 U571 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n489) );
  NOR2_X1 U572 ( .A1(n594), .A2(n369), .ZN(n492) );
  NAND2_X1 U573 ( .A1(n495), .A2(n492), .ZN(n493) );
  XNOR2_X2 U574 ( .A(n493), .B(KEYINPUT32), .ZN(n630) );
  INV_X1 U575 ( .A(n594), .ZN(n577) );
  INV_X1 U576 ( .A(n542), .ZN(n600) );
  NOR2_X1 U577 ( .A1(n577), .A2(n600), .ZN(n494) );
  NAND2_X1 U578 ( .A1(n495), .A2(n494), .ZN(n670) );
  NAND2_X1 U579 ( .A1(n630), .A2(n670), .ZN(n496) );
  NOR2_X2 U580 ( .A1(n733), .A2(n496), .ZN(n497) );
  XNOR2_X1 U581 ( .A(n497), .B(KEYINPUT44), .ZN(n518) );
  NOR2_X1 U582 ( .A1(n498), .A2(n542), .ZN(n602) );
  NAND2_X1 U583 ( .A1(n602), .A2(n499), .ZN(n500) );
  XNOR2_X1 U584 ( .A(n500), .B(KEYINPUT31), .ZN(n679) );
  NOR2_X1 U585 ( .A1(n543), .A2(n501), .ZN(n504) );
  INV_X1 U586 ( .A(n502), .ZN(n503) );
  NAND2_X1 U587 ( .A1(n504), .A2(n503), .ZN(n505) );
  NOR2_X1 U588 ( .A1(n600), .A2(n505), .ZN(n665) );
  NOR2_X1 U589 ( .A1(n679), .A2(n665), .ZN(n506) );
  XNOR2_X1 U590 ( .A(n506), .B(KEYINPUT93), .ZN(n512) );
  INV_X1 U591 ( .A(n507), .ZN(n510) );
  NAND2_X1 U592 ( .A1(n510), .A2(n509), .ZN(n508) );
  NOR2_X1 U593 ( .A1(n510), .A2(n509), .ZN(n678) );
  INV_X1 U594 ( .A(n678), .ZN(n511) );
  NAND2_X1 U595 ( .A1(n568), .A2(n511), .ZN(n546) );
  NAND2_X1 U596 ( .A1(n512), .A2(n546), .ZN(n516) );
  AND2_X1 U597 ( .A1(n594), .A2(n513), .ZN(n514) );
  INV_X1 U598 ( .A(n660), .ZN(n515) );
  AND2_X1 U599 ( .A1(n516), .A2(n515), .ZN(n517) );
  NAND2_X1 U600 ( .A1(n518), .A2(n517), .ZN(n520) );
  XNOR2_X1 U601 ( .A(KEYINPUT81), .B(KEYINPUT45), .ZN(n519) );
  XNOR2_X2 U602 ( .A(n520), .B(n519), .ZN(n634) );
  BUF_X2 U603 ( .A(n634), .Z(n709) );
  INV_X1 U604 ( .A(n568), .ZN(n675) );
  NOR2_X1 U605 ( .A1(G900), .A2(n521), .ZN(n522) );
  NAND2_X1 U606 ( .A1(G953), .A2(n522), .ZN(n523) );
  XOR2_X1 U607 ( .A(KEYINPUT104), .B(n523), .Z(n524) );
  NOR2_X1 U608 ( .A1(n525), .A2(n524), .ZN(n527) );
  INV_X1 U609 ( .A(n592), .ZN(n526) );
  NOR2_X1 U610 ( .A1(n527), .A2(n526), .ZN(n541) );
  INV_X1 U611 ( .A(n541), .ZN(n528) );
  NOR2_X1 U612 ( .A1(n543), .A2(n376), .ZN(n532) );
  XNOR2_X1 U613 ( .A(KEYINPUT30), .B(KEYINPUT105), .ZN(n530) );
  OR2_X2 U614 ( .A1(n542), .A2(n610), .ZN(n529) );
  XNOR2_X1 U615 ( .A(n530), .B(n529), .ZN(n531) );
  NAND2_X1 U616 ( .A1(n532), .A2(n531), .ZN(n547) );
  XNOR2_X1 U617 ( .A(KEYINPUT73), .B(KEYINPUT38), .ZN(n533) );
  XNOR2_X1 U618 ( .A(n581), .B(n533), .ZN(n607) );
  XOR2_X1 U619 ( .A(n534), .B(KEYINPUT39), .Z(n584) );
  AND2_X1 U620 ( .A1(n675), .A2(n584), .ZN(n536) );
  INV_X1 U621 ( .A(n607), .ZN(n611) );
  AND2_X1 U622 ( .A1(n579), .A2(n611), .ZN(n537) );
  NAND2_X1 U623 ( .A1(n612), .A2(n537), .ZN(n539) );
  INV_X1 U624 ( .A(KEYINPUT41), .ZN(n538) );
  XNOR2_X2 U625 ( .A(n539), .B(n538), .ZN(n591) );
  NAND2_X1 U626 ( .A1(n541), .A2(n540), .ZN(n566) );
  NOR2_X1 U627 ( .A1(n591), .A2(n557), .ZN(n544) );
  XNOR2_X1 U628 ( .A(KEYINPUT42), .B(n544), .ZN(n737) );
  NOR2_X1 U629 ( .A1(n734), .A2(n737), .ZN(n545) );
  XNOR2_X1 U630 ( .A(n545), .B(KEYINPUT46), .ZN(n565) );
  INV_X1 U631 ( .A(n546), .ZN(n606) );
  NAND2_X1 U632 ( .A1(n606), .A2(KEYINPUT47), .ZN(n553) );
  INV_X1 U633 ( .A(n547), .ZN(n551) );
  INV_X1 U634 ( .A(n548), .ZN(n549) );
  NOR2_X1 U635 ( .A1(n581), .A2(n549), .ZN(n550) );
  NAND2_X1 U636 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U637 ( .A(KEYINPUT106), .B(n552), .ZN(n736) );
  NAND2_X1 U638 ( .A1(n553), .A2(n736), .ZN(n554) );
  XOR2_X1 U639 ( .A(KEYINPUT80), .B(n554), .Z(n559) );
  INV_X1 U640 ( .A(n555), .ZN(n556) );
  NOR2_X1 U641 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U642 ( .A1(n559), .A2(n558), .ZN(n563) );
  AND2_X1 U643 ( .A1(n560), .A2(n678), .ZN(n671) );
  NOR2_X1 U644 ( .A1(n671), .A2(n674), .ZN(n561) );
  NOR2_X1 U645 ( .A1(KEYINPUT47), .A2(n561), .ZN(n562) );
  NOR2_X1 U646 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U647 ( .A1(n565), .A2(n564), .ZN(n574) );
  INV_X1 U648 ( .A(n566), .ZN(n570) );
  NOR2_X1 U649 ( .A1(n568), .A2(n567), .ZN(n569) );
  NAND2_X1 U650 ( .A1(n570), .A2(n569), .ZN(n576) );
  NOR2_X1 U651 ( .A1(n576), .A2(n571), .ZN(n572) );
  XNOR2_X1 U652 ( .A(n681), .B(KEYINPUT84), .ZN(n573) );
  XNOR2_X1 U653 ( .A(n575), .B(KEYINPUT48), .ZN(n583) );
  NOR2_X1 U654 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U655 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U656 ( .A(KEYINPUT43), .B(n580), .ZN(n582) );
  NAND2_X1 U657 ( .A1(n582), .A2(n581), .ZN(n629) );
  NAND2_X1 U658 ( .A1(n584), .A2(n678), .ZN(n683) );
  NAND2_X1 U659 ( .A1(n632), .A2(n683), .ZN(n725) );
  NOR2_X1 U660 ( .A1(n709), .A2(n725), .ZN(n585) );
  NOR2_X1 U661 ( .A1(n585), .A2(KEYINPUT2), .ZN(n590) );
  NAND2_X1 U662 ( .A1(KEYINPUT2), .A2(n683), .ZN(n586) );
  XNOR2_X1 U663 ( .A(KEYINPUT79), .B(n586), .ZN(n587) );
  XNOR2_X1 U664 ( .A(n348), .B(KEYINPUT82), .ZN(n588) );
  INV_X1 U665 ( .A(n588), .ZN(n589) );
  OR2_X1 U666 ( .A1(n590), .A2(n690), .ZN(n625) );
  XNOR2_X1 U667 ( .A(KEYINPUT49), .B(n593), .ZN(n598) );
  XOR2_X1 U668 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n596) );
  NAND2_X1 U669 ( .A1(n594), .A2(n501), .ZN(n595) );
  XNOR2_X1 U670 ( .A(n596), .B(n595), .ZN(n597) );
  NAND2_X1 U671 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U672 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U673 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U674 ( .A(KEYINPUT51), .B(n603), .Z(n604) );
  NOR2_X1 U675 ( .A1(n591), .A2(n604), .ZN(n605) );
  XNOR2_X1 U676 ( .A(KEYINPUT118), .B(n605), .ZN(n617) );
  NOR2_X1 U677 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U678 ( .A1(n612), .A2(n608), .ZN(n609) );
  NOR2_X1 U679 ( .A1(n610), .A2(n609), .ZN(n614) );
  AND2_X1 U680 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U681 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U682 ( .A1(n621), .A2(n615), .ZN(n616) );
  NOR2_X1 U683 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U684 ( .A(n618), .B(KEYINPUT52), .ZN(n619) );
  NOR2_X1 U685 ( .A1(n620), .A2(n619), .ZN(n623) );
  NOR2_X1 U686 ( .A1(n591), .A2(n621), .ZN(n622) );
  NOR2_X1 U687 ( .A1(G953), .A2(n378), .ZN(n624) );
  NAND2_X1 U688 ( .A1(n625), .A2(n624), .ZN(n627) );
  XNOR2_X1 U689 ( .A(KEYINPUT53), .B(KEYINPUT119), .ZN(n626) );
  XNOR2_X1 U690 ( .A(G140), .B(KEYINPUT116), .ZN(n628) );
  XNOR2_X1 U691 ( .A(n629), .B(n628), .ZN(G42) );
  XNOR2_X1 U692 ( .A(n630), .B(G119), .ZN(G21) );
  INV_X1 U693 ( .A(n683), .ZN(n631) );
  NAND2_X1 U694 ( .A1(n349), .A2(n632), .ZN(n633) );
  INV_X1 U695 ( .A(n635), .ZN(n636) );
  AND2_X1 U696 ( .A1(n636), .A2(KEYINPUT2), .ZN(n637) );
  NOR2_X1 U697 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X2 U698 ( .A(n639), .B(KEYINPUT64), .ZN(n692) );
  INV_X1 U699 ( .A(G210), .ZN(n640) );
  OR2_X2 U700 ( .A1(n692), .A2(n641), .ZN(n646) );
  XOR2_X1 U701 ( .A(KEYINPUT120), .B(KEYINPUT54), .Z(n642) );
  XNOR2_X1 U702 ( .A(n642), .B(KEYINPUT55), .ZN(n643) );
  XNOR2_X1 U703 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U704 ( .A(n646), .B(n645), .ZN(n649) );
  INV_X1 U705 ( .A(G952), .ZN(n647) );
  INV_X1 U706 ( .A(n708), .ZN(n648) );
  NAND2_X1 U707 ( .A1(n649), .A2(n648), .ZN(n651) );
  XNOR2_X1 U708 ( .A(KEYINPUT83), .B(KEYINPUT56), .ZN(n650) );
  XNOR2_X1 U709 ( .A(n651), .B(n650), .ZN(G51) );
  NOR2_X1 U710 ( .A1(n692), .A2(n652), .ZN(n656) );
  XOR2_X1 U711 ( .A(KEYINPUT109), .B(KEYINPUT62), .Z(n653) );
  XNOR2_X1 U712 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U713 ( .A(n656), .B(n655), .ZN(n657) );
  NOR2_X2 U714 ( .A1(n657), .A2(n708), .ZN(n659) );
  INV_X1 U715 ( .A(KEYINPUT63), .ZN(n658) );
  XNOR2_X1 U716 ( .A(n659), .B(n658), .ZN(G57) );
  XOR2_X1 U717 ( .A(G101), .B(n660), .Z(G3) );
  XNOR2_X1 U718 ( .A(G104), .B(KEYINPUT110), .ZN(n662) );
  NAND2_X1 U719 ( .A1(n665), .A2(n675), .ZN(n661) );
  XNOR2_X1 U720 ( .A(n662), .B(n661), .ZN(G6) );
  XOR2_X1 U721 ( .A(KEYINPUT113), .B(KEYINPUT27), .Z(n664) );
  XNOR2_X1 U722 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n663) );
  XNOR2_X1 U723 ( .A(n664), .B(n663), .ZN(n669) );
  XNOR2_X1 U724 ( .A(G107), .B(KEYINPUT26), .ZN(n667) );
  NAND2_X1 U725 ( .A1(n678), .A2(n665), .ZN(n666) );
  XNOR2_X1 U726 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U727 ( .A(n669), .B(n668), .ZN(G9) );
  XNOR2_X1 U728 ( .A(G110), .B(n670), .ZN(G12) );
  XNOR2_X1 U729 ( .A(n671), .B(KEYINPUT29), .ZN(n672) );
  XNOR2_X1 U730 ( .A(n672), .B(KEYINPUT114), .ZN(n673) );
  XNOR2_X1 U731 ( .A(G128), .B(n673), .ZN(G30) );
  XOR2_X1 U732 ( .A(G146), .B(n674), .Z(G48) );
  XOR2_X1 U733 ( .A(G113), .B(KEYINPUT115), .Z(n677) );
  NAND2_X1 U734 ( .A1(n679), .A2(n675), .ZN(n676) );
  XNOR2_X1 U735 ( .A(n677), .B(n676), .ZN(G15) );
  NAND2_X1 U736 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U737 ( .A(n680), .B(G116), .ZN(G18) );
  XNOR2_X1 U738 ( .A(G125), .B(n681), .ZN(n682) );
  XNOR2_X1 U739 ( .A(n682), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U740 ( .A(G134), .B(n683), .ZN(G36) );
  NAND2_X1 U741 ( .A1(n703), .A2(G469), .ZN(n687) );
  XNOR2_X1 U742 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n685) );
  XNOR2_X1 U743 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U744 ( .A(n687), .B(n686), .ZN(n688) );
  NOR2_X1 U745 ( .A1(n708), .A2(n688), .ZN(G54) );
  INV_X1 U746 ( .A(G475), .ZN(n689) );
  NOR2_X1 U747 ( .A1(n692), .A2(n691), .ZN(n697) );
  XOR2_X1 U748 ( .A(KEYINPUT67), .B(KEYINPUT59), .Z(n695) );
  XNOR2_X1 U749 ( .A(n693), .B(KEYINPUT122), .ZN(n694) );
  XNOR2_X1 U750 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U751 ( .A(n697), .B(n696), .ZN(n698) );
  NOR2_X2 U752 ( .A1(n698), .A2(n708), .ZN(n699) );
  XNOR2_X1 U753 ( .A(n699), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U754 ( .A1(n703), .A2(G478), .ZN(n701) );
  XNOR2_X1 U755 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U756 ( .A1(n708), .A2(n702), .ZN(G63) );
  NAND2_X1 U757 ( .A1(n703), .A2(G217), .ZN(n706) );
  XOR2_X1 U758 ( .A(n704), .B(KEYINPUT123), .Z(n705) );
  XNOR2_X1 U759 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U760 ( .A1(n708), .A2(n707), .ZN(G66) );
  NOR2_X1 U761 ( .A1(n709), .A2(G953), .ZN(n715) );
  XOR2_X1 U762 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n711) );
  NAND2_X1 U763 ( .A1(G224), .A2(G953), .ZN(n710) );
  XNOR2_X1 U764 ( .A(n711), .B(n710), .ZN(n712) );
  NOR2_X1 U765 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U766 ( .A1(n715), .A2(n714), .ZN(n722) );
  XOR2_X1 U767 ( .A(KEYINPUT126), .B(KEYINPUT125), .Z(n720) );
  XOR2_X1 U768 ( .A(n716), .B(G101), .Z(n718) );
  NAND2_X1 U769 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U770 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U771 ( .A(n722), .B(n721), .ZN(G69) );
  XOR2_X1 U772 ( .A(n724), .B(n723), .Z(n728) );
  XNOR2_X1 U773 ( .A(n725), .B(n728), .ZN(n727) );
  NAND2_X1 U774 ( .A1(n727), .A2(n726), .ZN(n732) );
  XNOR2_X1 U775 ( .A(G227), .B(n728), .ZN(n729) );
  NAND2_X1 U776 ( .A1(n729), .A2(G900), .ZN(n730) );
  NAND2_X1 U777 ( .A1(n730), .A2(G953), .ZN(n731) );
  NAND2_X1 U778 ( .A1(n732), .A2(n731), .ZN(G72) );
  XOR2_X1 U779 ( .A(G122), .B(n733), .Z(G24) );
  XNOR2_X1 U780 ( .A(n734), .B(G131), .ZN(n735) );
  XNOR2_X1 U781 ( .A(n735), .B(KEYINPUT127), .ZN(G33) );
  XNOR2_X1 U782 ( .A(G143), .B(n736), .ZN(G45) );
  XOR2_X1 U783 ( .A(n737), .B(G137), .Z(G39) );
endmodule

