

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U549 ( .A(KEYINPUT99), .B(n748), .Z(n513) );
  NOR2_X2 U550 ( .A1(G2104), .A2(n520), .ZN(n867) );
  XNOR2_X2 U551 ( .A(n534), .B(n533), .ZN(n635) );
  XNOR2_X1 U552 ( .A(n745), .B(KEYINPUT98), .ZN(n807) );
  NAND2_X1 U553 ( .A1(G8), .A2(n728), .ZN(n811) );
  AND2_X1 U554 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U555 ( .A1(n754), .A2(n753), .ZN(n791) );
  AND2_X1 U556 ( .A1(G114), .A2(n866), .ZN(n514) );
  AND2_X1 U557 ( .A1(G102), .A2(n871), .ZN(n515) );
  INV_X1 U558 ( .A(n728), .ZN(n707) );
  INV_X1 U559 ( .A(KEYINPUT28), .ZN(n701) );
  XNOR2_X1 U560 ( .A(n716), .B(KEYINPUT96), .ZN(n717) );
  XNOR2_X1 U561 ( .A(n718), .B(n717), .ZN(n719) );
  INV_X1 U562 ( .A(KEYINPUT31), .ZN(n723) );
  NOR2_X1 U563 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U564 ( .A1(n758), .A2(n756), .ZN(n728) );
  INV_X1 U565 ( .A(KEYINPUT13), .ZN(n537) );
  OR2_X1 U566 ( .A1(n676), .A2(n675), .ZN(n758) );
  XOR2_X1 U567 ( .A(G543), .B(KEYINPUT0), .Z(n613) );
  NOR2_X1 U568 ( .A1(n515), .A2(n514), .ZN(n550) );
  NAND2_X1 U569 ( .A1(n551), .A2(n550), .ZN(n673) );
  AND2_X1 U570 ( .A1(G452), .A2(G94), .ZN(G173) );
  NOR2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n516) );
  XOR2_X2 U572 ( .A(KEYINPUT17), .B(n516), .Z(n870) );
  NAND2_X1 U573 ( .A1(G135), .A2(n870), .ZN(n517) );
  XNOR2_X1 U574 ( .A(n517), .B(KEYINPUT78), .ZN(n525) );
  INV_X1 U575 ( .A(G2105), .ZN(n520) );
  AND2_X1 U576 ( .A1(n520), .A2(G2104), .ZN(n871) );
  NAND2_X1 U577 ( .A1(G99), .A2(n871), .ZN(n519) );
  AND2_X1 U578 ( .A1(G2104), .A2(G2105), .ZN(n866) );
  NAND2_X1 U579 ( .A1(G111), .A2(n866), .ZN(n518) );
  NAND2_X1 U580 ( .A1(n519), .A2(n518), .ZN(n523) );
  NAND2_X1 U581 ( .A1(n867), .A2(G123), .ZN(n521) );
  XOR2_X1 U582 ( .A(KEYINPUT18), .B(n521), .Z(n522) );
  NOR2_X1 U583 ( .A1(n523), .A2(n522), .ZN(n524) );
  NAND2_X1 U584 ( .A1(n525), .A2(n524), .ZN(n926) );
  XNOR2_X1 U585 ( .A(G2096), .B(n926), .ZN(n526) );
  OR2_X1 U586 ( .A1(G2100), .A2(n526), .ZN(G156) );
  INV_X1 U587 ( .A(G651), .ZN(n532) );
  NOR2_X1 U588 ( .A1(G543), .A2(n532), .ZN(n528) );
  XNOR2_X1 U589 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n527) );
  XNOR2_X1 U590 ( .A(n528), .B(n527), .ZN(n639) );
  NAND2_X1 U591 ( .A1(n639), .A2(G56), .ZN(n529) );
  XOR2_X1 U592 ( .A(KEYINPUT14), .B(n529), .Z(n540) );
  NOR2_X2 U593 ( .A1(G651), .A2(G543), .ZN(n631) );
  NAND2_X1 U594 ( .A1(G81), .A2(n631), .ZN(n530) );
  XOR2_X1 U595 ( .A(KEYINPUT12), .B(n530), .Z(n531) );
  XNOR2_X1 U596 ( .A(n531), .B(KEYINPUT73), .ZN(n536) );
  INV_X1 U597 ( .A(KEYINPUT65), .ZN(n534) );
  NOR2_X1 U598 ( .A1(n532), .A2(n613), .ZN(n533) );
  NAND2_X1 U599 ( .A1(G68), .A2(n635), .ZN(n535) );
  NAND2_X1 U600 ( .A1(n536), .A2(n535), .ZN(n538) );
  XNOR2_X1 U601 ( .A(n538), .B(n537), .ZN(n539) );
  NOR2_X1 U602 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U603 ( .A(n541), .B(KEYINPUT74), .ZN(n544) );
  NOR2_X1 U604 ( .A1(G651), .A2(n613), .ZN(n586) );
  BUF_X1 U605 ( .A(n586), .Z(n632) );
  NAND2_X1 U606 ( .A1(n632), .A2(G43), .ZN(n542) );
  XOR2_X1 U607 ( .A(KEYINPUT75), .B(n542), .Z(n543) );
  NAND2_X1 U608 ( .A1(n544), .A2(n543), .ZN(n685) );
  INV_X1 U609 ( .A(G860), .ZN(n595) );
  OR2_X1 U610 ( .A1(n685), .A2(n595), .ZN(G153) );
  INV_X1 U611 ( .A(G132), .ZN(G219) );
  NAND2_X1 U612 ( .A1(n870), .A2(G137), .ZN(n547) );
  NAND2_X1 U613 ( .A1(G101), .A2(n871), .ZN(n545) );
  XOR2_X1 U614 ( .A(KEYINPUT23), .B(n545), .Z(n546) );
  NAND2_X1 U615 ( .A1(n547), .A2(n546), .ZN(n680) );
  NAND2_X1 U616 ( .A1(G113), .A2(n866), .ZN(n549) );
  NAND2_X1 U617 ( .A1(G125), .A2(n867), .ZN(n548) );
  NAND2_X1 U618 ( .A1(n549), .A2(n548), .ZN(n678) );
  NOR2_X1 U619 ( .A1(n680), .A2(n678), .ZN(G160) );
  AND2_X1 U620 ( .A1(n870), .A2(G138), .ZN(n552) );
  NAND2_X1 U621 ( .A1(G126), .A2(n867), .ZN(n551) );
  NOR2_X1 U622 ( .A1(n552), .A2(n673), .ZN(G164) );
  NAND2_X1 U623 ( .A1(G51), .A2(n632), .ZN(n554) );
  NAND2_X1 U624 ( .A1(G63), .A2(n639), .ZN(n553) );
  NAND2_X1 U625 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U626 ( .A(KEYINPUT6), .B(n555), .ZN(n561) );
  NAND2_X1 U627 ( .A1(n631), .A2(G89), .ZN(n556) );
  XNOR2_X1 U628 ( .A(n556), .B(KEYINPUT4), .ZN(n558) );
  NAND2_X1 U629 ( .A1(G76), .A2(n635), .ZN(n557) );
  NAND2_X1 U630 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U631 ( .A(n559), .B(KEYINPUT5), .Z(n560) );
  NOR2_X1 U632 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U633 ( .A(KEYINPUT77), .B(n562), .Z(n563) );
  XOR2_X1 U634 ( .A(KEYINPUT7), .B(n563), .Z(G168) );
  XOR2_X1 U635 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U636 ( .A1(G7), .A2(G661), .ZN(n564) );
  XNOR2_X1 U637 ( .A(n564), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U638 ( .A(G223), .ZN(n821) );
  NAND2_X1 U639 ( .A1(n821), .A2(G567), .ZN(n565) );
  XOR2_X1 U640 ( .A(KEYINPUT11), .B(n565), .Z(G234) );
  NAND2_X1 U641 ( .A1(G52), .A2(n632), .ZN(n567) );
  NAND2_X1 U642 ( .A1(G64), .A2(n639), .ZN(n566) );
  NAND2_X1 U643 ( .A1(n567), .A2(n566), .ZN(n572) );
  NAND2_X1 U644 ( .A1(G90), .A2(n631), .ZN(n569) );
  NAND2_X1 U645 ( .A1(G77), .A2(n635), .ZN(n568) );
  NAND2_X1 U646 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U647 ( .A(KEYINPUT9), .B(n570), .Z(n571) );
  NOR2_X1 U648 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U649 ( .A(KEYINPUT68), .B(n573), .ZN(G171) );
  INV_X1 U650 ( .A(G171), .ZN(G301) );
  NAND2_X1 U651 ( .A1(G301), .A2(G868), .ZN(n583) );
  NAND2_X1 U652 ( .A1(n639), .A2(G66), .ZN(n580) );
  NAND2_X1 U653 ( .A1(G92), .A2(n631), .ZN(n575) );
  NAND2_X1 U654 ( .A1(G79), .A2(n635), .ZN(n574) );
  NAND2_X1 U655 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U656 ( .A1(n632), .A2(G54), .ZN(n576) );
  XOR2_X1 U657 ( .A(KEYINPUT76), .B(n576), .Z(n577) );
  NOR2_X1 U658 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U659 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U660 ( .A(KEYINPUT15), .B(n581), .Z(n691) );
  INV_X1 U661 ( .A(n691), .ZN(n601) );
  INV_X1 U662 ( .A(n601), .ZN(n967) );
  INV_X1 U663 ( .A(G868), .ZN(n653) );
  NAND2_X1 U664 ( .A1(n967), .A2(n653), .ZN(n582) );
  NAND2_X1 U665 ( .A1(n583), .A2(n582), .ZN(G284) );
  NAND2_X1 U666 ( .A1(G91), .A2(n631), .ZN(n585) );
  NAND2_X1 U667 ( .A1(G65), .A2(n639), .ZN(n584) );
  NAND2_X1 U668 ( .A1(n585), .A2(n584), .ZN(n589) );
  NAND2_X1 U669 ( .A1(G53), .A2(n586), .ZN(n587) );
  XNOR2_X1 U670 ( .A(KEYINPUT69), .B(n587), .ZN(n588) );
  NOR2_X1 U671 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U672 ( .A1(G78), .A2(n635), .ZN(n590) );
  NAND2_X1 U673 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U674 ( .A(n592), .B(KEYINPUT70), .ZN(G299) );
  NOR2_X1 U675 ( .A1(G286), .A2(n653), .ZN(n594) );
  NOR2_X1 U676 ( .A1(G299), .A2(G868), .ZN(n593) );
  NOR2_X1 U677 ( .A1(n594), .A2(n593), .ZN(G297) );
  NAND2_X1 U678 ( .A1(n595), .A2(G559), .ZN(n596) );
  NAND2_X1 U679 ( .A1(n596), .A2(n601), .ZN(n597) );
  XNOR2_X1 U680 ( .A(n597), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U681 ( .A1(G868), .A2(n685), .ZN(n600) );
  NAND2_X1 U682 ( .A1(G868), .A2(n601), .ZN(n598) );
  NOR2_X1 U683 ( .A1(G559), .A2(n598), .ZN(n599) );
  NOR2_X1 U684 ( .A1(n600), .A2(n599), .ZN(G282) );
  NAND2_X1 U685 ( .A1(n601), .A2(G559), .ZN(n650) );
  XNOR2_X1 U686 ( .A(n685), .B(n650), .ZN(n602) );
  NOR2_X1 U687 ( .A1(n602), .A2(G860), .ZN(n609) );
  NAND2_X1 U688 ( .A1(G93), .A2(n631), .ZN(n604) );
  NAND2_X1 U689 ( .A1(G80), .A2(n635), .ZN(n603) );
  NAND2_X1 U690 ( .A1(n604), .A2(n603), .ZN(n608) );
  NAND2_X1 U691 ( .A1(G55), .A2(n632), .ZN(n606) );
  NAND2_X1 U692 ( .A1(G67), .A2(n639), .ZN(n605) );
  NAND2_X1 U693 ( .A1(n606), .A2(n605), .ZN(n607) );
  OR2_X1 U694 ( .A1(n608), .A2(n607), .ZN(n652) );
  XOR2_X1 U695 ( .A(n609), .B(n652), .Z(G145) );
  NAND2_X1 U696 ( .A1(G49), .A2(n632), .ZN(n611) );
  NAND2_X1 U697 ( .A1(G74), .A2(G651), .ZN(n610) );
  NAND2_X1 U698 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U699 ( .A1(n639), .A2(n612), .ZN(n616) );
  NAND2_X1 U700 ( .A1(G87), .A2(n613), .ZN(n614) );
  XOR2_X1 U701 ( .A(KEYINPUT79), .B(n614), .Z(n615) );
  NAND2_X1 U702 ( .A1(n616), .A2(n615), .ZN(G288) );
  NAND2_X1 U703 ( .A1(G85), .A2(n631), .ZN(n618) );
  NAND2_X1 U704 ( .A1(G60), .A2(n639), .ZN(n617) );
  NAND2_X1 U705 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U706 ( .A1(G72), .A2(n635), .ZN(n619) );
  XOR2_X1 U707 ( .A(KEYINPUT66), .B(n619), .Z(n620) );
  NOR2_X1 U708 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U709 ( .A1(n632), .A2(G47), .ZN(n622) );
  NAND2_X1 U710 ( .A1(n623), .A2(n622), .ZN(G290) );
  NAND2_X1 U711 ( .A1(G88), .A2(n631), .ZN(n625) );
  NAND2_X1 U712 ( .A1(G75), .A2(n635), .ZN(n624) );
  NAND2_X1 U713 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U714 ( .A(KEYINPUT80), .B(n626), .ZN(n630) );
  NAND2_X1 U715 ( .A1(G50), .A2(n632), .ZN(n628) );
  NAND2_X1 U716 ( .A1(G62), .A2(n639), .ZN(n627) );
  NAND2_X1 U717 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U718 ( .A1(n630), .A2(n629), .ZN(G166) );
  NAND2_X1 U719 ( .A1(G86), .A2(n631), .ZN(n634) );
  NAND2_X1 U720 ( .A1(G48), .A2(n632), .ZN(n633) );
  NAND2_X1 U721 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U722 ( .A1(n635), .A2(G73), .ZN(n636) );
  XOR2_X1 U723 ( .A(KEYINPUT2), .B(n636), .Z(n637) );
  NOR2_X1 U724 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U725 ( .A1(n639), .A2(G61), .ZN(n640) );
  NAND2_X1 U726 ( .A1(n641), .A2(n640), .ZN(G305) );
  XNOR2_X1 U727 ( .A(KEYINPUT82), .B(KEYINPUT81), .ZN(n643) );
  XNOR2_X1 U728 ( .A(G288), .B(KEYINPUT19), .ZN(n642) );
  XNOR2_X1 U729 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U730 ( .A(G299), .B(n644), .ZN(n646) );
  XNOR2_X1 U731 ( .A(G290), .B(G166), .ZN(n645) );
  XNOR2_X1 U732 ( .A(n646), .B(n645), .ZN(n647) );
  XOR2_X1 U733 ( .A(n652), .B(n647), .Z(n648) );
  XNOR2_X1 U734 ( .A(n648), .B(G305), .ZN(n649) );
  XNOR2_X1 U735 ( .A(n685), .B(n649), .ZN(n885) );
  XNOR2_X1 U736 ( .A(n650), .B(n885), .ZN(n651) );
  NAND2_X1 U737 ( .A1(n651), .A2(G868), .ZN(n655) );
  NAND2_X1 U738 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U739 ( .A1(n655), .A2(n654), .ZN(G295) );
  NAND2_X1 U740 ( .A1(G2078), .A2(G2084), .ZN(n656) );
  XOR2_X1 U741 ( .A(KEYINPUT20), .B(n656), .Z(n657) );
  NAND2_X1 U742 ( .A1(G2090), .A2(n657), .ZN(n659) );
  XOR2_X1 U743 ( .A(KEYINPUT83), .B(KEYINPUT21), .Z(n658) );
  XNOR2_X1 U744 ( .A(n659), .B(n658), .ZN(n660) );
  NAND2_X1 U745 ( .A1(G2072), .A2(n660), .ZN(G158) );
  XNOR2_X1 U746 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U747 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  XNOR2_X1 U748 ( .A(KEYINPUT71), .B(G57), .ZN(G237) );
  INV_X1 U749 ( .A(G661), .ZN(n671) );
  NOR2_X1 U750 ( .A1(G220), .A2(G219), .ZN(n661) );
  XOR2_X1 U751 ( .A(KEYINPUT22), .B(n661), .Z(n662) );
  XNOR2_X1 U752 ( .A(n662), .B(KEYINPUT84), .ZN(n663) );
  NOR2_X1 U753 ( .A1(G218), .A2(n663), .ZN(n664) );
  NAND2_X1 U754 ( .A1(G96), .A2(n664), .ZN(n828) );
  NAND2_X1 U755 ( .A1(n828), .A2(G2106), .ZN(n668) );
  NAND2_X1 U756 ( .A1(G108), .A2(G120), .ZN(n665) );
  NOR2_X1 U757 ( .A1(G237), .A2(n665), .ZN(n666) );
  NAND2_X1 U758 ( .A1(G69), .A2(n666), .ZN(n827) );
  NAND2_X1 U759 ( .A1(G567), .A2(n827), .ZN(n667) );
  NAND2_X1 U760 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U761 ( .A(n669), .B(KEYINPUT85), .ZN(n884) );
  NAND2_X1 U762 ( .A1(n884), .A2(G483), .ZN(n670) );
  NOR2_X1 U763 ( .A1(n671), .A2(n670), .ZN(n825) );
  NAND2_X1 U764 ( .A1(n825), .A2(G36), .ZN(G176) );
  XOR2_X1 U765 ( .A(KEYINPUT86), .B(G166), .Z(G303) );
  INV_X1 U766 ( .A(G1384), .ZN(n674) );
  AND2_X1 U767 ( .A1(G138), .A2(n674), .ZN(n672) );
  AND2_X1 U768 ( .A1(n870), .A2(n672), .ZN(n676) );
  AND2_X1 U769 ( .A1(n674), .A2(n673), .ZN(n675) );
  INV_X1 U770 ( .A(G40), .ZN(n677) );
  OR2_X1 U771 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U772 ( .A1(n680), .A2(n679), .ZN(n756) );
  XNOR2_X1 U773 ( .A(KEYINPUT92), .B(KEYINPUT29), .ZN(n706) );
  INV_X1 U774 ( .A(G1996), .ZN(n942) );
  NOR2_X1 U775 ( .A1(n728), .A2(n942), .ZN(n681) );
  XOR2_X1 U776 ( .A(n681), .B(KEYINPUT26), .Z(n683) );
  NAND2_X1 U777 ( .A1(n728), .A2(G1341), .ZN(n682) );
  NAND2_X1 U778 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U779 ( .A1(n685), .A2(n684), .ZN(n689) );
  NAND2_X1 U780 ( .A1(G1348), .A2(n728), .ZN(n687) );
  NAND2_X1 U781 ( .A1(G2067), .A2(n707), .ZN(n686) );
  NAND2_X1 U782 ( .A1(n687), .A2(n686), .ZN(n690) );
  NOR2_X1 U783 ( .A1(n691), .A2(n690), .ZN(n688) );
  OR2_X1 U784 ( .A1(n689), .A2(n688), .ZN(n693) );
  NAND2_X1 U785 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U786 ( .A1(n693), .A2(n692), .ZN(n698) );
  NAND2_X1 U787 ( .A1(n707), .A2(G2072), .ZN(n694) );
  XNOR2_X1 U788 ( .A(n694), .B(KEYINPUT27), .ZN(n696) );
  INV_X1 U789 ( .A(G1956), .ZN(n991) );
  NOR2_X1 U790 ( .A1(n991), .A2(n707), .ZN(n695) );
  NOR2_X1 U791 ( .A1(n696), .A2(n695), .ZN(n700) );
  INV_X1 U792 ( .A(G299), .ZN(n699) );
  NAND2_X1 U793 ( .A1(n700), .A2(n699), .ZN(n697) );
  NAND2_X1 U794 ( .A1(n698), .A2(n697), .ZN(n704) );
  NOR2_X1 U795 ( .A1(n700), .A2(n699), .ZN(n702) );
  XNOR2_X1 U796 ( .A(n702), .B(n701), .ZN(n703) );
  NAND2_X1 U797 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U798 ( .A(n706), .B(n705), .ZN(n712) );
  XNOR2_X1 U799 ( .A(G1961), .B(KEYINPUT90), .ZN(n1001) );
  NAND2_X1 U800 ( .A1(n1001), .A2(n728), .ZN(n709) );
  XOR2_X1 U801 ( .A(G2078), .B(KEYINPUT25), .Z(n944) );
  NAND2_X1 U802 ( .A1(n707), .A2(n944), .ZN(n708) );
  NAND2_X1 U803 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U804 ( .A(n710), .B(KEYINPUT91), .Z(n720) );
  NOR2_X1 U805 ( .A1(G301), .A2(n720), .ZN(n711) );
  XNOR2_X1 U806 ( .A(n713), .B(KEYINPUT93), .ZN(n726) );
  NOR2_X1 U807 ( .A1(G1966), .A2(n811), .ZN(n739) );
  NOR2_X1 U808 ( .A1(G2084), .A2(n728), .ZN(n737) );
  NOR2_X1 U809 ( .A1(n739), .A2(n737), .ZN(n714) );
  XNOR2_X1 U810 ( .A(KEYINPUT94), .B(n714), .ZN(n715) );
  NAND2_X1 U811 ( .A1(n715), .A2(G8), .ZN(n718) );
  XOR2_X1 U812 ( .A(KEYINPUT30), .B(KEYINPUT95), .Z(n716) );
  NOR2_X1 U813 ( .A1(n719), .A2(G168), .ZN(n722) );
  AND2_X1 U814 ( .A1(n720), .A2(G301), .ZN(n721) );
  NOR2_X1 U815 ( .A1(n722), .A2(n721), .ZN(n724) );
  XNOR2_X1 U816 ( .A(n724), .B(n723), .ZN(n725) );
  NAND2_X1 U817 ( .A1(n726), .A2(n725), .ZN(n738) );
  NAND2_X1 U818 ( .A1(n738), .A2(G286), .ZN(n735) );
  INV_X1 U819 ( .A(G8), .ZN(n733) );
  NOR2_X1 U820 ( .A1(G1971), .A2(n811), .ZN(n727) );
  XOR2_X1 U821 ( .A(KEYINPUT97), .B(n727), .Z(n730) );
  NOR2_X1 U822 ( .A1(G2090), .A2(n728), .ZN(n729) );
  NOR2_X1 U823 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U824 ( .A1(G303), .A2(n731), .ZN(n732) );
  OR2_X1 U825 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U826 ( .A(n736), .B(KEYINPUT32), .ZN(n744) );
  NAND2_X1 U827 ( .A1(G8), .A2(n737), .ZN(n742) );
  INV_X1 U828 ( .A(n738), .ZN(n740) );
  NOR2_X1 U829 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U830 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U831 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n751) );
  NOR2_X1 U833 ( .A1(G303), .A2(G1971), .ZN(n746) );
  NOR2_X1 U834 ( .A1(n751), .A2(n746), .ZN(n977) );
  NAND2_X1 U835 ( .A1(n807), .A2(n977), .ZN(n747) );
  NAND2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n973) );
  NAND2_X1 U837 ( .A1(n747), .A2(n973), .ZN(n748) );
  NOR2_X1 U838 ( .A1(n811), .A2(n513), .ZN(n749) );
  XNOR2_X1 U839 ( .A(n749), .B(KEYINPUT64), .ZN(n750) );
  NOR2_X1 U840 ( .A1(KEYINPUT33), .A2(n750), .ZN(n754) );
  NAND2_X1 U841 ( .A1(n751), .A2(KEYINPUT33), .ZN(n752) );
  NOR2_X1 U842 ( .A1(n752), .A2(n811), .ZN(n753) );
  XOR2_X1 U843 ( .A(G1981), .B(KEYINPUT100), .Z(n755) );
  XNOR2_X1 U844 ( .A(G305), .B(n755), .ZN(n964) );
  XNOR2_X1 U845 ( .A(G1986), .B(G290), .ZN(n974) );
  INV_X1 U846 ( .A(n756), .ZN(n757) );
  NOR2_X1 U847 ( .A1(n758), .A2(n757), .ZN(n802) );
  AND2_X1 U848 ( .A1(n974), .A2(n802), .ZN(n789) );
  NAND2_X1 U849 ( .A1(G140), .A2(n870), .ZN(n760) );
  NAND2_X1 U850 ( .A1(G104), .A2(n871), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U852 ( .A(KEYINPUT34), .B(n761), .ZN(n767) );
  NAND2_X1 U853 ( .A1(G116), .A2(n866), .ZN(n763) );
  NAND2_X1 U854 ( .A1(G128), .A2(n867), .ZN(n762) );
  NAND2_X1 U855 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U856 ( .A(KEYINPUT35), .B(n764), .ZN(n765) );
  XNOR2_X1 U857 ( .A(KEYINPUT87), .B(n765), .ZN(n766) );
  NOR2_X1 U858 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U859 ( .A(n768), .B(KEYINPUT36), .ZN(n769) );
  XNOR2_X1 U860 ( .A(n769), .B(KEYINPUT88), .ZN(n882) );
  XNOR2_X1 U861 ( .A(KEYINPUT37), .B(G2067), .ZN(n800) );
  NOR2_X1 U862 ( .A1(n882), .A2(n800), .ZN(n929) );
  NAND2_X1 U863 ( .A1(n802), .A2(n929), .ZN(n798) );
  NAND2_X1 U864 ( .A1(G131), .A2(n870), .ZN(n771) );
  NAND2_X1 U865 ( .A1(G107), .A2(n866), .ZN(n770) );
  NAND2_X1 U866 ( .A1(n771), .A2(n770), .ZN(n775) );
  NAND2_X1 U867 ( .A1(G95), .A2(n871), .ZN(n773) );
  NAND2_X1 U868 ( .A1(G119), .A2(n867), .ZN(n772) );
  NAND2_X1 U869 ( .A1(n773), .A2(n772), .ZN(n774) );
  OR2_X1 U870 ( .A1(n775), .A2(n774), .ZN(n851) );
  NAND2_X1 U871 ( .A1(G1991), .A2(n851), .ZN(n776) );
  XNOR2_X1 U872 ( .A(n776), .B(KEYINPUT89), .ZN(n785) );
  NAND2_X1 U873 ( .A1(G141), .A2(n870), .ZN(n778) );
  NAND2_X1 U874 ( .A1(G117), .A2(n866), .ZN(n777) );
  NAND2_X1 U875 ( .A1(n778), .A2(n777), .ZN(n781) );
  NAND2_X1 U876 ( .A1(n871), .A2(G105), .ZN(n779) );
  XOR2_X1 U877 ( .A(KEYINPUT38), .B(n779), .Z(n780) );
  NOR2_X1 U878 ( .A1(n781), .A2(n780), .ZN(n783) );
  NAND2_X1 U879 ( .A1(n867), .A2(G129), .ZN(n782) );
  NAND2_X1 U880 ( .A1(n783), .A2(n782), .ZN(n863) );
  AND2_X1 U881 ( .A1(G1996), .A2(n863), .ZN(n784) );
  NOR2_X1 U882 ( .A1(n785), .A2(n784), .ZN(n931) );
  INV_X1 U883 ( .A(n802), .ZN(n786) );
  NOR2_X1 U884 ( .A1(n931), .A2(n786), .ZN(n794) );
  INV_X1 U885 ( .A(n794), .ZN(n787) );
  NAND2_X1 U886 ( .A1(n798), .A2(n787), .ZN(n788) );
  NOR2_X1 U887 ( .A1(n789), .A2(n788), .ZN(n804) );
  AND2_X1 U888 ( .A1(n964), .A2(n804), .ZN(n790) );
  NAND2_X1 U889 ( .A1(n791), .A2(n790), .ZN(n819) );
  NOR2_X1 U890 ( .A1(G1996), .A2(n863), .ZN(n920) );
  NOR2_X1 U891 ( .A1(G1991), .A2(n851), .ZN(n925) );
  NOR2_X1 U892 ( .A1(G1986), .A2(G290), .ZN(n792) );
  NOR2_X1 U893 ( .A1(n925), .A2(n792), .ZN(n793) );
  NOR2_X1 U894 ( .A1(n794), .A2(n793), .ZN(n795) );
  XOR2_X1 U895 ( .A(KEYINPUT101), .B(n795), .Z(n796) );
  NOR2_X1 U896 ( .A1(n920), .A2(n796), .ZN(n797) );
  XNOR2_X1 U897 ( .A(n797), .B(KEYINPUT39), .ZN(n799) );
  NAND2_X1 U898 ( .A1(n799), .A2(n798), .ZN(n801) );
  NAND2_X1 U899 ( .A1(n882), .A2(n800), .ZN(n936) );
  NAND2_X1 U900 ( .A1(n801), .A2(n936), .ZN(n803) );
  NAND2_X1 U901 ( .A1(n803), .A2(n802), .ZN(n817) );
  INV_X1 U902 ( .A(n804), .ZN(n815) );
  NOR2_X1 U903 ( .A1(G2090), .A2(G303), .ZN(n805) );
  NAND2_X1 U904 ( .A1(G8), .A2(n805), .ZN(n806) );
  NAND2_X1 U905 ( .A1(n807), .A2(n806), .ZN(n808) );
  AND2_X1 U906 ( .A1(n808), .A2(n811), .ZN(n813) );
  NOR2_X1 U907 ( .A1(G1981), .A2(G305), .ZN(n809) );
  XOR2_X1 U908 ( .A(n809), .B(KEYINPUT24), .Z(n810) );
  NOR2_X1 U909 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U910 ( .A1(n813), .A2(n812), .ZN(n814) );
  OR2_X1 U911 ( .A1(n815), .A2(n814), .ZN(n816) );
  AND2_X1 U912 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U914 ( .A(KEYINPUT40), .B(n820), .ZN(G329) );
  NAND2_X1 U915 ( .A1(n821), .A2(G2106), .ZN(n822) );
  XOR2_X1 U916 ( .A(KEYINPUT105), .B(n822), .Z(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n823) );
  NAND2_X1 U918 ( .A1(G661), .A2(n823), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n824) );
  XNOR2_X1 U920 ( .A(KEYINPUT106), .B(n824), .ZN(n826) );
  NAND2_X1 U921 ( .A1(n826), .A2(n825), .ZN(G188) );
  INV_X1 U923 ( .A(G120), .ZN(G236) );
  INV_X1 U924 ( .A(G108), .ZN(G238) );
  INV_X1 U925 ( .A(G69), .ZN(G235) );
  NOR2_X1 U926 ( .A1(n828), .A2(n827), .ZN(G325) );
  INV_X1 U927 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U928 ( .A(G2454), .B(G2451), .ZN(n837) );
  XNOR2_X1 U929 ( .A(G2430), .B(G2446), .ZN(n835) );
  XOR2_X1 U930 ( .A(G2435), .B(G2427), .Z(n830) );
  XNOR2_X1 U931 ( .A(KEYINPUT102), .B(G2438), .ZN(n829) );
  XNOR2_X1 U932 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U933 ( .A(n831), .B(G2443), .Z(n833) );
  XNOR2_X1 U934 ( .A(G1341), .B(G1348), .ZN(n832) );
  XNOR2_X1 U935 ( .A(n833), .B(n832), .ZN(n834) );
  XNOR2_X1 U936 ( .A(n835), .B(n834), .ZN(n836) );
  XNOR2_X1 U937 ( .A(n837), .B(n836), .ZN(n838) );
  NAND2_X1 U938 ( .A1(n838), .A2(G14), .ZN(n839) );
  XOR2_X1 U939 ( .A(KEYINPUT103), .B(n839), .Z(n911) );
  XOR2_X1 U940 ( .A(KEYINPUT104), .B(n911), .Z(G401) );
  NAND2_X1 U941 ( .A1(G100), .A2(n871), .ZN(n841) );
  NAND2_X1 U942 ( .A1(G112), .A2(n866), .ZN(n840) );
  NAND2_X1 U943 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U944 ( .A(KEYINPUT112), .B(n842), .ZN(n848) );
  NAND2_X1 U945 ( .A1(G124), .A2(n867), .ZN(n843) );
  XOR2_X1 U946 ( .A(KEYINPUT44), .B(n843), .Z(n844) );
  XNOR2_X1 U947 ( .A(n844), .B(KEYINPUT111), .ZN(n846) );
  NAND2_X1 U948 ( .A1(G136), .A2(n870), .ZN(n845) );
  NAND2_X1 U949 ( .A1(n846), .A2(n845), .ZN(n847) );
  NOR2_X1 U950 ( .A1(n848), .A2(n847), .ZN(G162) );
  XOR2_X1 U951 ( .A(KEYINPUT113), .B(KEYINPUT115), .Z(n849) );
  XNOR2_X1 U952 ( .A(n926), .B(n849), .ZN(n850) );
  XNOR2_X1 U953 ( .A(KEYINPUT48), .B(n850), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n851), .B(KEYINPUT46), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U956 ( .A(n854), .B(G162), .Z(n865) );
  NAND2_X1 U957 ( .A1(G139), .A2(n870), .ZN(n856) );
  NAND2_X1 U958 ( .A1(G103), .A2(n871), .ZN(n855) );
  NAND2_X1 U959 ( .A1(n856), .A2(n855), .ZN(n862) );
  NAND2_X1 U960 ( .A1(n866), .A2(G115), .ZN(n857) );
  XNOR2_X1 U961 ( .A(n857), .B(KEYINPUT114), .ZN(n859) );
  NAND2_X1 U962 ( .A1(G127), .A2(n867), .ZN(n858) );
  NAND2_X1 U963 ( .A1(n859), .A2(n858), .ZN(n860) );
  XOR2_X1 U964 ( .A(KEYINPUT47), .B(n860), .Z(n861) );
  NOR2_X1 U965 ( .A1(n862), .A2(n861), .ZN(n915) );
  XOR2_X1 U966 ( .A(n863), .B(n915), .Z(n864) );
  XNOR2_X1 U967 ( .A(n865), .B(n864), .ZN(n878) );
  NAND2_X1 U968 ( .A1(G118), .A2(n866), .ZN(n869) );
  NAND2_X1 U969 ( .A1(G130), .A2(n867), .ZN(n868) );
  NAND2_X1 U970 ( .A1(n869), .A2(n868), .ZN(n876) );
  NAND2_X1 U971 ( .A1(G142), .A2(n870), .ZN(n873) );
  NAND2_X1 U972 ( .A1(G106), .A2(n871), .ZN(n872) );
  NAND2_X1 U973 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U974 ( .A(KEYINPUT45), .B(n874), .Z(n875) );
  NOR2_X1 U975 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U976 ( .A(n878), .B(n877), .Z(n880) );
  XNOR2_X1 U977 ( .A(G164), .B(G160), .ZN(n879) );
  XNOR2_X1 U978 ( .A(n880), .B(n879), .ZN(n881) );
  XOR2_X1 U979 ( .A(n882), .B(n881), .Z(n883) );
  NOR2_X1 U980 ( .A1(G37), .A2(n883), .ZN(G395) );
  XOR2_X1 U981 ( .A(KEYINPUT107), .B(n884), .Z(G319) );
  XNOR2_X1 U982 ( .A(G286), .B(n967), .ZN(n886) );
  XNOR2_X1 U983 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U984 ( .A(n887), .B(G171), .ZN(n888) );
  NOR2_X1 U985 ( .A1(G37), .A2(n888), .ZN(G397) );
  XOR2_X1 U986 ( .A(G2096), .B(KEYINPUT43), .Z(n890) );
  XNOR2_X1 U987 ( .A(G2090), .B(G2678), .ZN(n889) );
  XNOR2_X1 U988 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U989 ( .A(n891), .B(KEYINPUT108), .Z(n893) );
  XNOR2_X1 U990 ( .A(G2067), .B(G2072), .ZN(n892) );
  XNOR2_X1 U991 ( .A(n893), .B(n892), .ZN(n897) );
  XOR2_X1 U992 ( .A(KEYINPUT42), .B(G2100), .Z(n895) );
  XNOR2_X1 U993 ( .A(G2078), .B(G2084), .ZN(n894) );
  XNOR2_X1 U994 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n897), .B(n896), .ZN(G227) );
  XOR2_X1 U996 ( .A(G2474), .B(G1976), .Z(n899) );
  XNOR2_X1 U997 ( .A(G1986), .B(G1956), .ZN(n898) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U999 ( .A(n900), .B(KEYINPUT109), .Z(n902) );
  XNOR2_X1 U1000 ( .A(G1996), .B(G1991), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n906) );
  XOR2_X1 U1002 ( .A(G1981), .B(G1971), .Z(n904) );
  XNOR2_X1 U1003 ( .A(G1966), .B(G1961), .ZN(n903) );
  XNOR2_X1 U1004 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1005 ( .A(n906), .B(n905), .Z(n908) );
  XNOR2_X1 U1006 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n907) );
  XNOR2_X1 U1007 ( .A(n908), .B(n907), .ZN(G229) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n909) );
  XOR2_X1 U1009 ( .A(KEYINPUT49), .B(n909), .Z(n910) );
  NAND2_X1 U1010 ( .A1(n911), .A2(n910), .ZN(n912) );
  NOR2_X1 U1011 ( .A1(G397), .A2(n912), .ZN(n913) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n913), .ZN(n914) );
  NOR2_X1 U1013 ( .A1(G395), .A2(n914), .ZN(G308) );
  INV_X1 U1014 ( .A(G308), .ZN(G225) );
  INV_X1 U1015 ( .A(G96), .ZN(G221) );
  XOR2_X1 U1016 ( .A(G2072), .B(n915), .Z(n917) );
  XOR2_X1 U1017 ( .A(G164), .B(G2078), .Z(n916) );
  NOR2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1019 ( .A(KEYINPUT50), .B(n918), .ZN(n923) );
  XOR2_X1 U1020 ( .A(G2090), .B(G162), .Z(n919) );
  NOR2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1022 ( .A(KEYINPUT51), .B(n921), .Z(n922) );
  NAND2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n935) );
  XOR2_X1 U1024 ( .A(G160), .B(G2084), .Z(n924) );
  NOR2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n927) );
  NAND2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1028 ( .A(KEYINPUT116), .B(n930), .ZN(n932) );
  NAND2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1030 ( .A(KEYINPUT117), .B(n933), .Z(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n937) );
  NAND2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1033 ( .A(KEYINPUT52), .B(n938), .ZN(n939) );
  NAND2_X1 U1034 ( .A1(n939), .A2(G29), .ZN(n1021) );
  XNOR2_X1 U1035 ( .A(G2067), .B(G26), .ZN(n941) );
  XNOR2_X1 U1036 ( .A(G33), .B(G2072), .ZN(n940) );
  NOR2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n949) );
  XNOR2_X1 U1038 ( .A(G32), .B(n942), .ZN(n943) );
  NAND2_X1 U1039 ( .A1(n943), .A2(G28), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(G27), .B(n944), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(KEYINPUT118), .B(n945), .ZN(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(G25), .B(G1991), .ZN(n950) );
  NOR2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1046 ( .A(KEYINPUT53), .B(n952), .Z(n956) );
  XNOR2_X1 U1047 ( .A(KEYINPUT54), .B(G34), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(n953), .B(KEYINPUT119), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(G2084), .B(n954), .ZN(n955) );
  NAND2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(G35), .B(G2090), .ZN(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(n959), .B(KEYINPUT120), .ZN(n960) );
  NOR2_X1 U1054 ( .A1(G29), .A2(n960), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(KEYINPUT55), .B(n961), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(n962), .A2(G11), .ZN(n1019) );
  INV_X1 U1057 ( .A(G16), .ZN(n1015) );
  XNOR2_X1 U1058 ( .A(KEYINPUT56), .B(KEYINPUT121), .ZN(n963) );
  XNOR2_X1 U1059 ( .A(n1015), .B(n963), .ZN(n990) );
  XNOR2_X1 U1060 ( .A(G1966), .B(G168), .ZN(n965) );
  NAND2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1062 ( .A(KEYINPUT57), .B(n966), .ZN(n988) );
  XOR2_X1 U1063 ( .A(n685), .B(G1341), .Z(n985) );
  XNOR2_X1 U1064 ( .A(n967), .B(G1348), .ZN(n969) );
  XNOR2_X1 U1065 ( .A(G301), .B(G1961), .ZN(n968) );
  NOR2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n970) );
  XOR2_X1 U1067 ( .A(KEYINPUT122), .B(n970), .Z(n982) );
  XNOR2_X1 U1068 ( .A(n991), .B(G299), .ZN(n972) );
  NAND2_X1 U1069 ( .A1(G1971), .A2(G303), .ZN(n971) );
  NAND2_X1 U1070 ( .A1(n972), .A2(n971), .ZN(n979) );
  INV_X1 U1071 ( .A(n973), .ZN(n975) );
  NOR2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(KEYINPUT123), .B(n980), .ZN(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(KEYINPUT124), .B(n983), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(KEYINPUT125), .B(n986), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n1017) );
  XNOR2_X1 U1082 ( .A(G20), .B(n991), .ZN(n995) );
  XNOR2_X1 U1083 ( .A(G1341), .B(G19), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(G1981), .B(G6), .ZN(n992) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n998) );
  XOR2_X1 U1087 ( .A(KEYINPUT59), .B(G1348), .Z(n996) );
  XNOR2_X1 U1088 ( .A(G4), .B(n996), .ZN(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1090 ( .A(KEYINPUT60), .B(n999), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(n1000), .B(KEYINPUT126), .ZN(n1005) );
  XNOR2_X1 U1092 ( .A(n1001), .B(G5), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(G21), .B(G1966), .ZN(n1002) );
  NOR2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1012) );
  XNOR2_X1 U1096 ( .A(G1971), .B(G22), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(G23), .B(G1976), .ZN(n1006) );
  NOR2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  XOR2_X1 U1099 ( .A(G1986), .B(G24), .Z(n1008) );
  NAND2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1101 ( .A(KEYINPUT58), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1103 ( .A(KEYINPUT61), .B(n1013), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1108 ( .A(n1022), .B(KEYINPUT127), .ZN(n1023) );
  XNOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1023), .ZN(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

