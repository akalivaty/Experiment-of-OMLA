//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT67), .B(G953), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G227), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n192), .B(KEYINPUT73), .ZN(new_n193));
  XNOR2_X1  g007(.A(G110), .B(G140), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n193), .B(new_n194), .ZN(new_n195));
  XOR2_X1   g009(.A(new_n195), .B(KEYINPUT74), .Z(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT10), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n199), .A2(KEYINPUT1), .A3(G146), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n200), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n205), .A2(KEYINPUT1), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(new_n202), .A3(new_n203), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n198), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  INV_X1    g024(.A(G104), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G107), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G104), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n210), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n213), .A2(G104), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT3), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n217), .B1(new_n211), .B2(G107), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n213), .A2(KEYINPUT3), .A3(G104), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n216), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n215), .B1(new_n220), .B2(new_n210), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n209), .A2(new_n221), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n213), .A2(KEYINPUT3), .A3(G104), .ZN(new_n223));
  AOI21_X1  g037(.A(KEYINPUT3), .B1(new_n213), .B2(G104), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n212), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT4), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(G101), .ZN(new_n227));
  XNOR2_X1  g041(.A(G143), .B(G146), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n229));
  OAI211_X1 g043(.A(KEYINPUT0), .B(G128), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  INV_X1    g045(.A(new_n229), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n204), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n227), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT4), .B1(new_n220), .B2(new_n210), .ZN(new_n235));
  AOI211_X1 g049(.A(G101), .B(new_n216), .C1(new_n218), .C2(new_n219), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT75), .B1(new_n234), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n225), .A2(G101), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n220), .A2(new_n210), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(KEYINPUT4), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n230), .A2(new_n233), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT75), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n241), .A2(new_n243), .A3(new_n244), .A4(new_n227), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n222), .B1(new_n238), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT76), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n208), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n228), .A2(KEYINPUT76), .A3(new_n207), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n206), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n221), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n198), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT77), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT77), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n251), .A2(new_n254), .A3(new_n198), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT11), .ZN(new_n257));
  INV_X1    g071(.A(G134), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n257), .B1(new_n258), .B2(G137), .ZN(new_n259));
  INV_X1    g073(.A(G137), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(KEYINPUT11), .A3(G134), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n258), .A2(G137), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G131), .ZN(new_n264));
  INV_X1    g078(.A(G131), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n259), .A2(new_n261), .A3(new_n265), .A4(new_n262), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n246), .A2(new_n256), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT78), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT78), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n246), .A2(new_n256), .A3(new_n271), .A4(new_n268), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n206), .A2(new_n208), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n251), .B1(new_n274), .B2(new_n221), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n267), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n276), .B(KEYINPUT12), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n197), .B1(new_n273), .B2(new_n278), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n246), .A2(new_n256), .ZN(new_n280));
  OR2_X1    g094(.A1(new_n280), .A2(new_n268), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n195), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n273), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT79), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n282), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AOI211_X1 g100(.A(new_n285), .B(new_n195), .C1(new_n270), .C2(new_n272), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n279), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(G469), .B1(new_n289), .B2(G902), .ZN(new_n290));
  INV_X1    g104(.A(G902), .ZN(new_n291));
  XNOR2_X1  g105(.A(KEYINPUT80), .B(G469), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n283), .B1(new_n273), .B2(new_n281), .ZN(new_n293));
  AOI211_X1 g107(.A(new_n195), .B(new_n277), .C1(new_n270), .C2(new_n272), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n291), .B(new_n292), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n190), .B1(new_n290), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT91), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT20), .ZN(new_n298));
  XNOR2_X1  g112(.A(G113), .B(G122), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n299), .B(new_n211), .ZN(new_n300));
  XOR2_X1   g114(.A(KEYINPUT71), .B(G125), .Z(new_n301));
  INV_X1    g115(.A(KEYINPUT16), .ZN(new_n302));
  INV_X1    g116(.A(G140), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  OR2_X1    g118(.A1(KEYINPUT71), .A2(G125), .ZN(new_n305));
  NAND2_X1  g119(.A1(KEYINPUT71), .A2(G125), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(G140), .A3(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(G125), .A2(G140), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g124(.A(G146), .B(new_n304), .C1(new_n310), .C2(new_n302), .ZN(new_n311));
  XNOR2_X1  g125(.A(G125), .B(G140), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT19), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT89), .ZN(new_n314));
  OR2_X1    g128(.A1(new_n313), .A2(KEYINPUT89), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n307), .A2(new_n309), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n201), .B(new_n316), .C1(new_n317), .C2(new_n313), .ZN(new_n318));
  INV_X1    g132(.A(G237), .ZN(new_n319));
  AND2_X1   g133(.A1(KEYINPUT67), .A2(G953), .ZN(new_n320));
  NOR2_X1   g134(.A1(KEYINPUT67), .A2(G953), .ZN(new_n321));
  OAI211_X1 g135(.A(G214), .B(new_n319), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n199), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n191), .A2(G143), .A3(G214), .A4(new_n319), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(new_n324), .A3(new_n265), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n265), .B1(new_n323), .B2(new_n324), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n311), .B(new_n318), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(KEYINPUT18), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n307), .A2(G146), .A3(new_n309), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT88), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AND2_X1   g146(.A1(G125), .A2(G140), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n201), .B1(new_n333), .B2(new_n308), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT72), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n312), .A2(KEYINPUT72), .A3(new_n201), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n307), .A2(KEYINPUT88), .A3(G146), .A4(new_n309), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n332), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(KEYINPUT18), .A2(G131), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n323), .A2(new_n324), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n329), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n300), .B1(new_n328), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n323), .A2(new_n324), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(KEYINPUT17), .A3(G131), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n302), .B1(new_n307), .B2(new_n309), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n305), .A2(new_n306), .ZN(new_n348));
  NOR3_X1   g162(.A1(new_n348), .A2(KEYINPUT16), .A3(G140), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n201), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n346), .A2(new_n350), .A3(new_n311), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n345), .A2(G131), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT17), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n353), .A3(new_n325), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n330), .A2(new_n331), .B1(new_n336), .B2(new_n337), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n323), .A2(new_n324), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n355), .A2(new_n339), .B1(new_n356), .B2(new_n341), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n351), .A2(new_n354), .B1(new_n357), .B2(new_n329), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n344), .B1(new_n358), .B2(new_n300), .ZN(new_n359));
  NOR2_X1   g173(.A1(G475), .A2(G902), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n298), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n328), .A2(new_n343), .ZN(new_n363));
  INV_X1    g177(.A(new_n300), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT17), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n346), .A2(new_n311), .A3(new_n350), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n300), .B(new_n343), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(KEYINPUT20), .A3(new_n360), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n362), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G475), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n354), .A2(new_n350), .A3(new_n311), .A4(new_n346), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n300), .B1(new_n373), .B2(new_n343), .ZN(new_n374));
  AOI21_X1  g188(.A(G902), .B1(new_n374), .B2(KEYINPUT90), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n343), .B1(new_n366), .B2(new_n367), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n364), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT90), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(new_n368), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n372), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n297), .B1(new_n371), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n375), .A2(new_n379), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G475), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT20), .B1(new_n369), .B2(new_n360), .ZN(new_n384));
  AOI211_X1 g198(.A(new_n298), .B(new_n361), .C1(new_n365), .C2(new_n368), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n383), .A2(new_n386), .A3(KEYINPUT91), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n381), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n205), .A2(G143), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n199), .A2(G128), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n258), .ZN(new_n392));
  OAI21_X1  g206(.A(G134), .B1(new_n389), .B2(new_n390), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT94), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AND2_X1   g210(.A1(KEYINPUT66), .A2(G116), .ZN(new_n397));
  NOR2_X1   g211(.A1(KEYINPUT66), .A2(G116), .ZN(new_n398));
  OAI21_X1  g212(.A(G122), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G122), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G116), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n213), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n392), .A2(KEYINPUT94), .A3(new_n393), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n396), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT95), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT66), .ZN(new_n406));
  INV_X1    g220(.A(G116), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(KEYINPUT66), .A2(G116), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n400), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT14), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n405), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n399), .A2(KEYINPUT95), .A3(KEYINPUT14), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n401), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT96), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n412), .A2(KEYINPUT96), .A3(new_n401), .A4(new_n413), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n410), .A2(new_n411), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n404), .B1(new_n419), .B2(G107), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n392), .B(KEYINPUT93), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT92), .ZN(new_n422));
  INV_X1    g236(.A(new_n389), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT13), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n390), .B1(new_n423), .B2(new_n424), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n389), .A2(KEYINPUT92), .A3(KEYINPUT13), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G134), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n399), .A2(new_n401), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G107), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n402), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n421), .A2(new_n429), .A3(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT97), .B1(new_n420), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT97), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n414), .A2(new_n415), .B1(new_n411), .B2(new_n410), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n213), .B1(new_n437), .B2(new_n417), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n436), .B(new_n433), .C1(new_n438), .C2(new_n404), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G217), .ZN(new_n441));
  NOR3_X1   g255(.A1(new_n188), .A2(new_n441), .A3(G953), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n435), .A2(new_n442), .A3(new_n439), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n291), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G478), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(KEYINPUT15), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n448), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n444), .A2(new_n291), .A3(new_n445), .A4(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n388), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n296), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(G234), .A2(G237), .ZN(new_n455));
  INV_X1    g269(.A(G953), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(G952), .A3(new_n456), .ZN(new_n457));
  XOR2_X1   g271(.A(new_n457), .B(KEYINPUT98), .Z(new_n458));
  XOR2_X1   g272(.A(KEYINPUT21), .B(G898), .Z(new_n459));
  INV_X1    g273(.A(new_n191), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(G902), .A3(new_n455), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n458), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(G214), .B1(G237), .B2(G902), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n242), .A2(new_n301), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n206), .A2(new_n208), .A3(new_n348), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT7), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n456), .A2(G224), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n470), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(G110), .B(G122), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n475), .B(KEYINPUT8), .ZN(new_n476));
  OAI21_X1  g290(.A(G119), .B1(new_n397), .B2(new_n398), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n407), .A2(G119), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(KEYINPUT5), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G113), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT5), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n481), .B1(new_n478), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  AND2_X1   g298(.A1(KEYINPUT2), .A2(G113), .ZN(new_n485));
  NOR2_X1   g299(.A1(KEYINPUT2), .A2(G113), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n477), .A2(new_n479), .A3(new_n487), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n484), .A2(new_n488), .A3(new_n221), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n221), .B1(new_n484), .B2(new_n488), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n476), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n468), .A2(KEYINPUT7), .A3(new_n472), .A4(new_n469), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n474), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n488), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n487), .B1(new_n477), .B2(new_n479), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n227), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT81), .B1(new_n496), .B2(new_n237), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT81), .ZN(new_n498));
  OR2_X1    g312(.A1(new_n485), .A2(new_n486), .ZN(new_n499));
  INV_X1    g313(.A(G119), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n500), .B1(new_n408), .B2(new_n409), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n499), .B1(new_n501), .B2(new_n478), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n488), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n241), .A2(new_n498), .A3(new_n503), .A4(new_n227), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n484), .A2(new_n221), .A3(new_n488), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n497), .A2(new_n475), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT82), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n503), .B(new_n227), .C1(new_n236), .C2(new_n235), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n489), .B1(new_n509), .B2(KEYINPUT81), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n510), .A2(KEYINPUT82), .A3(new_n475), .A4(new_n504), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n493), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT84), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n512), .A2(new_n513), .A3(G902), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n513), .B1(new_n512), .B2(G902), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n475), .B1(new_n510), .B2(new_n504), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n518), .A2(KEYINPUT6), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n518), .B1(new_n508), .B2(new_n511), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT6), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT83), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n470), .B(new_n472), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n522), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n523), .B1(new_n522), .B2(new_n525), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n517), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(G210), .B1(G237), .B2(G902), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(KEYINPUT85), .ZN(new_n530));
  XOR2_X1   g344(.A(new_n530), .B(KEYINPUT86), .Z(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT87), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n530), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n534), .B(new_n517), .C1(new_n526), .C2(new_n527), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n508), .A2(new_n511), .ZN(new_n536));
  INV_X1    g350(.A(new_n493), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT84), .B1(new_n538), .B2(new_n291), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n539), .A2(new_n514), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n522), .A2(new_n525), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT83), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n522), .A2(new_n523), .A3(new_n525), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n535), .B1(new_n544), .B2(new_n531), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n533), .B1(new_n545), .B2(KEYINPUT87), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n454), .A2(new_n467), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n267), .A2(new_n230), .A3(new_n233), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT65), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n243), .A2(KEYINPUT65), .A3(new_n267), .ZN(new_n551));
  INV_X1    g365(.A(new_n262), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n258), .A2(G137), .ZN(new_n553));
  OAI21_X1  g367(.A(G131), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n554), .A2(new_n266), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n274), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n550), .A2(new_n551), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT30), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n548), .A2(new_n556), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n560), .A2(new_n558), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n559), .A2(new_n503), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n503), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n548), .A2(new_n564), .A3(new_n556), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n191), .A2(G210), .A3(new_n319), .ZN(new_n566));
  XOR2_X1   g380(.A(KEYINPUT26), .B(G101), .Z(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n568), .B(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n563), .A2(new_n565), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT31), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT31), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n563), .A2(new_n573), .A3(new_n565), .A4(new_n570), .ZN(new_n574));
  INV_X1    g388(.A(new_n570), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT28), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n565), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n548), .A2(new_n564), .A3(new_n556), .A4(KEYINPUT28), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n548), .A2(new_n549), .B1(new_n274), .B2(new_n555), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n564), .B1(new_n580), .B2(new_n551), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n575), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n572), .A2(new_n574), .A3(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(G472), .A2(G902), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT32), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n557), .A2(new_n503), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n588), .A2(new_n570), .A3(new_n577), .A4(new_n578), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT69), .ZN(new_n590));
  AOI21_X1  g404(.A(KEYINPUT29), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n563), .A2(new_n565), .A3(new_n575), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n570), .B1(new_n579), .B2(new_n581), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT69), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n591), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT70), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n548), .A2(new_n564), .A3(new_n556), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n564), .B1(new_n548), .B2(new_n556), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT28), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n596), .B1(new_n599), .B2(new_n577), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n577), .A2(new_n596), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n570), .A2(KEYINPUT29), .ZN(new_n604));
  AOI21_X1  g418(.A(G902), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n595), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(G472), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n583), .A2(KEYINPUT32), .A3(new_n584), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n587), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n441), .B1(G234), .B2(new_n291), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n500), .A2(G128), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT23), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n615), .B1(G119), .B2(new_n205), .ZN(new_n616));
  XNOR2_X1  g430(.A(G119), .B(G128), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT24), .B(G110), .Z(new_n618));
  OAI22_X1  g432(.A1(new_n616), .A2(G110), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(new_n311), .A3(new_n338), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n616), .A2(G110), .B1(new_n617), .B2(new_n618), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n311), .A2(new_n350), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT22), .B(G137), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n620), .A2(new_n623), .ZN(new_n629));
  INV_X1    g443(.A(new_n627), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n632), .A2(KEYINPUT25), .A3(new_n291), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n628), .A2(new_n291), .A3(new_n631), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT25), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n612), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n632), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n611), .A2(G902), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n610), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n547), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G101), .ZN(G3));
  INV_X1    g460(.A(G469), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n273), .A2(new_n278), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n196), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n195), .B1(new_n270), .B2(new_n272), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n281), .B1(new_n650), .B2(KEYINPUT79), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n649), .B1(new_n651), .B2(new_n287), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n647), .B1(new_n652), .B2(new_n291), .ZN(new_n653));
  INV_X1    g467(.A(new_n295), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n189), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(G472), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n656), .B1(new_n583), .B2(new_n291), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT99), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n585), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n657), .A2(new_n659), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n661), .A2(new_n642), .A3(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n655), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT100), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(KEYINPUT100), .B1(new_n655), .B2(new_n663), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n528), .A2(new_n530), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n535), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n435), .A2(new_n442), .A3(new_n439), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n442), .B1(new_n435), .B2(new_n439), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n672), .A2(new_n673), .A3(G902), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n671), .B1(new_n674), .B2(G478), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n446), .A2(KEYINPUT101), .A3(new_n447), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT33), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n678), .B1(new_n672), .B2(new_n673), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n444), .A2(KEYINPUT33), .A3(new_n445), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n447), .A2(G902), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n677), .A2(new_n683), .ZN(new_n684));
  AND4_X1   g498(.A1(new_n466), .A2(new_n670), .A3(new_n388), .A4(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n668), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT34), .B(G104), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G6));
  NOR2_X1   g502(.A1(new_n371), .A2(new_n380), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n452), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n668), .A2(new_n466), .A3(new_n670), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G107), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT102), .B(KEYINPUT35), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G9));
  NAND2_X1  g508(.A1(new_n661), .A2(new_n662), .ZN(new_n695));
  OR2_X1    g509(.A1(new_n629), .A2(KEYINPUT103), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n630), .A2(KEYINPUT36), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n629), .A2(KEYINPUT103), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n697), .B1(new_n696), .B2(new_n698), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n699), .A2(new_n700), .A3(new_n640), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n637), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n695), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n547), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(KEYINPUT37), .B(G110), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G12));
  OAI211_X1 g520(.A(new_n609), .B(new_n189), .C1(new_n653), .C2(new_n654), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  AOI211_X1 g522(.A(new_n465), .B(new_n702), .C1(new_n669), .C2(new_n535), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT104), .B(G900), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n458), .B1(new_n461), .B2(new_n710), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n452), .A2(new_n689), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n708), .A2(new_n709), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G128), .ZN(G30));
  XNOR2_X1  g528(.A(new_n711), .B(KEYINPUT39), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n296), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(KEYINPUT40), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n716), .B(KEYINPUT106), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT40), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n546), .B(KEYINPUT38), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n388), .A2(new_n452), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT105), .ZN(new_n725));
  OR3_X1    g539(.A1(new_n570), .A2(new_n597), .A3(new_n598), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n561), .B1(new_n558), .B2(new_n557), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n597), .B1(new_n727), .B2(new_n503), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n725), .B(new_n726), .C1(new_n728), .C2(new_n575), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n291), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n563), .A2(new_n565), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n570), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n725), .B1(new_n732), .B2(new_n726), .ZN(new_n733));
  OAI21_X1  g547(.A(G472), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n587), .A2(new_n608), .A3(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n724), .A2(new_n735), .A3(new_n464), .A4(new_n702), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n723), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n719), .A2(new_n722), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(KEYINPUT107), .B(G143), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G45));
  AOI22_X1  g554(.A1(new_n675), .A2(new_n676), .B1(new_n681), .B2(new_n682), .ZN(new_n741));
  INV_X1    g555(.A(new_n388), .ZN(new_n742));
  INV_X1    g556(.A(new_n711), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n708), .A2(new_n709), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G146), .ZN(G48));
  OAI21_X1  g560(.A(new_n291), .B1(new_n293), .B2(new_n294), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(G469), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(new_n189), .A3(new_n295), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n610), .A2(new_n749), .A3(new_n643), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n685), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g565(.A(KEYINPUT41), .B(G113), .Z(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT108), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n751), .B(new_n753), .ZN(G15));
  INV_X1    g568(.A(KEYINPUT109), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n465), .B1(new_n669), .B2(new_n535), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n748), .A2(new_n189), .A3(new_n295), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n690), .A2(new_n609), .A3(new_n642), .A4(new_n462), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n755), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n759), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n761), .A2(KEYINPUT109), .A3(new_n756), .A4(new_n757), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G116), .ZN(G18));
  NAND2_X1  g578(.A1(new_n453), .A2(new_n462), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n765), .A2(new_n610), .A3(new_n749), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n709), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G119), .ZN(G21));
  INV_X1    g582(.A(new_n584), .ZN(new_n769));
  INV_X1    g583(.A(new_n574), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n599), .A2(new_n577), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT70), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT110), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n773), .A3(new_n601), .ZN(new_n774));
  OAI21_X1  g588(.A(KEYINPUT110), .B1(new_n600), .B2(new_n602), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(new_n775), .A3(new_n575), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n572), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT111), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n770), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n776), .A2(KEYINPUT111), .A3(new_n572), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n769), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n388), .A2(new_n452), .A3(new_n462), .ZN(new_n782));
  NOR4_X1   g596(.A1(new_n781), .A2(new_n782), .A3(new_n643), .A4(new_n657), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT112), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n783), .A2(new_n784), .A3(new_n756), .A4(new_n757), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n777), .A2(new_n778), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n574), .A3(new_n780), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n584), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n388), .A2(new_n452), .A3(new_n462), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n788), .A2(new_n789), .A3(new_n642), .A4(new_n658), .ZN(new_n790));
  OAI21_X1  g604(.A(KEYINPUT112), .B1(new_n758), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n785), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G122), .ZN(G24));
  NOR3_X1   g607(.A1(new_n781), .A2(new_n657), .A3(new_n702), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n794), .A2(new_n756), .A3(new_n744), .A4(new_n757), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G125), .ZN(G27));
  AND3_X1   g610(.A1(new_n546), .A2(new_n464), .A3(new_n296), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n797), .A2(KEYINPUT42), .A3(new_n644), .A4(new_n744), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT42), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n546), .A2(new_n644), .A3(new_n296), .A4(new_n464), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n684), .A2(new_n388), .A3(new_n711), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G131), .ZN(G33));
  XNOR2_X1  g618(.A(new_n712), .B(KEYINPUT113), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n800), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(new_n258), .ZN(G36));
  INV_X1    g621(.A(KEYINPUT87), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n528), .A2(new_n532), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n808), .B1(new_n809), .B2(new_n535), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n810), .A2(new_n465), .A3(new_n533), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n741), .A2(new_n388), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(KEYINPUT43), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n684), .A2(KEYINPUT43), .A3(new_n742), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n695), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n815), .A2(new_n816), .A3(new_n702), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n811), .B1(new_n817), .B2(KEYINPUT44), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n818), .B1(KEYINPUT44), .B2(new_n817), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT45), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n647), .B1(new_n652), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n289), .A2(KEYINPUT45), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n821), .A2(new_n822), .B1(G469), .B2(G902), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n823), .A2(KEYINPUT46), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n295), .B1(new_n823), .B2(KEYINPUT46), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n189), .A3(new_n715), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT114), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT114), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n826), .A2(new_n829), .A3(new_n189), .A4(new_n715), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n819), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(G137), .ZN(G39));
  INV_X1    g647(.A(KEYINPUT47), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n834), .B1(new_n826), .B2(new_n189), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n834), .B(new_n189), .C1(new_n824), .C2(new_n825), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n811), .A2(new_n610), .A3(new_n643), .A4(new_n744), .ZN(new_n838));
  OR3_X1    g652(.A1(new_n835), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(G140), .ZN(G42));
  NOR2_X1   g654(.A1(new_n815), .A2(new_n458), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n781), .A2(new_n643), .A3(new_n657), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(new_n756), .A3(new_n757), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n844), .A2(G952), .A3(new_n456), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n545), .A2(KEYINPUT87), .ZN(new_n846));
  INV_X1    g660(.A(new_n533), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n848), .A2(new_n465), .A3(new_n749), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n841), .A2(new_n644), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT48), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n735), .A2(new_n643), .A3(new_n458), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n855), .A2(new_n388), .A3(new_n684), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n845), .A2(new_n852), .A3(new_n853), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(KEYINPUT119), .A2(KEYINPUT50), .ZN(new_n858));
  OR2_X1    g672(.A1(KEYINPUT119), .A2(KEYINPUT50), .ZN(new_n859));
  AND4_X1   g673(.A1(new_n465), .A2(new_n723), .A3(new_n757), .A4(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n858), .B1(new_n860), .B2(new_n843), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n841), .A2(new_n794), .A3(new_n849), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n855), .A2(new_n742), .A3(new_n741), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n748), .A2(new_n295), .ZN(new_n866));
  OAI22_X1  g680(.A1(new_n835), .A2(new_n837), .B1(new_n189), .B2(new_n866), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n867), .A2(new_n811), .B1(new_n858), .B2(new_n860), .ZN(new_n868));
  INV_X1    g682(.A(new_n843), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n865), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT51), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n857), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n872), .B1(new_n871), .B2(new_n870), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n874));
  INV_X1    g688(.A(new_n702), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n788), .A2(new_n658), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n876), .A2(new_n801), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n689), .A2(new_n711), .ZN(new_n878));
  NOR4_X1   g692(.A1(new_n610), .A2(new_n452), .A3(new_n702), .A4(new_n878), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n296), .B(new_n811), .C1(new_n877), .C2(new_n879), .ZN(new_n880));
  AOI22_X1  g694(.A1(new_n685), .A2(new_n750), .B1(new_n766), .B2(new_n709), .ZN(new_n881));
  AND4_X1   g695(.A1(new_n763), .A2(new_n792), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n806), .B1(new_n798), .B2(new_n802), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n388), .B1(new_n449), .B2(new_n451), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n466), .B(new_n884), .C1(new_n810), .C2(new_n533), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT116), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT116), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n848), .A2(new_n887), .A3(new_n466), .A4(new_n884), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n886), .A2(new_n888), .A3(new_n666), .A4(new_n667), .ZN(new_n889));
  INV_X1    g703(.A(new_n454), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n546), .A2(new_n467), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n890), .B(new_n891), .C1(new_n644), .C2(new_n703), .ZN(new_n892));
  OR3_X1    g706(.A1(new_n741), .A2(KEYINPUT115), .A3(new_n742), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT115), .B1(new_n741), .B2(new_n742), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n666), .A2(new_n891), .A3(new_n667), .A4(new_n895), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n882), .A2(new_n883), .A3(new_n889), .A4(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n542), .A2(new_n543), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n534), .B1(new_n900), .B2(new_n517), .ZN(new_n901));
  INV_X1    g715(.A(new_n535), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n464), .B(new_n724), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n711), .B(KEYINPUT117), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n637), .A2(new_n701), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n735), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n655), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n899), .B1(new_n904), .B2(new_n909), .ZN(new_n910));
  NOR4_X1   g724(.A1(new_n903), .A2(new_n655), .A3(KEYINPUT118), .A4(new_n908), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n713), .A2(new_n745), .A3(new_n795), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT52), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n713), .A2(new_n745), .A3(new_n795), .ZN(new_n916));
  INV_X1    g730(.A(new_n908), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n296), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT118), .B1(new_n918), .B2(new_n903), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n904), .A2(new_n909), .A3(new_n899), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT52), .B1(new_n916), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n915), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n874), .B1(new_n898), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n889), .A2(new_n896), .A3(new_n892), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n792), .A2(new_n880), .A3(new_n763), .A4(new_n881), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n914), .B1(new_n912), .B2(new_n913), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n916), .A2(KEYINPUT52), .A3(new_n921), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n927), .A2(new_n930), .A3(KEYINPUT53), .A4(new_n883), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n924), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT54), .ZN(new_n933));
  OAI22_X1  g747(.A1(new_n873), .A2(new_n933), .B1(G952), .B2(G953), .ZN(new_n934));
  NOR4_X1   g748(.A1(new_n735), .A2(new_n643), .A3(new_n465), .A4(new_n190), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n866), .B(KEYINPUT49), .Z(new_n936));
  NAND4_X1  g750(.A1(new_n723), .A2(new_n812), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n934), .A2(new_n937), .ZN(G75));
  NOR2_X1   g752(.A1(new_n191), .A2(G952), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n291), .B1(new_n924), .B2(new_n931), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n941), .A2(new_n532), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n522), .B(new_n525), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT55), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT56), .B1(new_n945), .B2(KEYINPUT121), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n946), .B1(KEYINPUT121), .B2(new_n945), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n940), .B1(new_n942), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT56), .B1(new_n941), .B2(new_n530), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT120), .ZN(new_n950));
  OR3_X1    g764(.A1(new_n949), .A2(new_n950), .A3(new_n945), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n950), .B1(new_n949), .B2(new_n945), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n948), .B1(new_n951), .B2(new_n952), .ZN(G51));
  NAND2_X1  g767(.A1(G469), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT57), .Z(new_n955));
  AND2_X1   g769(.A1(new_n932), .A2(KEYINPUT54), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n932), .A2(KEYINPUT54), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n958), .B1(new_n293), .B2(new_n294), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n941), .A2(new_n822), .A3(new_n821), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n939), .B1(new_n959), .B2(new_n960), .ZN(G54));
  NAND3_X1  g775(.A1(new_n941), .A2(KEYINPUT58), .A3(G475), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n962), .A2(new_n359), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n962), .A2(new_n359), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n963), .A2(new_n964), .A3(new_n939), .ZN(G60));
  NAND2_X1  g779(.A1(G478), .A2(G902), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT59), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n681), .B(new_n967), .C1(new_n956), .C2(new_n957), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n940), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n681), .B1(new_n933), .B2(new_n967), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(G63));
  INV_X1    g785(.A(KEYINPUT61), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT123), .ZN(new_n973));
  NAND2_X1  g787(.A1(G217), .A2(G902), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT122), .Z(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT60), .Z(new_n976));
  INV_X1    g790(.A(new_n806), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n803), .A2(new_n977), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n978), .A2(new_n925), .A3(new_n926), .ZN(new_n979));
  AOI21_X1  g793(.A(KEYINPUT53), .B1(new_n979), .B2(new_n930), .ZN(new_n980));
  INV_X1    g794(.A(new_n931), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n976), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n638), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n973), .B1(new_n983), .B2(new_n940), .ZN(new_n984));
  INV_X1    g798(.A(new_n976), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n985), .B1(new_n924), .B2(new_n931), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n973), .B(new_n940), .C1(new_n986), .C2(new_n632), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n699), .A2(new_n700), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n932), .A2(new_n988), .A3(new_n976), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n972), .B1(new_n984), .B2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT124), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n989), .A2(KEYINPUT61), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n940), .B1(new_n986), .B2(new_n632), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n972), .B1(new_n986), .B2(new_n988), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n996), .A2(new_n983), .A3(KEYINPUT124), .A4(new_n940), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n991), .A2(new_n998), .ZN(G66));
  AOI21_X1  g813(.A(new_n456), .B1(new_n459), .B2(G224), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n792), .A2(new_n763), .A3(new_n881), .ZN(new_n1001));
  OR2_X1    g815(.A1(new_n925), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1000), .B1(new_n1002), .B2(new_n191), .ZN(new_n1003));
  INV_X1    g817(.A(new_n522), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1004), .B1(G898), .B2(new_n191), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT125), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1003), .B(new_n1006), .ZN(G69));
  NAND2_X1  g821(.A1(new_n738), .A2(new_n916), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT62), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n738), .A2(KEYINPUT62), .A3(new_n916), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1012), .ZN(new_n1013));
  OR2_X1    g827(.A1(new_n895), .A2(new_n884), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n720), .A2(new_n644), .A3(new_n811), .A4(new_n1014), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n832), .A2(new_n839), .A3(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n191), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(new_n316), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1018), .B1(KEYINPUT19), .B2(new_n310), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n727), .B(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(KEYINPUT126), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1017), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n831), .A2(new_n644), .A3(new_n904), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n978), .A2(new_n913), .ZN(new_n1024));
  AND4_X1   g838(.A1(new_n832), .A2(new_n1023), .A3(new_n839), .A4(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1025), .A2(new_n191), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1020), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1027), .B1(G900), .B2(new_n460), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n191), .B1(G227), .B2(G900), .ZN(new_n1030));
  NAND4_X1  g844(.A1(new_n1022), .A2(new_n1029), .A3(KEYINPUT127), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1030), .A2(KEYINPUT127), .ZN(new_n1032));
  OR2_X1    g846(.A1(new_n1030), .A2(KEYINPUT127), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1021), .ZN(new_n1034));
  NAND4_X1  g848(.A1(new_n1012), .A2(new_n832), .A3(new_n839), .A4(new_n1015), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1034), .B1(new_n1035), .B2(new_n191), .ZN(new_n1036));
  INV_X1    g850(.A(new_n1028), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1037), .B1(new_n1025), .B2(new_n191), .ZN(new_n1038));
  OAI211_X1 g852(.A(new_n1032), .B(new_n1033), .C1(new_n1036), .C2(new_n1038), .ZN(new_n1039));
  AND2_X1   g853(.A1(new_n1031), .A2(new_n1039), .ZN(G72));
  OR2_X1    g854(.A1(new_n1035), .A2(new_n732), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1025), .A2(new_n592), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n1002), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g857(.A1(G472), .A2(G902), .ZN(new_n1044));
  XOR2_X1   g858(.A(new_n1044), .B(KEYINPUT63), .Z(new_n1045));
  INV_X1    g859(.A(new_n732), .ZN(new_n1046));
  NOR2_X1   g860(.A1(new_n1046), .A2(new_n592), .ZN(new_n1047));
  AND3_X1   g861(.A1(new_n932), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n940), .B1(new_n1047), .B2(new_n1045), .ZN(new_n1049));
  NOR3_X1   g863(.A1(new_n1043), .A2(new_n1048), .A3(new_n1049), .ZN(G57));
endmodule


