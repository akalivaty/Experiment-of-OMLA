//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1217, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1272, new_n1273, new_n1274, new_n1275;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G13), .ZN(new_n205));
  OAI211_X1 g0005(.A(new_n205), .B(G250), .C1(G257), .C2(G264), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT0), .ZN(new_n207));
  OAI21_X1  g0007(.A(G50), .B1(G58), .B2(G68), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT65), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT66), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n204), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n207), .B(new_n213), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT67), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n232), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XOR2_X1   g0038(.A(G50), .B(G58), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  AOI21_X1  g0044(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(KEYINPUT3), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT3), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G1698), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G222), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT3), .B(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G223), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(G1698), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n253), .B1(new_n217), .B2(new_n254), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n246), .B1(new_n257), .B2(KEYINPUT68), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(KEYINPUT68), .B2(new_n257), .ZN(new_n259));
  INV_X1    g0059(.A(G274), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n245), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  INV_X1    g0062(.A(G45), .ZN(new_n263));
  AOI21_X1  g0063(.A(G1), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n245), .A2(new_n264), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G226), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n259), .A2(G190), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT71), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n271), .B(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n259), .A2(new_n270), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT70), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(new_n275), .A3(G200), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G50), .A2(G58), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n211), .B1(new_n277), .B2(new_n215), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G20), .A2(G33), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G150), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XOR2_X1   g0082(.A(KEYINPUT8), .B(G58), .Z(new_n283));
  NOR2_X1   g0083(.A1(new_n247), .A2(G20), .ZN(new_n284));
  AOI211_X1 g0084(.A(new_n278), .B(new_n282), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n210), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G13), .ZN(new_n290));
  NOR3_X1   g0090(.A1(new_n290), .A2(new_n211), .A3(G1), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(new_n287), .ZN(new_n292));
  INV_X1    g0092(.A(G1), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G20), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n292), .A2(G50), .A3(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n290), .A2(G1), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G20), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n295), .B1(G50), .B2(new_n297), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n289), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT9), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n276), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n274), .A2(G200), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT70), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n273), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT10), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT10), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n273), .A2(new_n301), .A3(new_n306), .A4(new_n303), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n299), .ZN(new_n309));
  INV_X1    g0109(.A(G169), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n309), .B1(new_n274), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G179), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n259), .A2(new_n312), .A3(new_n270), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n279), .A2(G50), .B1(G20), .B2(new_n215), .ZN(new_n316));
  INV_X1    g0116(.A(new_n284), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n316), .B1(new_n317), .B2(new_n217), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n287), .ZN(new_n319));
  XOR2_X1   g0119(.A(new_n319), .B(KEYINPUT11), .Z(new_n320));
  NAND3_X1  g0120(.A1(new_n292), .A2(G68), .A3(new_n294), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n296), .A2(G20), .A3(new_n215), .ZN(new_n322));
  NAND2_X1  g0122(.A1(KEYINPUT74), .A2(KEYINPUT12), .ZN(new_n323));
  OR2_X1    g0123(.A1(KEYINPUT74), .A2(KEYINPUT12), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n321), .B(new_n325), .C1(new_n323), .C2(new_n322), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n320), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n265), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n328), .B1(G238), .B2(new_n266), .ZN(new_n329));
  NAND2_X1  g0129(.A1(G33), .A2(G97), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n330), .B(KEYINPUT72), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(new_n252), .B2(G226), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n254), .A2(G232), .A3(G1698), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n245), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT73), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT73), .B1(new_n334), .B2(new_n245), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n329), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT13), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT13), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n341), .B(new_n329), .C1(new_n337), .C2(new_n338), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G190), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n327), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G200), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(new_n340), .B2(new_n342), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n335), .B(new_n336), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n341), .B1(new_n349), .B2(new_n329), .ZN(new_n350));
  INV_X1    g0150(.A(new_n342), .ZN(new_n351));
  OAI21_X1  g0151(.A(G169), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT14), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n340), .A2(G179), .A3(new_n342), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT14), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n343), .A2(new_n355), .A3(G169), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n353), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n327), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n348), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT15), .B(G87), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n361), .A2(new_n284), .B1(G20), .B2(G77), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n283), .A2(new_n279), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n288), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n292), .A2(G77), .A3(new_n294), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(G77), .B2(new_n297), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n251), .A2(G107), .ZN(new_n368));
  INV_X1    g0168(.A(G1698), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n254), .A2(new_n369), .ZN(new_n370));
  OAI221_X1 g0170(.A(new_n368), .B1(new_n370), .B2(new_n229), .C1(new_n216), .C2(new_n256), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n245), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n328), .B1(G244), .B2(new_n266), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT69), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT69), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n372), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n367), .B1(new_n378), .B2(new_n312), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n375), .A2(new_n310), .A3(new_n377), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n378), .A2(G190), .ZN(new_n383));
  INV_X1    g0183(.A(new_n367), .ZN(new_n384));
  INV_X1    g0184(.A(new_n378), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n384), .B1(new_n385), .B2(G200), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n382), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n308), .A2(new_n315), .A3(new_n359), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n283), .A2(new_n294), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n288), .A2(new_n297), .ZN(new_n390));
  OAI22_X1  g0190(.A1(new_n389), .A2(new_n390), .B1(new_n297), .B2(new_n283), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n254), .B2(G20), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n211), .A2(KEYINPUT7), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n251), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n215), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  AND2_X1   g0197(.A1(G58), .A2(G68), .ZN(new_n398));
  NOR2_X1   g0198(.A1(G58), .A2(G68), .ZN(new_n399));
  OAI21_X1  g0199(.A(G20), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT75), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT75), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n402), .B(G20), .C1(new_n398), .C2(new_n399), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n279), .A2(G159), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n401), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n397), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n288), .B1(new_n406), .B2(KEYINPUT16), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT77), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n400), .A2(KEYINPUT75), .B1(G159), .B2(new_n279), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n249), .A2(G33), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n247), .A2(KEYINPUT3), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n211), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT76), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n249), .B2(G33), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n247), .A2(KEYINPUT76), .A3(KEYINPUT3), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(new_n250), .A3(new_n415), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n392), .A2(new_n412), .B1(new_n416), .B2(new_n395), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n403), .B(new_n409), .C1(new_n417), .C2(new_n215), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT16), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n408), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n416), .A2(new_n395), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n215), .B1(new_n421), .B2(new_n393), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n408), .B(new_n419), .C1(new_n422), .C2(new_n405), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n407), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT78), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n419), .B1(new_n422), .B2(new_n405), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT77), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n423), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n430), .A2(KEYINPUT78), .A3(new_n407), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n391), .B1(new_n427), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n266), .A2(G232), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n433), .B(KEYINPUT79), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n268), .A2(G1698), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(G223), .B2(G1698), .ZN(new_n436));
  INV_X1    g0236(.A(G87), .ZN(new_n437));
  OAI22_X1  g0237(.A1(new_n436), .A2(new_n251), .B1(new_n247), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n328), .B1(new_n438), .B2(new_n245), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(G169), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n434), .A2(new_n439), .A3(G179), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT18), .B1(new_n432), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n440), .A2(new_n346), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(G190), .B2(new_n440), .ZN(new_n447));
  INV_X1    g0247(.A(new_n391), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n401), .A2(new_n403), .A3(new_n404), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT7), .B1(new_n251), .B2(new_n211), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n254), .A2(new_n394), .ZN(new_n451));
  OAI21_X1  g0251(.A(G68), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(new_n452), .A3(KEYINPUT16), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n287), .ZN(new_n454));
  AOI211_X1 g0254(.A(new_n426), .B(new_n454), .C1(new_n429), .C2(new_n423), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT78), .B1(new_n430), .B2(new_n407), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n447), .B(new_n448), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT17), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n448), .B1(new_n455), .B2(new_n456), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT18), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n460), .A2(new_n461), .A3(new_n443), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n427), .A2(new_n431), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n463), .A2(KEYINPUT17), .A3(new_n448), .A4(new_n447), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n445), .A2(new_n459), .A3(new_n462), .A4(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n388), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n254), .A2(new_n211), .A3(G87), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n467), .B(KEYINPUT22), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT23), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(new_n211), .B2(G107), .ZN(new_n470));
  INV_X1    g0270(.A(G107), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(KEYINPUT23), .A3(G20), .ZN(new_n472));
  NAND2_X1  g0272(.A1(G33), .A2(G116), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n470), .A2(new_n472), .B1(new_n474), .B2(new_n211), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n468), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(KEYINPUT24), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT24), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n478), .B1(new_n468), .B2(new_n475), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n287), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n292), .B1(G1), .B2(new_n247), .ZN(new_n481));
  XNOR2_X1  g0281(.A(new_n481), .B(KEYINPUT80), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G107), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n297), .A2(G107), .ZN(new_n484));
  XNOR2_X1  g0284(.A(new_n484), .B(KEYINPUT25), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n480), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n262), .A2(KEYINPUT5), .ZN(new_n487));
  XNOR2_X1  g0287(.A(new_n487), .B(KEYINPUT83), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n262), .A2(KEYINPUT5), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n489), .A2(G1), .A3(new_n263), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n261), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n245), .B1(new_n490), .B2(new_n487), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G264), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n254), .A2(G257), .ZN(new_n494));
  INV_X1    g0294(.A(G294), .ZN(new_n495));
  OAI22_X1  g0295(.A1(new_n494), .A2(new_n369), .B1(new_n247), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G250), .ZN(new_n497));
  OR3_X1    g0297(.A1(new_n370), .A2(KEYINPUT87), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(KEYINPUT87), .B1(new_n370), .B2(new_n497), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n496), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n491), .B(new_n493), .C1(new_n500), .C2(new_n246), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT88), .ZN(new_n502));
  OR3_X1    g0302(.A1(new_n501), .A2(new_n502), .A3(new_n312), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n501), .A2(G169), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n502), .B1(new_n501), .B2(new_n312), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n486), .B(new_n503), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n483), .A2(new_n485), .ZN(new_n507));
  XNOR2_X1  g0307(.A(new_n476), .B(KEYINPUT24), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(new_n287), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n501), .A2(G200), .ZN(new_n510));
  OR2_X1    g0310(.A1(new_n501), .A2(new_n344), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G283), .ZN(new_n514));
  INV_X1    g0314(.A(G97), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n514), .B(new_n211), .C1(G33), .C2(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n516), .B(new_n287), .C1(new_n211), .C2(G116), .ZN(new_n517));
  XNOR2_X1  g0317(.A(new_n517), .B(KEYINPUT20), .ZN(new_n518));
  INV_X1    g0318(.A(G116), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n291), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n481), .B2(new_n519), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g0322(.A(new_n522), .B(KEYINPUT85), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n492), .A2(G270), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n524), .A2(new_n491), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n254), .A2(G264), .A3(G1698), .ZN(new_n526));
  INV_X1    g0326(.A(G303), .ZN(new_n527));
  OAI221_X1 g0327(.A(new_n526), .B1(new_n527), .B2(new_n254), .C1(new_n494), .C2(G1698), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n245), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n310), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n523), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT86), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n532), .A2(KEYINPUT21), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n525), .A2(new_n529), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n534), .A2(new_n312), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n531), .A2(new_n533), .B1(new_n523), .B2(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n523), .B(new_n530), .C1(new_n532), .C2(KEYINPUT21), .ZN(new_n537));
  INV_X1    g0337(.A(new_n523), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n534), .A2(G200), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n538), .B(new_n539), .C1(new_n344), .C2(new_n534), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n536), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  OAI221_X1 g0341(.A(new_n473), .B1(new_n370), .B2(new_n216), .C1(new_n218), .C2(new_n256), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n245), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n293), .A2(new_n260), .A3(G45), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n497), .B1(new_n263), .B2(G1), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n246), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(G190), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n543), .A2(new_n546), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G200), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n254), .A2(new_n211), .A3(G68), .ZN(new_n551));
  XNOR2_X1  g0351(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n317), .A2(new_n515), .ZN(new_n553));
  AOI21_X1  g0353(.A(G20), .B1(new_n331), .B2(new_n552), .ZN(new_n554));
  NOR3_X1   g0354(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n555));
  OAI221_X1 g0355(.A(new_n551), .B1(new_n552), .B2(new_n553), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n556), .A2(new_n287), .B1(new_n291), .B2(new_n360), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n482), .A2(G87), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n548), .A2(new_n550), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n547), .A2(new_n312), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n482), .A2(new_n361), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n549), .A2(new_n310), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n492), .A2(G257), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n491), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n370), .A2(new_n218), .ZN(new_n570));
  OAI221_X1 g0370(.A(new_n514), .B1(new_n497), .B2(new_n256), .C1(new_n570), .C2(KEYINPUT4), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n252), .A2(KEYINPUT4), .A3(G244), .ZN(new_n572));
  OR2_X1    g0372(.A1(new_n572), .A2(KEYINPUT82), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(KEYINPUT82), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n571), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n569), .B1(new_n575), .B2(new_n246), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n310), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n573), .A2(new_n574), .ZN(new_n578));
  INV_X1    g0378(.A(new_n571), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n568), .B1(new_n580), .B2(new_n245), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n312), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT81), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT80), .ZN(new_n584));
  OR2_X1    g0384(.A1(new_n481), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n481), .A2(new_n584), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n515), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n291), .A2(G97), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n583), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n588), .ZN(new_n590));
  OAI211_X1 g0390(.A(KEYINPUT81), .B(new_n590), .C1(new_n482), .C2(new_n515), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n471), .A2(KEYINPUT6), .A3(G97), .ZN(new_n593));
  XOR2_X1   g0393(.A(G97), .B(G107), .Z(new_n594));
  OAI21_X1  g0394(.A(new_n593), .B1(new_n594), .B2(KEYINPUT6), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n595), .A2(G20), .B1(G77), .B2(new_n279), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n471), .B2(new_n417), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n597), .A2(new_n287), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n577), .B(new_n582), .C1(new_n592), .C2(new_n598), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n589), .A2(new_n591), .B1(new_n287), .B2(new_n597), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n581), .A2(G190), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n576), .A2(G200), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n566), .A2(new_n599), .A3(new_n603), .ZN(new_n604));
  AND4_X1   g0404(.A1(new_n466), .A2(new_n513), .A3(new_n541), .A4(new_n604), .ZN(G372));
  NAND3_X1  g0405(.A1(new_n536), .A2(new_n506), .A3(new_n537), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n599), .A2(new_n512), .A3(new_n603), .ZN(new_n608));
  INV_X1    g0408(.A(new_n550), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n557), .A2(new_n558), .ZN(new_n610));
  OAI21_X1  g0410(.A(KEYINPUT89), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT89), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n550), .A2(new_n612), .A3(new_n557), .A4(new_n558), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n611), .A2(new_n548), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n564), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n608), .A2(KEYINPUT90), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT90), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n599), .A2(new_n512), .A3(new_n603), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n618), .B1(new_n619), .B2(new_n615), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n607), .B1(new_n617), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n615), .A2(new_n599), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT26), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT26), .B1(new_n599), .B2(new_n565), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(new_n564), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n466), .B1(new_n621), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n356), .A2(new_n354), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n355), .B1(new_n343), .B2(G169), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n358), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n348), .B2(new_n381), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n459), .A2(new_n464), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n445), .A2(KEYINPUT91), .A3(new_n462), .ZN(new_n634));
  AOI21_X1  g0434(.A(KEYINPUT91), .B1(new_n445), .B2(new_n462), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n314), .B1(new_n637), .B2(new_n308), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n627), .A2(new_n638), .ZN(G369));
  NAND2_X1  g0439(.A1(new_n531), .A2(new_n533), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n523), .A2(new_n535), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(new_n537), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n296), .A2(new_n211), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(G213), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(G343), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n523), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n642), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(KEYINPUT92), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n649), .B1(new_n536), .B2(new_n537), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT92), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n536), .A2(new_n540), .A3(new_n537), .A4(new_n649), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n652), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G330), .ZN(new_n658));
  INV_X1    g0458(.A(new_n648), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT93), .B1(new_n509), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT93), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n486), .A2(new_n661), .A3(new_n648), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n506), .A2(new_n660), .A3(new_n512), .A4(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT94), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n504), .A2(new_n505), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n665), .A2(new_n503), .A3(new_n486), .A4(new_n648), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n663), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n664), .B1(new_n663), .B2(new_n666), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n658), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n642), .A2(new_n659), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n668), .B2(new_n669), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n506), .A2(new_n648), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n671), .A2(new_n677), .ZN(G399));
  INV_X1    g0478(.A(new_n205), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(G41), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  AND4_X1   g0481(.A1(G1), .A2(new_n681), .A3(new_n519), .A4(new_n555), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n682), .B1(new_n209), .B2(new_n680), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n683), .B(KEYINPUT28), .Z(new_n684));
  INV_X1    g0484(.A(G330), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n604), .A2(new_n541), .A3(new_n513), .A4(new_n659), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT31), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n534), .A2(new_n549), .A3(new_n312), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n500), .A2(new_n246), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n689), .B1(G264), .B2(new_n492), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n581), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT30), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n581), .A2(new_n688), .A3(KEYINPUT30), .A4(new_n690), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n547), .A2(G179), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n576), .A2(new_n695), .A3(new_n501), .A4(new_n534), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n693), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n648), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n687), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n697), .A2(KEYINPUT31), .A3(new_n648), .ZN(new_n700));
  XOR2_X1   g0500(.A(new_n700), .B(KEYINPUT95), .Z(new_n701));
  AOI21_X1  g0501(.A(new_n685), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n659), .B1(new_n621), .B2(new_n626), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT29), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n608), .A2(new_n606), .A3(new_n616), .ZN(new_n706));
  INV_X1    g0506(.A(new_n564), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n599), .A2(new_n565), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n707), .B1(new_n708), .B2(new_n623), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n706), .B(new_n709), .C1(new_n623), .C2(new_n622), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(KEYINPUT29), .A3(new_n659), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n702), .B1(new_n705), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n684), .B1(new_n712), .B2(G1), .ZN(G364));
  NOR2_X1   g0513(.A1(new_n290), .A2(G20), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n293), .B1(new_n714), .B2(G45), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n680), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n717), .B1(new_n657), .B2(G330), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(G330), .B2(new_n657), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n290), .A2(new_n247), .A3(KEYINPUT96), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT96), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(G13), .B2(G33), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G20), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n210), .B1(G20), .B2(new_n310), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n679), .A2(new_n254), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(G45), .B2(new_n208), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(G45), .B2(new_n240), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n205), .A2(G355), .A3(new_n254), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(G116), .B2(new_n205), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n727), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n717), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n211), .A2(new_n312), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n736), .A2(G190), .A3(new_n346), .ZN(new_n737));
  INV_X1    g0537(.A(G317), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(KEYINPUT33), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n738), .A2(KEYINPUT33), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n737), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NOR4_X1   g0541(.A1(new_n211), .A2(new_n344), .A3(new_n346), .A4(G179), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G326), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n736), .A2(new_n344), .A3(new_n346), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI221_X1 g0546(.A(new_n741), .B1(new_n527), .B2(new_n743), .C1(new_n744), .C2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G179), .A2(G200), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n211), .B1(new_n748), .B2(G190), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n254), .B(new_n747), .C1(G294), .C2(new_n750), .ZN(new_n751));
  NOR4_X1   g0551(.A1(new_n211), .A2(new_n346), .A3(G179), .A4(G190), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G283), .ZN(new_n754));
  INV_X1    g0554(.A(G329), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n748), .A2(G20), .A3(new_n344), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n753), .A2(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT99), .ZN(new_n758));
  AOI21_X1  g0558(.A(G200), .B1(new_n736), .B2(KEYINPUT97), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n759), .B1(KEYINPUT97), .B2(new_n736), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G190), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n344), .ZN(new_n762));
  AOI22_X1  g0562(.A1(G311), .A2(new_n761), .B1(new_n762), .B2(G322), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n751), .A2(new_n758), .A3(new_n763), .ZN(new_n764));
  AOI22_X1  g0564(.A1(G58), .A2(new_n762), .B1(new_n761), .B2(G77), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT98), .Z(new_n766));
  INV_X1    g0566(.A(new_n737), .ZN(new_n767));
  INV_X1    g0567(.A(new_n756), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G159), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n767), .A2(new_n215), .B1(KEYINPUT32), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n753), .A2(new_n471), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n770), .A2(new_n251), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n743), .A2(new_n437), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(G50), .B2(new_n745), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n749), .A2(new_n515), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(new_n769), .B2(KEYINPUT32), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n772), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n764), .B1(new_n766), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n734), .B1(new_n778), .B2(new_n726), .ZN(new_n779));
  INV_X1    g0579(.A(new_n725), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n779), .B1(new_n657), .B2(new_n780), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n719), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(G396));
  INV_X1    g0583(.A(KEYINPUT101), .ZN(new_n784));
  AND3_X1   g0584(.A1(new_n379), .A2(new_n784), .A3(new_n380), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n784), .B1(new_n379), .B2(new_n380), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n384), .A2(new_n648), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT102), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n789), .B1(new_n386), .B2(new_n383), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n659), .B(new_n792), .C1(new_n621), .C2(new_n626), .ZN(new_n793));
  AOI21_X1  g0593(.A(KEYINPUT90), .B1(new_n608), .B2(new_n616), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n619), .A2(new_n615), .A3(new_n618), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n606), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n625), .A2(new_n564), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(new_n623), .B2(new_n622), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n648), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n787), .A2(new_n790), .B1(new_n382), .B2(new_n648), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n793), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n698), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(new_n686), .B2(KEYINPUT31), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n700), .B(KEYINPUT95), .ZN(new_n805));
  OAI21_X1  g0605(.A(G330), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n717), .B1(new_n802), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n806), .B2(new_n802), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n723), .A2(new_n726), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n717), .B1(G77), .B2(new_n809), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT100), .Z(new_n811));
  AOI22_X1  g0611(.A1(G116), .A2(new_n761), .B1(new_n762), .B2(G294), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n254), .B(new_n775), .C1(G311), .C2(new_n768), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n753), .A2(new_n437), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G303), .B2(new_n745), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n737), .A2(G283), .B1(G107), .B2(new_n742), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n812), .A2(new_n813), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n762), .A2(G143), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n737), .A2(G150), .B1(new_n745), .B2(G137), .ZN(new_n819));
  INV_X1    g0619(.A(new_n761), .ZN(new_n820));
  INV_X1    g0620(.A(G159), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n818), .B(new_n819), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT34), .Z(new_n823));
  INV_X1    g0623(.A(G50), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n743), .A2(new_n824), .B1(new_n753), .B2(new_n215), .ZN(new_n825));
  INV_X1    g0625(.A(G132), .ZN(new_n826));
  INV_X1    g0626(.A(G58), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n254), .B1(new_n756), .B2(new_n826), .C1(new_n827), .C2(new_n749), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n817), .B1(new_n823), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n811), .B1(new_n830), .B2(new_n726), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n801), .B2(new_n724), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n808), .A2(new_n832), .ZN(G384));
  NOR2_X1   g0633(.A1(new_n714), .A2(new_n293), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n406), .A2(KEYINPUT16), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n448), .B1(new_n454), .B2(new_n835), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT105), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n837), .A2(new_n646), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n465), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT106), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n465), .A2(KEYINPUT106), .A3(new_n838), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n432), .A2(new_n646), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT37), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n460), .A2(new_n443), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n457), .ZN(new_n848));
  INV_X1    g0648(.A(new_n646), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n443), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n457), .B1(new_n837), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(KEYINPUT37), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT38), .B1(new_n843), .B2(new_n853), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n465), .A2(KEYINPUT106), .A3(new_n838), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT106), .B1(new_n465), .B2(new_n838), .ZN(new_n856));
  OAI211_X1 g0656(.A(KEYINPUT38), .B(new_n853), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT39), .B1(new_n854), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT39), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n847), .A2(new_n457), .ZN(new_n862));
  OAI21_X1  g0662(.A(KEYINPUT37), .B1(new_n862), .B2(new_n844), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n861), .A2(new_n844), .B1(new_n848), .B2(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n857), .B(new_n860), .C1(new_n864), .C2(KEYINPUT38), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n859), .A2(KEYINPUT107), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n357), .A2(new_n358), .A3(new_n659), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n853), .B1(new_n855), .B2(new_n856), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT38), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n857), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT107), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n872), .A2(new_n873), .A3(KEYINPUT39), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n866), .A2(new_n868), .A3(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n636), .A2(new_n849), .ZN(new_n876));
  INV_X1    g0676(.A(new_n348), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n327), .A2(new_n659), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n630), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n358), .B(new_n648), .C1(new_n357), .C2(new_n348), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n659), .B1(new_n785), .B2(new_n786), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n884), .B(KEYINPUT104), .Z(new_n885));
  AOI21_X1  g0685(.A(new_n883), .B1(new_n793), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n876), .B1(new_n886), .B2(new_n872), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n875), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n705), .A2(new_n466), .A3(new_n711), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n638), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n888), .B(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n699), .A2(new_n700), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n466), .A2(new_n892), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n893), .B(KEYINPUT108), .Z(new_n894));
  INV_X1    g0694(.A(KEYINPUT40), .ZN(new_n895));
  INV_X1    g0695(.A(new_n700), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n804), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n800), .B1(new_n880), .B2(new_n881), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n857), .B1(new_n864), .B2(KEYINPUT38), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n895), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n898), .B(new_n895), .C1(new_n804), .C2(new_n896), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n857), .B2(new_n871), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n894), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n894), .A2(new_n905), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(G330), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n834), .B1(new_n891), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n891), .B2(new_n908), .ZN(new_n910));
  NOR3_X1   g0710(.A1(new_n208), .A2(new_n398), .A3(new_n217), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n215), .A2(G50), .ZN(new_n912));
  OAI211_X1 g0712(.A(G1), .B(new_n290), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  OR2_X1    g0713(.A1(new_n595), .A2(KEYINPUT35), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n595), .A2(KEYINPUT35), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n914), .A2(G116), .A3(new_n212), .A4(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(KEYINPUT103), .B(KEYINPUT36), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n916), .B(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n910), .A2(new_n913), .A3(new_n918), .ZN(G367));
  INV_X1    g0719(.A(new_n669), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n672), .B1(new_n920), .B2(new_n667), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n599), .A2(new_n659), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n599), .B(new_n603), .C1(new_n600), .C2(new_n659), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n925), .A2(KEYINPUT42), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n599), .B1(new_n923), .B2(new_n506), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n925), .A2(KEYINPUT42), .B1(new_n659), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n610), .A2(new_n648), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n564), .A2(new_n929), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(KEYINPUT109), .Z(new_n931));
  NAND2_X1  g0731(.A1(new_n616), .A2(new_n929), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n926), .A2(new_n928), .B1(KEYINPUT43), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n933), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT43), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n671), .ZN(new_n939));
  INV_X1    g0739(.A(new_n924), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n926), .A2(new_n928), .A3(new_n936), .A4(new_n935), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n938), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n941), .B1(new_n938), .B2(new_n942), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n680), .B(KEYINPUT41), .Z(new_n946));
  AOI21_X1  g0746(.A(new_n924), .B1(new_n674), .B2(new_n676), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT44), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n947), .B(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n674), .A2(new_n676), .A3(new_n924), .ZN(new_n950));
  XOR2_X1   g0750(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n950), .B(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n671), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n670), .A2(new_n672), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT111), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n656), .B1(new_n653), .B2(new_n654), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n651), .A2(KEYINPUT92), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n956), .B(G330), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n956), .B1(new_n657), .B2(G330), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n674), .B(new_n955), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n668), .A2(new_n669), .A3(new_n673), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n959), .B1(new_n921), .B2(new_n963), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n965), .A2(KEYINPUT112), .A3(new_n712), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT112), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n711), .B1(new_n799), .B2(KEYINPUT29), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n806), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n962), .A2(new_n964), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n950), .B(new_n951), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n940), .B1(new_n921), .B2(new_n675), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n948), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n947), .A2(KEYINPUT44), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n972), .A2(new_n976), .A3(new_n939), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n954), .A2(new_n966), .A3(new_n971), .A4(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n946), .B1(new_n978), .B2(new_n712), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n945), .B1(new_n979), .B2(new_n716), .ZN(new_n980));
  INV_X1    g0780(.A(new_n728), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n981), .A2(new_n236), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n727), .B1(new_n205), .B2(new_n360), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n717), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n767), .A2(new_n495), .B1(new_n749), .B2(new_n471), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(G311), .B2(new_n745), .ZN(new_n986));
  INV_X1    g0786(.A(new_n762), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n986), .B1(new_n987), .B2(new_n527), .C1(new_n754), .C2(new_n820), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n251), .B1(new_n756), .B2(new_n738), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n753), .A2(new_n515), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT46), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n742), .A2(G116), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n989), .B(new_n990), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n991), .B2(new_n992), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n742), .A2(G58), .B1(new_n768), .B2(G137), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT113), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n987), .B2(new_n281), .C1(new_n824), .C2(new_n820), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n737), .A2(G159), .B1(new_n745), .B2(G143), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n753), .A2(new_n217), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n999), .A2(new_n251), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n998), .B(new_n1000), .C1(new_n215), .C2(new_n749), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n988), .A2(new_n994), .B1(new_n997), .B2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT47), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n984), .B1(new_n1003), .B2(new_n726), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n933), .B2(new_n780), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n980), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(KEYINPUT114), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT114), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n980), .A2(new_n1008), .A3(new_n1005), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(G387));
  NAND2_X1  g0811(.A1(new_n966), .A2(new_n971), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1012), .B(new_n680), .C1(new_n712), .C2(new_n965), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n670), .A2(new_n725), .ZN(new_n1014));
  OR3_X1    g0814(.A1(new_n232), .A2(new_n263), .A3(new_n254), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n263), .B1(new_n215), .B2(new_n217), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT50), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n283), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1017), .B1(new_n1018), .B2(G50), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n283), .A2(KEYINPUT50), .A3(new_n824), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1016), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n519), .B(new_n555), .C1(new_n1021), .C2(new_n254), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n679), .B1(new_n1015), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n727), .B1(new_n471), .B2(new_n205), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n717), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G50), .A2(new_n762), .B1(new_n761), .B2(G68), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n251), .B(new_n990), .C1(G150), .C2(new_n768), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n749), .A2(new_n360), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G77), .B2(new_n742), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G159), .A2(new_n745), .B1(new_n737), .B2(new_n283), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1026), .A2(new_n1027), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n743), .A2(new_n495), .B1(new_n754), .B2(new_n749), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n737), .A2(G311), .B1(new_n745), .B2(G322), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(new_n987), .B2(new_n738), .C1(new_n527), .C2(new_n820), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT48), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1032), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n1035), .B2(new_n1034), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT49), .Z(new_n1038));
  OAI221_X1 g0838(.A(new_n251), .B1(new_n744), .B2(new_n756), .C1(new_n753), .C2(new_n519), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1031), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1025), .B1(new_n1040), .B2(new_n726), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n965), .A2(new_n716), .B1(new_n1014), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1013), .A2(new_n1042), .ZN(G393));
  NAND2_X1  g0843(.A1(new_n954), .A2(new_n977), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n1012), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1045), .A2(new_n680), .A3(new_n978), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n954), .A2(new_n977), .A3(new_n716), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n981), .A2(new_n243), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n727), .B1(new_n515), .B2(new_n205), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n717), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n762), .A2(G311), .B1(G317), .B2(new_n745), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT52), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n254), .B(new_n771), .C1(G322), .C2(new_n768), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n761), .A2(G294), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n737), .A2(G303), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n742), .A2(G283), .B1(new_n750), .B2(G116), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n762), .A2(G159), .B1(G150), .B2(new_n745), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT51), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n251), .B(new_n814), .C1(G143), .C2(new_n768), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n761), .A2(new_n283), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n737), .A2(G50), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n749), .A2(new_n217), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(G68), .B2(new_n742), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .A4(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n1052), .A2(new_n1057), .B1(new_n1059), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1050), .B1(new_n1066), .B2(new_n726), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n924), .B2(new_n780), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1047), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1046), .A2(new_n1069), .ZN(G390));
  NAND3_X1  g0870(.A1(new_n892), .A2(G330), .A3(new_n898), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n886), .A2(new_n868), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n866), .B2(new_n874), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n710), .A2(new_n659), .A3(new_n792), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n884), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n868), .B1(new_n1076), .B2(new_n882), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n901), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1072), .B1(new_n1074), .B2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g0880(.A(G330), .B(new_n801), .C1(new_n804), .C2(new_n805), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n882), .ZN(new_n1083));
  AOI211_X1 g0883(.A(KEYINPUT107), .B(new_n860), .C1(new_n871), .C2(new_n857), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n873), .B1(new_n872), .B2(KEYINPUT39), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1084), .B1(new_n1085), .B2(new_n865), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1078), .B(new_n1083), .C1(new_n1086), .C2(new_n1073), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1080), .A2(new_n1087), .A3(new_n716), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n717), .B1(new_n283), .B2(new_n809), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G97), .A2(new_n761), .B1(new_n762), .B2(G116), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n254), .B(new_n773), .C1(G294), .C2(new_n768), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1063), .B1(G68), .B2(new_n752), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n737), .A2(G107), .B1(new_n745), .B2(G283), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(KEYINPUT54), .B(G143), .ZN(new_n1095));
  INV_X1    g0895(.A(G137), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n820), .A2(new_n1095), .B1(new_n1096), .B2(new_n767), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT115), .Z(new_n1098));
  INV_X1    g0898(.A(G125), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n254), .B1(new_n1099), .B2(new_n756), .C1(new_n753), .C2(new_n824), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT116), .Z(new_n1101));
  NAND2_X1  g0901(.A1(new_n742), .A2(G150), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT53), .Z(new_n1103));
  NAND2_X1  g0903(.A1(new_n762), .A2(G132), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n745), .A2(G128), .B1(new_n750), .B2(G159), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1101), .A2(new_n1103), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1094), .B1(new_n1098), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1089), .B1(new_n1107), .B2(new_n726), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT117), .Z(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n1086), .B2(new_n724), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1088), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1080), .A2(new_n1087), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n793), .A2(new_n885), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1071), .B1(new_n1082), .B2(new_n882), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1076), .B1(new_n1082), .B2(new_n882), .ZN(new_n1115));
  OAI211_X1 g0915(.A(G330), .B(new_n801), .C1(new_n804), .C2(new_n896), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n883), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1113), .A2(new_n1114), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n466), .A2(new_n892), .A3(G330), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n889), .A2(new_n1119), .A3(new_n638), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n681), .B1(new_n1112), .B2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1080), .A2(new_n1087), .A3(new_n1121), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1111), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(G378));
  XNOR2_X1  g0926(.A(new_n1120), .B(KEYINPUT119), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(G330), .B1(new_n902), .B2(new_n904), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n308), .A2(new_n315), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n299), .A2(new_n849), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n1131), .B(KEYINPUT55), .Z(new_n1132));
  AND2_X1   g0932(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1134));
  XOR2_X1   g0934(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  OR3_X1    g0936(.A1(new_n1133), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1136), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1129), .A2(new_n1140), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1139), .B(G330), .C1(new_n902), .C2(new_n904), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n888), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1141), .A2(new_n1142), .A3(new_n875), .A4(new_n887), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1128), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT57), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1148), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n681), .B1(new_n1150), .B2(new_n1128), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1140), .A2(new_n723), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n717), .B1(G50), .B2(new_n809), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n824), .B1(G33), .B2(G41), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(new_n251), .B2(new_n262), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(G107), .A2(new_n762), .B1(new_n761), .B2(new_n361), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n251), .B(new_n262), .C1(new_n756), .C2(new_n754), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(G68), .B2(new_n750), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n745), .A2(G116), .B1(G77), .B2(new_n742), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n753), .A2(new_n827), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G97), .B2(new_n737), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1157), .A2(new_n1159), .A3(new_n1160), .A4(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT58), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1156), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n767), .A2(new_n826), .B1(new_n749), .B2(new_n281), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n746), .A2(new_n1099), .B1(new_n743), .B2(new_n1095), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(G128), .C2(new_n762), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n1096), .B2(new_n820), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n752), .A2(G159), .ZN(new_n1171));
  AOI211_X1 g0971(.A(G33), .B(G41), .C1(new_n768), .C2(G124), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1165), .B1(new_n1164), .B2(new_n1163), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1154), .B1(new_n1175), .B2(new_n726), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1146), .A2(new_n716), .B1(new_n1153), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1152), .A2(new_n1177), .ZN(G375));
  OAI21_X1  g0978(.A(KEYINPUT120), .B1(new_n1118), .B2(new_n715), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1114), .A2(new_n1113), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n715), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT120), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n717), .B1(G68), .B2(new_n809), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(G137), .A2(new_n762), .B1(new_n761), .B2(G150), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n251), .B(new_n1161), .C1(G128), .C2(new_n768), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n746), .A2(new_n826), .B1(new_n821), .B2(new_n743), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n767), .A2(new_n1095), .B1(new_n824), .B2(new_n749), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1186), .A2(new_n1187), .A3(new_n1190), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n254), .B(new_n999), .C1(G303), .C2(new_n768), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1028), .B1(new_n745), .B2(G294), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n737), .A2(G116), .B1(G97), .B2(new_n742), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n471), .A2(new_n820), .B1(new_n987), .B2(new_n754), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1191), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1185), .B1(new_n1197), .B2(new_n726), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n882), .B2(new_n724), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1179), .A2(new_n1184), .A3(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n946), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1122), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1200), .A2(new_n1203), .ZN(G381));
  NAND3_X1  g1004(.A1(new_n1013), .A2(new_n782), .A3(new_n1042), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1205), .A2(G384), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT121), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(G381), .A2(G390), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1207), .A2(new_n1010), .A3(new_n1208), .ZN(new_n1209));
  XOR2_X1   g1009(.A(new_n1209), .B(KEYINPUT122), .Z(new_n1210));
  NAND2_X1  g1010(.A1(new_n1146), .A2(new_n716), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1153), .A2(new_n1176), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n1125), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1210), .A2(new_n1215), .ZN(G407));
  NAND3_X1  g1016(.A1(new_n1214), .A2(new_n647), .A3(new_n1125), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(G407), .A2(G213), .A3(new_n1217), .ZN(G409));
  NAND3_X1  g1018(.A1(G387), .A2(new_n1046), .A3(new_n1069), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n980), .A2(new_n1005), .A3(G390), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(G393), .B(new_n782), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1219), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(G390), .B1(new_n980), .B2(new_n1005), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1221), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(KEYINPUT127), .B1(new_n1226), .B2(new_n1222), .ZN(new_n1227));
  OAI211_X1 g1027(.A(KEYINPUT127), .B(new_n1222), .C1(new_n1221), .C2(new_n1225), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1224), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT124), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1128), .A2(new_n1201), .A3(new_n1146), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1125), .A2(new_n1177), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n647), .A2(G213), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1234), .B(new_n1235), .C1(new_n1214), .C2(new_n1125), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n680), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1202), .A2(KEYINPUT60), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT60), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1118), .A2(new_n1239), .A3(new_n1120), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1237), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1184), .A2(new_n1179), .A3(new_n1199), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT123), .B1(new_n808), .B2(new_n832), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n808), .A2(KEYINPUT123), .A3(new_n832), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n1241), .A2(new_n1242), .B1(new_n1243), .B2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1239), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1247));
  AND4_X1   g1047(.A1(new_n1239), .A2(new_n1180), .A3(new_n1181), .A4(new_n1120), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1122), .B(new_n680), .C1(new_n1247), .C2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1249), .A2(new_n1200), .A3(new_n1244), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1246), .A2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1232), .B1(new_n1236), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G375), .A2(G378), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1251), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1253), .A2(new_n1254), .A3(KEYINPUT124), .A4(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT62), .B1(new_n1252), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1235), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(KEYINPUT126), .A3(G2897), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1246), .A2(new_n1250), .A3(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT126), .B1(new_n1258), .B2(G2897), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1260), .B(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT61), .B1(new_n1236), .B2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(KEYINPUT62), .B1(new_n1236), .B2(new_n1251), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1231), .B1(new_n1257), .B2(new_n1265), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1252), .A2(new_n1256), .A3(new_n1267), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1253), .A2(new_n1254), .A3(KEYINPUT63), .A4(new_n1255), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1268), .A2(new_n1263), .A3(new_n1230), .A4(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1266), .A2(new_n1270), .ZN(G405));
  NAND2_X1  g1071(.A1(new_n1253), .A2(new_n1215), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1255), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1253), .A2(new_n1215), .A3(new_n1251), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1275), .B(new_n1230), .ZN(G402));
endmodule


