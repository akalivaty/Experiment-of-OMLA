

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754;

  XNOR2_X1 U373 ( .A(n523), .B(KEYINPUT33), .ZN(n691) );
  XNOR2_X2 U374 ( .A(n391), .B(n559), .ZN(n722) );
  AND2_X2 U375 ( .A1(n577), .A2(n427), .ZN(n523) );
  NOR2_X1 U376 ( .A1(n692), .A2(n608), .ZN(n602) );
  XNOR2_X1 U377 ( .A(n376), .B(n497), .ZN(n667) );
  NOR2_X1 U378 ( .A1(n628), .A2(n721), .ZN(n630) );
  AND2_X2 U379 ( .A1(n409), .A2(n408), .ZN(n706) );
  AND2_X1 U380 ( .A1(n687), .A2(n617), .ZN(n408) );
  OR2_X1 U381 ( .A1(n686), .A2(KEYINPUT2), .ZN(n409) );
  NAND2_X1 U382 ( .A1(n377), .A2(n386), .ZN(n740) );
  NOR2_X1 U383 ( .A1(KEYINPUT65), .A2(n555), .ZN(n557) );
  NOR2_X1 U384 ( .A1(G902), .A2(n700), .ZN(n522) );
  XNOR2_X1 U385 ( .A(n471), .B(KEYINPUT10), .ZN(n488) );
  INV_X2 U386 ( .A(G953), .ZN(n742) );
  XOR2_X1 U387 ( .A(G146), .B(G125), .Z(n471) );
  NOR2_X1 U388 ( .A1(n749), .A2(n639), .ZN(n556) );
  NAND2_X1 U389 ( .A1(n388), .A2(n387), .ZN(n386) );
  NOR2_X1 U390 ( .A1(n615), .A2(n364), .ZN(n387) );
  INV_X1 U391 ( .A(n616), .ZN(n388) );
  XNOR2_X1 U392 ( .A(G134), .B(n472), .ZN(n503) );
  NOR2_X1 U393 ( .A1(n385), .A2(n652), .ZN(n384) );
  AND2_X1 U394 ( .A1(n615), .A2(n364), .ZN(n385) );
  NAND2_X1 U395 ( .A1(n616), .A2(n364), .ZN(n383) );
  INV_X1 U396 ( .A(KEYINPUT39), .ZN(n372) );
  XNOR2_X1 U397 ( .A(n513), .B(G472), .ZN(n595) );
  XNOR2_X1 U398 ( .A(n595), .B(KEYINPUT6), .ZN(n577) );
  XOR2_X1 U399 ( .A(G101), .B(G110), .Z(n517) );
  XNOR2_X1 U400 ( .A(n448), .B(n447), .ZN(n542) );
  XNOR2_X1 U401 ( .A(KEYINPUT46), .B(KEYINPUT64), .ZN(n605) );
  AND2_X1 U402 ( .A1(n406), .A2(n481), .ZN(n405) );
  INV_X1 U403 ( .A(n683), .ZN(n406) );
  XNOR2_X1 U404 ( .A(G116), .B(G101), .ZN(n504) );
  XNOR2_X1 U405 ( .A(KEYINPUT4), .B(G131), .ZN(n502) );
  XNOR2_X1 U406 ( .A(n514), .B(KEYINPUT72), .ZN(n515) );
  AND2_X1 U407 ( .A1(G227), .A2(n742), .ZN(n514) );
  XNOR2_X1 U408 ( .A(G137), .B(G140), .ZN(n518) );
  XNOR2_X1 U409 ( .A(n733), .B(G146), .ZN(n516) );
  INV_X1 U410 ( .A(n386), .ZN(n380) );
  NOR2_X1 U411 ( .A1(G237), .A2(G902), .ZN(n474) );
  NOR2_X1 U412 ( .A1(n667), .A2(n668), .ZN(n665) );
  AND2_X1 U413 ( .A1(n378), .A2(n383), .ZN(n377) );
  NOR2_X1 U414 ( .A1(n382), .A2(n381), .ZN(n378) );
  INV_X1 U415 ( .A(n754), .ZN(n381) );
  XNOR2_X1 U416 ( .A(n491), .B(n375), .ZN(n374) );
  XNOR2_X1 U417 ( .A(G128), .B(KEYINPUT24), .ZN(n491) );
  XNOR2_X1 U418 ( .A(KEYINPUT23), .B(KEYINPUT85), .ZN(n375) );
  XNOR2_X1 U419 ( .A(G119), .B(G110), .ZN(n490) );
  XNOR2_X1 U420 ( .A(n449), .B(n414), .ZN(n493) );
  INV_X1 U421 ( .A(KEYINPUT8), .ZN(n414) );
  NAND2_X1 U422 ( .A1(n493), .A2(G217), .ZN(n413) );
  XNOR2_X1 U423 ( .A(n450), .B(n412), .ZN(n411) );
  INV_X1 U424 ( .A(KEYINPUT7), .ZN(n412) );
  XNOR2_X1 U425 ( .A(G131), .B(G140), .ZN(n437) );
  XOR2_X1 U426 ( .A(KEYINPUT17), .B(KEYINPUT73), .Z(n466) );
  XNOR2_X1 U427 ( .A(n467), .B(KEYINPUT4), .ZN(n468) );
  AND2_X1 U428 ( .A1(G224), .A2(n742), .ZN(n467) );
  NAND2_X1 U429 ( .A1(n454), .A2(n453), .ZN(n472) );
  NAND2_X1 U430 ( .A1(n421), .A2(n418), .ZN(n692) );
  NAND2_X1 U431 ( .A1(n416), .A2(n415), .ZN(n421) );
  INV_X1 U432 ( .A(n594), .ZN(n415) );
  NAND2_X1 U433 ( .A1(n592), .A2(n372), .ZN(n370) );
  NAND2_X1 U434 ( .A1(n369), .A2(n368), .ZN(n365) );
  NOR2_X1 U435 ( .A1(n592), .A2(n372), .ZN(n368) );
  NAND2_X1 U436 ( .A1(n647), .A2(n359), .ZN(n582) );
  XNOR2_X1 U437 ( .A(G478), .B(n459), .ZN(n543) );
  XNOR2_X1 U438 ( .A(KEYINPUT104), .B(KEYINPUT28), .ZN(n597) );
  XNOR2_X1 U439 ( .A(n533), .B(n532), .ZN(n539) );
  XNOR2_X1 U440 ( .A(n531), .B(KEYINPUT67), .ZN(n532) );
  NOR2_X1 U441 ( .A1(n539), .A2(n577), .ZN(n553) );
  XNOR2_X1 U442 ( .A(n393), .B(n510), .ZN(n426) );
  XNOR2_X1 U443 ( .A(n517), .B(n463), .ZN(n393) );
  INV_X1 U444 ( .A(n750), .ZN(n555) );
  XNOR2_X1 U445 ( .A(n485), .B(n484), .ZN(n498) );
  XOR2_X1 U446 ( .A(KEYINPUT87), .B(KEYINPUT20), .Z(n483) );
  INV_X1 U447 ( .A(n384), .ZN(n382) );
  AND2_X1 U448 ( .A1(n556), .A2(n528), .ZN(n424) );
  AND2_X1 U449 ( .A1(n355), .A2(n390), .ZN(n389) );
  NOR2_X1 U450 ( .A1(G953), .A2(G237), .ZN(n507) );
  XOR2_X1 U451 ( .A(KEYINPUT98), .B(KEYINPUT12), .Z(n440) );
  XNOR2_X1 U452 ( .A(KEYINPUT11), .B(KEYINPUT96), .ZN(n439) );
  XOR2_X1 U453 ( .A(KEYINPUT97), .B(KEYINPUT95), .Z(n438) );
  INV_X1 U454 ( .A(n653), .ZN(n422) );
  INV_X1 U455 ( .A(KEYINPUT0), .ZN(n403) );
  NAND2_X1 U456 ( .A1(n402), .A2(n400), .ZN(n397) );
  NOR2_X1 U457 ( .A1(n401), .A2(KEYINPUT0), .ZN(n400) );
  INV_X1 U458 ( .A(n405), .ZN(n401) );
  XNOR2_X1 U459 ( .A(n516), .B(n430), .ZN(n625) );
  XNOR2_X1 U460 ( .A(n512), .B(n506), .ZN(n430) );
  XNOR2_X1 U461 ( .A(n392), .B(G119), .ZN(n510) );
  XNOR2_X1 U462 ( .A(G113), .B(KEYINPUT3), .ZN(n392) );
  XNOR2_X1 U463 ( .A(G902), .B(KEYINPUT15), .ZN(n434) );
  NOR2_X1 U464 ( .A1(n740), .A2(n722), .ZN(n686) );
  XNOR2_X1 U465 ( .A(n516), .B(n431), .ZN(n700) );
  XNOR2_X1 U466 ( .A(n432), .B(n520), .ZN(n431) );
  XNOR2_X1 U467 ( .A(n515), .B(n517), .ZN(n432) );
  NAND2_X1 U468 ( .A1(G234), .A2(G237), .ZN(n480) );
  NOR2_X1 U469 ( .A1(n380), .A2(n379), .ZN(n618) );
  NAND2_X1 U470 ( .A1(n383), .A2(n384), .ZN(n379) );
  AND2_X1 U471 ( .A1(n534), .A2(n665), .ZN(n427) );
  XNOR2_X1 U472 ( .A(n583), .B(n479), .ZN(n607) );
  INV_X1 U473 ( .A(KEYINPUT19), .ZN(n479) );
  NAND2_X1 U474 ( .A1(n665), .A2(n545), .ZN(n561) );
  INV_X1 U475 ( .A(n595), .ZN(n670) );
  XNOR2_X1 U476 ( .A(n492), .B(n374), .ZN(n495) );
  XNOR2_X1 U477 ( .A(n458), .B(n457), .ZN(n714) );
  XNOR2_X1 U478 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U479 ( .A(n413), .B(n411), .ZN(n458) );
  XNOR2_X1 U480 ( .A(n446), .B(n445), .ZN(n708) );
  XNOR2_X1 U481 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U482 ( .A(G113), .B(G143), .ZN(n443) );
  XNOR2_X1 U483 ( .A(n728), .B(n425), .ZN(n620) );
  XNOR2_X1 U484 ( .A(n470), .B(n473), .ZN(n425) );
  NOR2_X1 U485 ( .A1(G952), .A2(n742), .ZN(n721) );
  NAND2_X1 U486 ( .A1(n358), .A2(n365), .ZN(n604) );
  XNOR2_X1 U487 ( .A(n373), .B(KEYINPUT40), .ZN(n753) );
  NAND2_X1 U488 ( .A1(n360), .A2(n365), .ZN(n373) );
  NOR2_X1 U489 ( .A1(n367), .A2(n603), .ZN(n366) );
  XNOR2_X1 U490 ( .A(KEYINPUT107), .B(n587), .ZN(n746) );
  XNOR2_X1 U491 ( .A(n538), .B(n537), .ZN(n749) );
  XNOR2_X1 U492 ( .A(n536), .B(KEYINPUT74), .ZN(n537) );
  INV_X1 U493 ( .A(KEYINPUT32), .ZN(n536) );
  XNOR2_X1 U494 ( .A(n603), .B(KEYINPUT101), .ZN(n647) );
  OR2_X1 U495 ( .A1(n395), .A2(n394), .ZN(n632) );
  OR2_X1 U496 ( .A1(n664), .A2(n667), .ZN(n394) );
  XNOR2_X1 U497 ( .A(n553), .B(n396), .ZN(n395) );
  INV_X1 U498 ( .A(KEYINPUT80), .ZN(n396) );
  AND2_X1 U499 ( .A1(n357), .A2(n397), .ZN(n352) );
  OR2_X1 U500 ( .A1(n612), .A2(n552), .ZN(n353) );
  XOR2_X1 U501 ( .A(KEYINPUT75), .B(n574), .Z(n354) );
  AND2_X1 U502 ( .A1(n632), .A2(n353), .ZN(n355) );
  AND2_X1 U503 ( .A1(n609), .A2(KEYINPUT47), .ZN(n356) );
  AND2_X1 U504 ( .A1(n404), .A2(n398), .ZN(n357) );
  AND2_X1 U505 ( .A1(n371), .A2(n370), .ZN(n358) );
  AND2_X1 U506 ( .A1(n410), .A2(n577), .ZN(n359) );
  AND2_X1 U507 ( .A1(n371), .A2(n366), .ZN(n360) );
  OR2_X1 U508 ( .A1(n405), .A2(n403), .ZN(n361) );
  AND2_X1 U509 ( .A1(n404), .A2(n361), .ZN(n362) );
  XOR2_X1 U510 ( .A(n527), .B(n526), .Z(n363) );
  XOR2_X1 U511 ( .A(KEYINPUT48), .B(KEYINPUT79), .Z(n364) );
  XNOR2_X1 U512 ( .A(n426), .B(n464), .ZN(n728) );
  XNOR2_X1 U513 ( .A(n503), .B(n502), .ZN(n733) );
  INV_X1 U514 ( .A(n370), .ZN(n367) );
  INV_X1 U515 ( .A(n589), .ZN(n369) );
  NAND2_X1 U516 ( .A1(n589), .A2(n372), .ZN(n371) );
  NOR2_X1 U517 ( .A1(n719), .A2(G902), .ZN(n376) );
  NAND2_X1 U518 ( .A1(n389), .A2(n423), .ZN(n391) );
  NAND2_X1 U519 ( .A1(n558), .A2(KEYINPUT44), .ZN(n390) );
  NAND2_X1 U520 ( .A1(n362), .A2(n397), .ZN(n549) );
  NOR2_X1 U521 ( .A1(n668), .A2(n399), .ZN(n398) );
  INV_X1 U522 ( .A(n361), .ZN(n399) );
  INV_X1 U523 ( .A(n607), .ZN(n402) );
  NAND2_X1 U524 ( .A1(n607), .A2(KEYINPUT0), .ZN(n404) );
  NAND2_X1 U525 ( .A1(n407), .A2(n618), .ZN(n687) );
  NOR2_X1 U526 ( .A1(n722), .A2(n354), .ZN(n407) );
  INV_X1 U527 ( .A(n582), .ZN(n581) );
  INV_X1 U528 ( .A(n596), .ZN(n410) );
  NOR2_X1 U529 ( .A1(n656), .A2(n422), .ZN(n417) );
  NAND2_X1 U530 ( .A1(n654), .A2(n417), .ZN(n416) );
  INV_X1 U531 ( .A(n592), .ZN(n654) );
  NAND2_X1 U532 ( .A1(n654), .A2(n653), .ZN(n658) );
  NAND2_X1 U533 ( .A1(n654), .A2(n419), .ZN(n418) );
  NOR2_X1 U534 ( .A1(n656), .A2(n420), .ZN(n419) );
  NAND2_X1 U535 ( .A1(n653), .A2(n594), .ZN(n420) );
  NAND2_X1 U536 ( .A1(n529), .A2(n424), .ZN(n423) );
  XNOR2_X2 U537 ( .A(n428), .B(n363), .ZN(n750) );
  NAND2_X1 U538 ( .A1(n525), .A2(n429), .ZN(n428) );
  INV_X1 U539 ( .A(n588), .ZN(n429) );
  NOR2_X1 U540 ( .A1(n623), .A2(n721), .ZN(n624) );
  BUF_X1 U541 ( .A(n560), .Z(n590) );
  NOR2_X1 U542 ( .A1(n610), .A2(n356), .ZN(n611) );
  XNOR2_X1 U543 ( .A(n606), .B(n605), .ZN(n610) );
  XNOR2_X2 U544 ( .A(n522), .B(n521), .ZN(n600) );
  AND2_X1 U545 ( .A1(n746), .A2(n644), .ZN(n433) );
  XNOR2_X1 U546 ( .A(n483), .B(KEYINPUT86), .ZN(n484) );
  XNOR2_X1 U547 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U548 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U549 ( .A(n598), .B(n597), .ZN(n599) );
  INV_X1 U550 ( .A(KEYINPUT35), .ZN(n526) );
  XNOR2_X1 U551 ( .A(n714), .B(n713), .ZN(n715) );
  XNOR2_X1 U552 ( .A(n716), .B(n715), .ZN(n717) );
  XNOR2_X1 U553 ( .A(n434), .B(KEYINPUT83), .ZN(n617) );
  XOR2_X1 U554 ( .A(G122), .B(G104), .Z(n461) );
  NAND2_X1 U555 ( .A1(G214), .A2(n507), .ZN(n435) );
  XOR2_X1 U556 ( .A(n435), .B(n488), .Z(n436) );
  XOR2_X1 U557 ( .A(n461), .B(n436), .Z(n446) );
  XNOR2_X1 U558 ( .A(n438), .B(n437), .ZN(n442) );
  XNOR2_X1 U559 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U560 ( .A(n442), .B(n441), .Z(n444) );
  NOR2_X1 U561 ( .A1(G902), .A2(n708), .ZN(n448) );
  XNOR2_X1 U562 ( .A(KEYINPUT13), .B(G475), .ZN(n447) );
  XOR2_X1 U563 ( .A(KEYINPUT9), .B(KEYINPUT99), .Z(n450) );
  NAND2_X1 U564 ( .A1(G234), .A2(n742), .ZN(n449) );
  XOR2_X1 U565 ( .A(G116), .B(G107), .Z(n462) );
  XNOR2_X1 U566 ( .A(G122), .B(n462), .ZN(n456) );
  INV_X1 U567 ( .A(G128), .ZN(n451) );
  NAND2_X1 U568 ( .A1(G143), .A2(n451), .ZN(n454) );
  INV_X1 U569 ( .A(G143), .ZN(n452) );
  NAND2_X1 U570 ( .A1(n452), .A2(G128), .ZN(n453) );
  INV_X1 U571 ( .A(n503), .ZN(n455) );
  NOR2_X1 U572 ( .A1(G902), .A2(n714), .ZN(n459) );
  INV_X1 U573 ( .A(n543), .ZN(n530) );
  NAND2_X1 U574 ( .A1(n542), .A2(n530), .ZN(n588) );
  NOR2_X1 U575 ( .A1(G898), .A2(n742), .ZN(n730) );
  NAND2_X1 U576 ( .A1(n730), .A2(G902), .ZN(n460) );
  NAND2_X1 U577 ( .A1(G952), .A2(n742), .ZN(n565) );
  NAND2_X1 U578 ( .A1(n460), .A2(n565), .ZN(n481) );
  XOR2_X1 U579 ( .A(n462), .B(n461), .Z(n464) );
  XNOR2_X1 U580 ( .A(KEYINPUT68), .B(KEYINPUT16), .ZN(n463) );
  XNOR2_X1 U581 ( .A(KEYINPUT82), .B(KEYINPUT18), .ZN(n465) );
  XOR2_X1 U582 ( .A(n466), .B(n465), .Z(n469) );
  XNOR2_X1 U583 ( .A(n472), .B(n471), .ZN(n473) );
  NOR2_X1 U584 ( .A1(n620), .A2(n617), .ZN(n477) );
  XOR2_X1 U585 ( .A(KEYINPUT70), .B(n474), .Z(n478) );
  NAND2_X1 U586 ( .A1(n478), .A2(G210), .ZN(n475) );
  XNOR2_X1 U587 ( .A(n475), .B(KEYINPUT84), .ZN(n476) );
  XNOR2_X1 U588 ( .A(n477), .B(n476), .ZN(n560) );
  NAND2_X1 U589 ( .A1(n478), .A2(G214), .ZN(n653) );
  NAND2_X1 U590 ( .A1(n560), .A2(n653), .ZN(n583) );
  XOR2_X1 U591 ( .A(KEYINPUT14), .B(n480), .Z(n683) );
  XOR2_X1 U592 ( .A(KEYINPUT88), .B(KEYINPUT25), .Z(n487) );
  INV_X1 U593 ( .A(n617), .ZN(n482) );
  NAND2_X1 U594 ( .A1(G234), .A2(n482), .ZN(n485) );
  NAND2_X1 U595 ( .A1(G217), .A2(n498), .ZN(n486) );
  XNOR2_X1 U596 ( .A(n487), .B(n486), .ZN(n497) );
  INV_X1 U597 ( .A(n518), .ZN(n489) );
  XNOR2_X1 U598 ( .A(n489), .B(n488), .ZN(n734) );
  XNOR2_X1 U599 ( .A(n490), .B(KEYINPUT71), .ZN(n492) );
  NAND2_X1 U600 ( .A1(G221), .A2(n493), .ZN(n494) );
  XNOR2_X1 U601 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U602 ( .A(n734), .B(n496), .ZN(n719) );
  XOR2_X1 U603 ( .A(KEYINPUT90), .B(KEYINPUT21), .Z(n500) );
  NAND2_X1 U604 ( .A1(G221), .A2(n498), .ZN(n499) );
  XNOR2_X1 U605 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U606 ( .A(KEYINPUT89), .B(n501), .ZN(n668) );
  XOR2_X1 U607 ( .A(KEYINPUT92), .B(G137), .Z(n505) );
  XNOR2_X1 U608 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U609 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n509) );
  NAND2_X1 U610 ( .A1(n507), .A2(G210), .ZN(n508) );
  XNOR2_X1 U611 ( .A(n509), .B(n508), .ZN(n511) );
  NOR2_X1 U612 ( .A1(n625), .A2(G902), .ZN(n513) );
  XNOR2_X1 U613 ( .A(G104), .B(G107), .ZN(n519) );
  XNOR2_X1 U614 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U615 ( .A(KEYINPUT66), .B(G469), .ZN(n521) );
  XOR2_X1 U616 ( .A(n600), .B(KEYINPUT1), .Z(n534) );
  NOR2_X1 U617 ( .A1(n549), .A2(n691), .ZN(n524) );
  XNOR2_X1 U618 ( .A(n524), .B(KEYINPUT34), .ZN(n525) );
  INV_X1 U619 ( .A(KEYINPUT78), .ZN(n527) );
  XNOR2_X1 U620 ( .A(n555), .B(KEYINPUT65), .ZN(n529) );
  INV_X1 U621 ( .A(KEYINPUT44), .ZN(n528) );
  NOR2_X1 U622 ( .A1(n542), .A2(n530), .ZN(n593) );
  NAND2_X1 U623 ( .A1(n593), .A2(n352), .ZN(n533) );
  INV_X1 U624 ( .A(KEYINPUT22), .ZN(n531) );
  BUF_X1 U625 ( .A(n534), .Z(n664) );
  INV_X1 U626 ( .A(n664), .ZN(n586) );
  INV_X1 U627 ( .A(n667), .ZN(n554) );
  NOR2_X1 U628 ( .A1(n586), .A2(n554), .ZN(n535) );
  NAND2_X1 U629 ( .A1(n553), .A2(n535), .ZN(n538) );
  NOR2_X1 U630 ( .A1(n664), .A2(n539), .ZN(n540) );
  NAND2_X1 U631 ( .A1(n540), .A2(n667), .ZN(n541) );
  NOR2_X1 U632 ( .A1(n670), .A2(n541), .ZN(n639) );
  NAND2_X1 U633 ( .A1(n542), .A2(n543), .ZN(n603) );
  NOR2_X1 U634 ( .A1(n543), .A2(n542), .ZN(n649) );
  INV_X1 U635 ( .A(n649), .ZN(n572) );
  NAND2_X1 U636 ( .A1(n603), .A2(n572), .ZN(n544) );
  XNOR2_X1 U637 ( .A(n544), .B(KEYINPUT100), .ZN(n657) );
  XNOR2_X1 U638 ( .A(n657), .B(KEYINPUT77), .ZN(n612) );
  INV_X1 U639 ( .A(n600), .ZN(n545) );
  NOR2_X1 U640 ( .A1(n549), .A2(n561), .ZN(n546) );
  XNOR2_X1 U641 ( .A(n546), .B(KEYINPUT91), .ZN(n547) );
  NOR2_X1 U642 ( .A1(n670), .A2(n547), .ZN(n634) );
  AND2_X1 U643 ( .A1(n665), .A2(n664), .ZN(n548) );
  NAND2_X1 U644 ( .A1(n670), .A2(n548), .ZN(n675) );
  NOR2_X1 U645 ( .A1(n549), .A2(n675), .ZN(n551) );
  XOR2_X1 U646 ( .A(KEYINPUT31), .B(KEYINPUT94), .Z(n550) );
  XNOR2_X1 U647 ( .A(n551), .B(n550), .ZN(n650) );
  NOR2_X1 U648 ( .A1(n634), .A2(n650), .ZN(n552) );
  NAND2_X1 U649 ( .A1(n557), .A2(n556), .ZN(n558) );
  INV_X1 U650 ( .A(KEYINPUT45), .ZN(n559) );
  XNOR2_X1 U651 ( .A(KEYINPUT38), .B(n590), .ZN(n592) );
  XNOR2_X1 U652 ( .A(KEYINPUT103), .B(n561), .ZN(n571) );
  NAND2_X1 U653 ( .A1(G953), .A2(G902), .ZN(n562) );
  NOR2_X1 U654 ( .A1(n683), .A2(n562), .ZN(n563) );
  XOR2_X1 U655 ( .A(KEYINPUT102), .B(n563), .Z(n564) );
  NOR2_X1 U656 ( .A1(G900), .A2(n564), .ZN(n567) );
  NOR2_X1 U657 ( .A1(n683), .A2(n565), .ZN(n566) );
  NOR2_X1 U658 ( .A1(n567), .A2(n566), .ZN(n575) );
  NAND2_X1 U659 ( .A1(n670), .A2(n653), .ZN(n568) );
  XNOR2_X1 U660 ( .A(KEYINPUT30), .B(n568), .ZN(n569) );
  NOR2_X1 U661 ( .A1(n575), .A2(n569), .ZN(n570) );
  NAND2_X1 U662 ( .A1(n571), .A2(n570), .ZN(n589) );
  OR2_X1 U663 ( .A1(n572), .A2(n604), .ZN(n573) );
  XNOR2_X1 U664 ( .A(n573), .B(KEYINPUT108), .ZN(n754) );
  NAND2_X1 U665 ( .A1(KEYINPUT2), .A2(n754), .ZN(n574) );
  NOR2_X1 U666 ( .A1(n575), .A2(n668), .ZN(n576) );
  NAND2_X1 U667 ( .A1(n576), .A2(n667), .ZN(n596) );
  NAND2_X1 U668 ( .A1(n581), .A2(n653), .ZN(n578) );
  NOR2_X1 U669 ( .A1(n664), .A2(n578), .ZN(n579) );
  XNOR2_X1 U670 ( .A(n579), .B(KEYINPUT43), .ZN(n580) );
  NOR2_X1 U671 ( .A1(n590), .A2(n580), .ZN(n652) );
  NOR2_X1 U672 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U673 ( .A(KEYINPUT36), .B(n584), .Z(n585) );
  NOR2_X1 U674 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U675 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U676 ( .A1(n591), .A2(n590), .ZN(n644) );
  INV_X1 U677 ( .A(n593), .ZN(n656) );
  XNOR2_X1 U678 ( .A(KEYINPUT41), .B(KEYINPUT106), .ZN(n594) );
  OR2_X1 U679 ( .A1(n596), .A2(n595), .ZN(n598) );
  NOR2_X1 U680 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U681 ( .A(KEYINPUT105), .B(n601), .ZN(n608) );
  XOR2_X1 U682 ( .A(KEYINPUT42), .B(n602), .Z(n752) );
  NAND2_X1 U683 ( .A1(n752), .A2(n753), .ZN(n606) );
  NOR2_X1 U684 ( .A1(n608), .A2(n607), .ZN(n645) );
  NAND2_X1 U685 ( .A1(n657), .A2(n645), .ZN(n609) );
  NAND2_X1 U686 ( .A1(n433), .A2(n611), .ZN(n616) );
  NOR2_X1 U687 ( .A1(KEYINPUT47), .A2(n612), .ZN(n613) );
  NAND2_X1 U688 ( .A1(n613), .A2(n645), .ZN(n614) );
  XNOR2_X1 U689 ( .A(KEYINPUT69), .B(n614), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n706), .A2(G210), .ZN(n622) );
  XOR2_X1 U691 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n619) );
  XNOR2_X1 U692 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U693 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U694 ( .A(n624), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U695 ( .A(n625), .B(KEYINPUT62), .ZN(n627) );
  NAND2_X1 U696 ( .A1(n706), .A2(G472), .ZN(n626) );
  XNOR2_X1 U697 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U698 ( .A(KEYINPUT63), .B(KEYINPUT81), .ZN(n629) );
  XNOR2_X1 U699 ( .A(n630), .B(n629), .ZN(G57) );
  XOR2_X1 U700 ( .A(G101), .B(KEYINPUT109), .Z(n631) );
  XNOR2_X1 U701 ( .A(n632), .B(n631), .ZN(G3) );
  NAND2_X1 U702 ( .A1(n634), .A2(n647), .ZN(n633) );
  XNOR2_X1 U703 ( .A(n633), .B(G104), .ZN(G6) );
  XNOR2_X1 U704 ( .A(G107), .B(KEYINPUT27), .ZN(n638) );
  XOR2_X1 U705 ( .A(KEYINPUT110), .B(KEYINPUT26), .Z(n636) );
  NAND2_X1 U706 ( .A1(n634), .A2(n649), .ZN(n635) );
  XNOR2_X1 U707 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U708 ( .A(n638), .B(n637), .ZN(G9) );
  XOR2_X1 U709 ( .A(G110), .B(n639), .Z(G12) );
  XOR2_X1 U710 ( .A(KEYINPUT29), .B(KEYINPUT112), .Z(n641) );
  NAND2_X1 U711 ( .A1(n645), .A2(n649), .ZN(n640) );
  XNOR2_X1 U712 ( .A(n641), .B(n640), .ZN(n643) );
  XOR2_X1 U713 ( .A(G128), .B(KEYINPUT111), .Z(n642) );
  XNOR2_X1 U714 ( .A(n643), .B(n642), .ZN(G30) );
  XNOR2_X1 U715 ( .A(G143), .B(n644), .ZN(G45) );
  NAND2_X1 U716 ( .A1(n647), .A2(n645), .ZN(n646) );
  XNOR2_X1 U717 ( .A(n646), .B(G146), .ZN(G48) );
  NAND2_X1 U718 ( .A1(n650), .A2(n647), .ZN(n648) );
  XNOR2_X1 U719 ( .A(n648), .B(G113), .ZN(G15) );
  NAND2_X1 U720 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U721 ( .A(n651), .B(G116), .ZN(G18) );
  XOR2_X1 U722 ( .A(G140), .B(n652), .Z(G42) );
  XOR2_X1 U723 ( .A(KEYINPUT116), .B(KEYINPUT53), .Z(n697) );
  NOR2_X1 U724 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U725 ( .A1(n656), .A2(n655), .ZN(n661) );
  INV_X1 U726 ( .A(n657), .ZN(n659) );
  NOR2_X1 U727 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U728 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U729 ( .A1(n662), .A2(n691), .ZN(n663) );
  XOR2_X1 U730 ( .A(KEYINPUT115), .B(n663), .Z(n680) );
  NOR2_X1 U731 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U732 ( .A(KEYINPUT50), .B(n666), .Z(n673) );
  NAND2_X1 U733 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U734 ( .A(n669), .B(KEYINPUT49), .ZN(n671) );
  NOR2_X1 U735 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U736 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U737 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U738 ( .A(KEYINPUT51), .B(n676), .ZN(n677) );
  NOR2_X1 U739 ( .A1(n692), .A2(n677), .ZN(n678) );
  XNOR2_X1 U740 ( .A(KEYINPUT114), .B(n678), .ZN(n679) );
  NOR2_X1 U741 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U742 ( .A(n681), .B(KEYINPUT52), .ZN(n682) );
  NOR2_X1 U743 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U744 ( .A1(G952), .A2(n684), .ZN(n690) );
  XNOR2_X1 U745 ( .A(KEYINPUT2), .B(KEYINPUT76), .ZN(n685) );
  OR2_X1 U746 ( .A1(n686), .A2(n685), .ZN(n688) );
  NAND2_X1 U747 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U748 ( .A1(n690), .A2(n689), .ZN(n694) );
  NOR2_X1 U749 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U750 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U751 ( .A1(n695), .A2(n742), .ZN(n696) );
  XNOR2_X1 U752 ( .A(n697), .B(n696), .ZN(G75) );
  XNOR2_X1 U753 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n698) );
  XNOR2_X1 U754 ( .A(n698), .B(KEYINPUT117), .ZN(n699) );
  XNOR2_X1 U755 ( .A(KEYINPUT57), .B(n699), .ZN(n702) );
  XNOR2_X1 U756 ( .A(n700), .B(KEYINPUT58), .ZN(n701) );
  XNOR2_X1 U757 ( .A(n702), .B(n701), .ZN(n704) );
  NAND2_X1 U758 ( .A1(n706), .A2(G469), .ZN(n703) );
  XOR2_X1 U759 ( .A(n704), .B(n703), .Z(n705) );
  NOR2_X1 U760 ( .A1(n721), .A2(n705), .ZN(G54) );
  NAND2_X1 U761 ( .A1(n706), .A2(G475), .ZN(n710) );
  XOR2_X1 U762 ( .A(KEYINPUT120), .B(KEYINPUT59), .Z(n707) );
  XNOR2_X1 U763 ( .A(n708), .B(n707), .ZN(n709) );
  XNOR2_X1 U764 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X2 U765 ( .A1(n721), .A2(n711), .ZN(n712) );
  XNOR2_X1 U766 ( .A(KEYINPUT60), .B(n712), .ZN(G60) );
  NAND2_X1 U767 ( .A1(n706), .A2(G478), .ZN(n716) );
  INV_X1 U768 ( .A(KEYINPUT121), .ZN(n713) );
  NOR2_X1 U769 ( .A1(n721), .A2(n717), .ZN(G63) );
  NAND2_X1 U770 ( .A1(G217), .A2(n706), .ZN(n718) );
  XNOR2_X1 U771 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U772 ( .A1(n721), .A2(n720), .ZN(G66) );
  OR2_X1 U773 ( .A1(G953), .A2(n722), .ZN(n727) );
  NAND2_X1 U774 ( .A1(G224), .A2(G953), .ZN(n723) );
  XNOR2_X1 U775 ( .A(n723), .B(KEYINPUT61), .ZN(n724) );
  XNOR2_X1 U776 ( .A(KEYINPUT122), .B(n724), .ZN(n725) );
  NAND2_X1 U777 ( .A1(n725), .A2(G898), .ZN(n726) );
  NAND2_X1 U778 ( .A1(n727), .A2(n726), .ZN(n732) );
  XOR2_X1 U779 ( .A(n728), .B(KEYINPUT123), .Z(n729) );
  NOR2_X1 U780 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U781 ( .A(n732), .B(n731), .ZN(G69) );
  XOR2_X1 U782 ( .A(n734), .B(KEYINPUT124), .Z(n735) );
  XOR2_X1 U783 ( .A(n733), .B(n735), .Z(n741) );
  XOR2_X1 U784 ( .A(n741), .B(KEYINPUT125), .Z(n736) );
  XNOR2_X1 U785 ( .A(G227), .B(n736), .ZN(n737) );
  NAND2_X1 U786 ( .A1(G900), .A2(n737), .ZN(n738) );
  NAND2_X1 U787 ( .A1(G953), .A2(n738), .ZN(n739) );
  XNOR2_X1 U788 ( .A(n739), .B(KEYINPUT126), .ZN(n745) );
  XNOR2_X1 U789 ( .A(n741), .B(n740), .ZN(n743) );
  NAND2_X1 U790 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U791 ( .A1(n745), .A2(n744), .ZN(G72) );
  XNOR2_X1 U792 ( .A(KEYINPUT37), .B(KEYINPUT113), .ZN(n747) );
  XNOR2_X1 U793 ( .A(n747), .B(n746), .ZN(n748) );
  XNOR2_X1 U794 ( .A(G125), .B(n748), .ZN(G27) );
  XOR2_X1 U795 ( .A(n749), .B(G119), .Z(G21) );
  XNOR2_X1 U796 ( .A(G122), .B(KEYINPUT127), .ZN(n751) );
  XOR2_X1 U797 ( .A(n751), .B(n750), .Z(G24) );
  XNOR2_X1 U798 ( .A(G137), .B(n752), .ZN(G39) );
  XNOR2_X1 U799 ( .A(G131), .B(n753), .ZN(G33) );
  XNOR2_X1 U800 ( .A(G134), .B(n754), .ZN(G36) );
endmodule

