//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n187));
  INV_X1    g001(.A(G469), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G137), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT11), .A3(G134), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(G137), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G131), .ZN(new_n196));
  INV_X1    g010(.A(G131), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n191), .A2(new_n193), .A3(new_n197), .A4(new_n194), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G107), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G104), .ZN(new_n201));
  AND2_X1   g015(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n202));
  NOR2_X1   g016(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n201), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G101), .ZN(new_n205));
  INV_X1    g019(.A(G104), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G107), .ZN(new_n207));
  NAND2_X1  g021(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(G104), .A3(new_n200), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n204), .A2(new_n205), .A3(new_n207), .A4(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n201), .A2(new_n207), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G101), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(G146), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT64), .B1(new_n216), .B2(G143), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(new_n214), .A3(G146), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n215), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT1), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(G128), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n216), .A2(G143), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n214), .A2(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n226), .B(KEYINPUT1), .C1(new_n214), .C2(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G128), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n226), .B1(new_n223), .B2(KEYINPUT1), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n225), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n213), .A2(new_n222), .A3(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n223), .A2(KEYINPUT79), .A3(KEYINPUT1), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G128), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n221), .B1(G143), .B2(new_n216), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n234), .A2(KEYINPUT79), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n217), .A2(new_n219), .ZN(new_n236));
  OAI22_X1  g050(.A1(new_n233), .A2(new_n235), .B1(new_n236), .B2(new_n215), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n213), .B1(new_n222), .B2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n199), .B1(new_n231), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT12), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI211_X1 g055(.A(KEYINPUT12), .B(new_n199), .C1(new_n231), .C2(new_n238), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  OR2_X1    g057(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n244), .A2(new_n208), .B1(G104), .B2(new_n200), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n209), .A2(new_n207), .ZN(new_n246));
  OAI21_X1  g060(.A(G101), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n247), .A2(KEYINPUT4), .A3(new_n210), .ZN(new_n248));
  AND2_X1   g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  NOR2_X1   g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n220), .A2(new_n249), .B1(new_n225), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n253), .B(G101), .C1(new_n245), .C2(new_n246), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT78), .B1(new_n248), .B2(new_n255), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n252), .A2(new_n254), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT78), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n247), .A2(KEYINPUT4), .A3(new_n210), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT80), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n210), .A2(new_n262), .A3(new_n212), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n262), .B1(new_n210), .B2(new_n212), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT10), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n266), .B1(new_n222), .B2(new_n230), .ZN(new_n267));
  INV_X1    g081(.A(G128), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n268), .B1(new_n234), .B2(KEYINPUT79), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT79), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(new_n215), .B2(new_n221), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n220), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n221), .A2(G128), .ZN(new_n273));
  AOI211_X1 g087(.A(new_n273), .B(new_n215), .C1(new_n217), .C2(new_n219), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n210), .B(new_n212), .C1(new_n272), .C2(new_n274), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n265), .A2(new_n267), .B1(new_n275), .B2(new_n266), .ZN(new_n276));
  INV_X1    g090(.A(new_n199), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n261), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n243), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G953), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT69), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT69), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G953), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G227), .ZN(new_n285));
  XOR2_X1   g099(.A(G110), .B(G140), .Z(new_n286));
  XNOR2_X1  g100(.A(new_n285), .B(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n279), .A2(new_n287), .ZN(new_n288));
  NOR3_X1   g102(.A1(new_n248), .A2(new_n255), .A3(KEYINPUT78), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n258), .B1(new_n257), .B2(new_n259), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n213), .A2(KEYINPUT80), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n210), .A2(new_n262), .A3(new_n212), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n267), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n294), .B1(KEYINPUT10), .B2(new_n238), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n199), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n287), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(new_n278), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n288), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G902), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n188), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n243), .A2(new_n278), .A3(new_n297), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n297), .B1(new_n296), .B2(new_n278), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n188), .B(new_n300), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT81), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n261), .A2(new_n276), .A3(new_n277), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n277), .B1(new_n261), .B2(new_n276), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n287), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(G902), .B1(new_n310), .B2(new_n302), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(KEYINPUT81), .A3(new_n188), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n301), .B1(new_n307), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT9), .B(G234), .ZN(new_n314));
  OAI21_X1  g128(.A(G221), .B1(new_n314), .B2(G902), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n187), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n308), .A2(new_n287), .ZN(new_n318));
  AOI22_X1  g132(.A1(new_n318), .A2(new_n296), .B1(new_n279), .B2(new_n287), .ZN(new_n319));
  OAI21_X1  g133(.A(G469), .B1(new_n319), .B2(G902), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n310), .A2(new_n302), .ZN(new_n321));
  AND4_X1   g135(.A1(KEYINPUT81), .A2(new_n321), .A3(new_n188), .A4(new_n300), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT81), .B1(new_n311), .B2(new_n188), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(KEYINPUT82), .A3(new_n315), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n317), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT23), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT66), .B(G119), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n327), .B1(new_n328), .B2(G128), .ZN(new_n329));
  INV_X1    g143(.A(G119), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n268), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n331), .B1(new_n328), .B2(new_n268), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n329), .B1(new_n332), .B2(new_n327), .ZN(new_n333));
  XOR2_X1   g147(.A(KEYINPUT24), .B(G110), .Z(new_n334));
  OAI22_X1  g148(.A1(new_n333), .A2(G110), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(G125), .B(G140), .ZN(new_n336));
  OR2_X1    g150(.A1(new_n336), .A2(KEYINPUT72), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(KEYINPUT72), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n216), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT16), .ZN(new_n340));
  INV_X1    g154(.A(G140), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(G125), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(G125), .ZN(new_n343));
  INV_X1    g157(.A(G125), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G140), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g160(.A(G146), .B(new_n342), .C1(new_n346), .C2(new_n340), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n339), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n335), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n342), .B1(new_n346), .B2(new_n340), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n216), .ZN(new_n351));
  AOI22_X1  g165(.A1(new_n351), .A2(new_n347), .B1(new_n332), .B2(new_n334), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n333), .A2(G110), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT73), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n284), .A2(G221), .A3(G234), .ZN(new_n357));
  XNOR2_X1  g171(.A(KEYINPUT22), .B(G137), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n357), .B(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n355), .A2(new_n356), .A3(new_n360), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n335), .A2(new_n348), .B1(new_n352), .B2(new_n353), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT73), .B1(new_n362), .B2(new_n359), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n349), .A2(new_n354), .A3(new_n359), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT74), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT74), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n362), .A2(new_n367), .A3(new_n359), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n364), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G217), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n371), .B1(G234), .B2(new_n300), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(G902), .ZN(new_n373));
  XOR2_X1   g187(.A(new_n373), .B(KEYINPUT76), .Z(new_n374));
  NOR2_X1   g188(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n364), .A2(new_n369), .A3(new_n300), .ZN(new_n376));
  NOR2_X1   g190(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n377), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n364), .A2(new_n369), .A3(new_n300), .A4(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n378), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n375), .B1(new_n382), .B2(new_n372), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n330), .A2(KEYINPUT66), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT66), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G119), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(new_n387), .A3(G116), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n330), .A2(G116), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(KEYINPUT2), .B(G113), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n392), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(new_n388), .A3(new_n390), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT67), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n391), .A2(KEYINPUT67), .A3(new_n392), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n222), .A2(new_n230), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n190), .A2(G137), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n192), .A2(G134), .ZN(new_n402));
  OAI21_X1  g216(.A(G131), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n198), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n400), .A2(new_n405), .B1(new_n199), .B2(new_n252), .ZN(new_n406));
  OR2_X1    g220(.A1(KEYINPUT68), .A2(KEYINPUT30), .ZN(new_n407));
  NAND2_X1  g221(.A1(KEYINPUT68), .A2(KEYINPUT30), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n199), .A2(new_n252), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n404), .B1(new_n222), .B2(new_n230), .ZN(new_n411));
  OAI211_X1 g225(.A(KEYINPUT68), .B(KEYINPUT30), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n399), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n406), .A2(new_n399), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G237), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n284), .A2(G210), .A3(new_n416), .ZN(new_n417));
  OR2_X1    g231(.A1(new_n417), .A2(KEYINPUT27), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(KEYINPUT27), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT26), .B(G101), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT70), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n418), .A2(new_n419), .A3(new_n421), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT31), .B1(new_n415), .B2(new_n426), .ZN(new_n427));
  NOR4_X1   g241(.A1(new_n413), .A2(KEYINPUT31), .A3(new_n426), .A4(new_n414), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n423), .A2(new_n425), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n414), .A2(KEYINPUT28), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT28), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n398), .B(new_n397), .C1(new_n410), .C2(new_n411), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n406), .A2(new_n399), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n430), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n427), .A2(new_n429), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(G472), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n438), .A3(new_n300), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT32), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT32), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n437), .A2(new_n441), .A3(new_n438), .A4(new_n300), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n431), .A2(new_n435), .ZN(new_n444));
  INV_X1    g258(.A(new_n430), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT29), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n300), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT71), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n413), .A2(new_n414), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n446), .B(new_n447), .C1(new_n450), .C2(new_n445), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT71), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n452), .B(new_n300), .C1(new_n446), .C2(new_n447), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n449), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G472), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n384), .B1(new_n443), .B2(new_n455), .ZN(new_n456));
  XOR2_X1   g270(.A(KEYINPUT94), .B(G475), .Z(new_n457));
  NAND4_X1  g271(.A1(new_n284), .A2(G143), .A3(G214), .A4(new_n416), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n281), .A2(new_n283), .A3(G214), .A4(new_n416), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n214), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G131), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT17), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n458), .A2(new_n197), .A3(new_n460), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT93), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n351), .A2(new_n347), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT93), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n462), .A2(new_n468), .A3(new_n463), .A4(new_n464), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n461), .A2(KEYINPUT17), .A3(G131), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n466), .A2(new_n467), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT91), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n346), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n336), .A2(KEYINPUT91), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n339), .B1(new_n475), .B2(new_n216), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n461), .A2(KEYINPUT18), .A3(G131), .ZN(new_n477));
  NAND2_X1  g291(.A1(KEYINPUT18), .A2(G131), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n458), .A2(new_n460), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n476), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT92), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT92), .A4(new_n479), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n471), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(G113), .B(G122), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(new_n206), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(KEYINPUT95), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n300), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n470), .A2(new_n467), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n491), .B1(KEYINPUT93), .B2(new_n465), .ZN(new_n492));
  AOI22_X1  g306(.A1(new_n492), .A2(new_n469), .B1(new_n482), .B2(new_n483), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(new_n488), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n457), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT20), .ZN(new_n496));
  INV_X1    g310(.A(new_n487), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n462), .A2(new_n464), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n473), .A2(new_n474), .A3(KEYINPUT19), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n336), .B(KEYINPUT72), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n500), .B1(new_n501), .B2(KEYINPUT19), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n347), .B1(new_n502), .B2(G146), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n497), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  AOI22_X1  g319(.A1(new_n485), .A2(new_n487), .B1(new_n484), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(G475), .A2(G902), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n496), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n497), .B1(new_n471), .B2(new_n484), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n504), .B1(new_n482), .B2(new_n483), .ZN(new_n510));
  INV_X1    g324(.A(new_n507), .ZN(new_n511));
  NOR4_X1   g325(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT20), .A4(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n495), .B1(new_n508), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT98), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n314), .A2(new_n371), .A3(G953), .ZN(new_n515));
  XOR2_X1   g329(.A(new_n515), .B(KEYINPUT97), .Z(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  XOR2_X1   g331(.A(G128), .B(G143), .Z(new_n518));
  INV_X1    g332(.A(KEYINPUT96), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(G128), .B(G143), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT96), .ZN(new_n522));
  AOI21_X1  g336(.A(G134), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT13), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(new_n214), .A3(G128), .ZN(new_n526));
  OAI211_X1 g340(.A(G134), .B(new_n526), .C1(new_n518), .C2(new_n525), .ZN(new_n527));
  XNOR2_X1  g341(.A(G116), .B(G122), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(new_n200), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n524), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  XOR2_X1   g344(.A(G116), .B(G122), .Z(new_n531));
  INV_X1    g345(.A(G122), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G116), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n200), .B1(new_n533), .B2(KEYINPUT14), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n531), .B(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n520), .A2(G134), .A3(new_n522), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n536), .B1(new_n538), .B2(new_n523), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n517), .A2(new_n530), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n535), .B1(new_n524), .B2(new_n537), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n529), .A2(new_n527), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(new_n523), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n516), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n300), .ZN(new_n546));
  INV_X1    g360(.A(G478), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n547), .A2(KEYINPUT15), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n545), .B(new_n300), .C1(KEYINPUT15), .C2(new_n547), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n514), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n549), .A2(KEYINPUT98), .A3(new_n551), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G952), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(G953), .ZN(new_n557));
  INV_X1    g371(.A(G234), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n557), .B1(new_n558), .B2(new_n416), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  AOI211_X1 g374(.A(new_n300), .B(new_n284), .C1(G234), .C2(G237), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT21), .B(G898), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n513), .A2(new_n555), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(G214), .B1(G237), .B2(G902), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  XOR2_X1   g380(.A(G110), .B(G122), .Z(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(KEYINPUT83), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n397), .A2(new_n259), .A3(new_n398), .A4(new_n254), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT5), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n385), .A2(new_n387), .A3(new_n570), .A4(G116), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n571), .A2(G113), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n388), .A2(KEYINPUT5), .A3(new_n390), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n389), .B1(new_n328), .B2(G116), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n572), .A2(new_n573), .B1(new_n574), .B2(new_n394), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n292), .A2(new_n575), .A3(new_n293), .ZN(new_n576));
  AOI211_X1 g390(.A(KEYINPUT6), .B(new_n568), .C1(new_n569), .C2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n569), .A2(new_n576), .A3(new_n568), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT84), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n569), .A2(new_n576), .A3(KEYINPUT84), .A4(new_n568), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n568), .B1(new_n569), .B2(new_n576), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT6), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n577), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  OR3_X1    g400(.A1(new_n252), .A2(KEYINPUT85), .A3(new_n344), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT85), .B1(new_n252), .B2(new_n344), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n222), .A2(new_n230), .A3(new_n344), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(KEYINPUT86), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n592), .A2(G224), .A3(new_n280), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n280), .A2(G224), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n589), .A2(new_n594), .A3(new_n591), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n586), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n594), .A2(KEYINPUT7), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT86), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n590), .B(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n589), .B1(new_n600), .B2(KEYINPUT88), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT88), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n591), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n598), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n598), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n589), .A2(new_n591), .A3(KEYINPUT89), .A4(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT89), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n587), .A2(new_n605), .A3(new_n588), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n607), .B1(new_n600), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n575), .A2(new_n213), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n568), .B(KEYINPUT8), .ZN(new_n612));
  INV_X1    g426(.A(new_n572), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n613), .B1(new_n573), .B2(KEYINPUT87), .ZN(new_n614));
  OR2_X1    g428(.A1(new_n573), .A2(KEYINPUT87), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n614), .A2(new_n615), .B1(new_n574), .B2(new_n394), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n611), .B(new_n612), .C1(new_n616), .C2(new_n213), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n604), .A2(new_n610), .A3(new_n582), .A4(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n597), .A2(new_n300), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(G210), .B1(G237), .B2(G902), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(G902), .B1(new_n586), .B2(new_n596), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(new_n618), .A3(new_n620), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n566), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n625), .A2(KEYINPUT90), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT90), .ZN(new_n627));
  AOI211_X1 g441(.A(new_n627), .B(new_n566), .C1(new_n622), .C2(new_n624), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n326), .A2(new_n456), .A3(new_n564), .A4(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G101), .ZN(G3));
  NOR3_X1   g445(.A1(new_n413), .A2(new_n414), .A3(new_n426), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT31), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n436), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n634), .A2(new_n428), .ZN(new_n635));
  OAI21_X1  g449(.A(G472), .B1(new_n635), .B2(G902), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n383), .A2(new_n439), .A3(new_n636), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n317), .A2(new_n325), .A3(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n563), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n625), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT99), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n641), .B1(new_n541), .B2(new_n543), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n539), .A2(KEYINPUT99), .A3(new_n530), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n642), .A2(new_n643), .A3(new_n516), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(KEYINPUT100), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT100), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n642), .A2(new_n643), .A3(new_n646), .A4(new_n516), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n540), .A2(KEYINPUT33), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT33), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n545), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n547), .A2(G902), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n650), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n546), .A2(new_n547), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n513), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n640), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n638), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT101), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT34), .B(G104), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G6));
  NAND2_X1  g476(.A1(new_n505), .A2(new_n484), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n663), .B(new_n507), .C1(new_n493), .C2(new_n497), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(KEYINPUT20), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n506), .A2(new_n496), .A3(new_n507), .ZN(new_n666));
  AOI21_X1  g480(.A(G902), .B1(new_n493), .B2(new_n488), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n667), .B1(new_n493), .B2(new_n488), .ZN(new_n668));
  AOI22_X1  g482(.A1(new_n665), .A2(new_n666), .B1(new_n668), .B2(new_n457), .ZN(new_n669));
  AND4_X1   g483(.A1(new_n669), .A2(new_n625), .A3(new_n639), .A4(new_n555), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n638), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT35), .B(G107), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  NOR2_X1   g487(.A1(new_n360), .A2(KEYINPUT36), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n355), .B(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n374), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(new_n382), .B2(new_n372), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  AND4_X1   g493(.A1(new_n439), .A2(new_n564), .A3(new_n636), .A4(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n326), .A2(new_n629), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT37), .B(G110), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT102), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n681), .B(new_n683), .ZN(G12));
  NAND2_X1  g498(.A1(new_n443), .A2(new_n455), .ZN(new_n685));
  AND4_X1   g499(.A1(new_n300), .A2(new_n597), .A3(new_n618), .A4(new_n620), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n620), .B1(new_n623), .B2(new_n618), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n565), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n678), .ZN(new_n689));
  AND4_X1   g503(.A1(new_n685), .A2(new_n689), .A3(new_n317), .A4(new_n325), .ZN(new_n690));
  INV_X1    g504(.A(G900), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n561), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n559), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n669), .A2(new_n555), .A3(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G128), .ZN(G30));
  XNOR2_X1  g511(.A(new_n693), .B(KEYINPUT39), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n326), .A2(new_n698), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n699), .A2(KEYINPUT40), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(KEYINPUT40), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n415), .A2(new_n445), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n433), .A2(new_n434), .ZN(new_n703));
  AOI21_X1  g517(.A(G902), .B1(new_n703), .B2(new_n430), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n438), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(new_n705), .B(KEYINPUT103), .Z(new_n706));
  AOI21_X1  g520(.A(new_n706), .B1(new_n440), .B2(new_n442), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(new_n679), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n622), .A2(new_n624), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT38), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n513), .A2(new_n555), .A3(new_n565), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n700), .A2(new_n701), .A3(new_n708), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G143), .ZN(G45));
  INV_X1    g529(.A(new_n693), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n657), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n690), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G146), .ZN(G48));
  NAND2_X1  g533(.A1(new_n307), .A2(new_n312), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n311), .A2(new_n188), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n720), .A2(new_n315), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n658), .A2(new_n456), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT41), .B(G113), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G15));
  NAND3_X1  g539(.A1(new_n670), .A2(new_n456), .A3(new_n722), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G116), .ZN(G18));
  NAND3_X1  g541(.A1(new_n720), .A2(new_n315), .A3(new_n721), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n688), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n729), .A2(new_n685), .A3(new_n564), .A4(new_n679), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G119), .ZN(G21));
  INV_X1    g545(.A(KEYINPUT104), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n636), .A2(new_n439), .A3(new_n732), .ZN(new_n733));
  OAI211_X1 g547(.A(KEYINPUT104), .B(G472), .C1(new_n635), .C2(G902), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n384), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n712), .B1(new_n622), .B2(new_n624), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n735), .A2(new_n736), .A3(new_n639), .A4(new_n722), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  INV_X1    g552(.A(KEYINPUT105), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n733), .A2(new_n734), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n717), .A3(new_n679), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n722), .A2(new_n625), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n739), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n678), .B1(new_n733), .B2(new_n734), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n729), .A2(new_n744), .A3(KEYINPUT105), .A4(new_n717), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G125), .ZN(G27));
  NAND3_X1  g561(.A1(new_n622), .A2(new_n565), .A3(new_n624), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n748), .A2(new_n313), .A3(new_n316), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n456), .A2(new_n717), .A3(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT42), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n456), .A2(new_n749), .A3(KEYINPUT42), .A4(new_n717), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G131), .ZN(G33));
  NAND3_X1  g569(.A1(new_n456), .A2(new_n695), .A3(new_n749), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G134), .ZN(G36));
  AOI22_X1  g571(.A1(new_n648), .A2(new_n649), .B1(new_n651), .B2(new_n545), .ZN(new_n758));
  AOI22_X1  g572(.A1(new_n758), .A2(new_n653), .B1(new_n547), .B2(new_n546), .ZN(new_n759));
  OAI21_X1  g573(.A(KEYINPUT43), .B1(new_n513), .B2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n669), .A2(new_n656), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n678), .B1(new_n439), .B2(new_n636), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT44), .ZN(new_n767));
  XOR2_X1   g581(.A(new_n748), .B(KEYINPUT107), .Z(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(G469), .B1(new_n319), .B2(KEYINPUT45), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT106), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT106), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n772), .B(G469), .C1(new_n319), .C2(KEYINPUT45), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n319), .A2(KEYINPUT45), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n771), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(G469), .A2(G902), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT46), .ZN(new_n778));
  AOI22_X1  g592(.A1(new_n777), .A2(new_n778), .B1(new_n307), .B2(new_n312), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n775), .A2(KEYINPUT46), .A3(new_n776), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n316), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n698), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n769), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(new_n192), .ZN(G39));
  NAND2_X1  g598(.A1(new_n777), .A2(new_n778), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n785), .A2(new_n720), .A3(new_n780), .ZN(new_n786));
  XOR2_X1   g600(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n786), .A2(new_n315), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n789), .B1(new_n781), .B2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n748), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n717), .A2(new_n792), .A3(new_n384), .ZN(new_n793));
  OR3_X1    g607(.A1(new_n791), .A2(new_n685), .A3(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G140), .ZN(G42));
  INV_X1    g609(.A(KEYINPUT112), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n688), .A2(new_n627), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n709), .A2(KEYINPUT90), .A3(new_n565), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n550), .A2(new_n552), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n513), .A2(new_n799), .A3(new_n563), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT111), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT111), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n797), .A2(new_n798), .A3(new_n803), .A4(new_n800), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n802), .A2(new_n638), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n796), .B1(new_n805), .B2(new_n681), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n805), .A2(new_n681), .A3(new_n796), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n669), .A2(new_n759), .A3(new_n563), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n797), .A2(new_n798), .A3(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT109), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n797), .A2(new_n798), .A3(KEYINPUT109), .A4(new_n810), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n638), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n630), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT110), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT110), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n815), .A2(new_n630), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  AND4_X1   g634(.A1(new_n723), .A2(new_n726), .A3(new_n730), .A4(new_n737), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n821), .A2(new_n754), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n749), .A2(new_n717), .A3(new_n744), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n756), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n669), .A2(new_n799), .A3(new_n693), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n825), .A2(new_n748), .A3(new_n678), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n326), .A2(new_n685), .A3(new_n826), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n827), .A2(KEYINPUT113), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(KEYINPUT113), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n824), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AND4_X1   g644(.A1(new_n809), .A2(new_n820), .A3(new_n822), .A4(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n746), .A2(new_n696), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n313), .A2(new_n316), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n693), .B(KEYINPUT114), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n736), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n708), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n718), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n833), .B1(new_n834), .B2(new_n839), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n690), .A2(new_n717), .B1(new_n837), .B2(new_n708), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(KEYINPUT52), .A3(new_n696), .A4(new_n746), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n831), .A2(new_n832), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n807), .A2(new_n808), .B1(new_n817), .B2(new_n819), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n847), .A2(new_n843), .A3(new_n830), .A4(new_n822), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT116), .B1(new_n848), .B2(new_n844), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT53), .B1(new_n831), .B2(new_n843), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n846), .B(KEYINPUT54), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n805), .A2(new_n796), .A3(new_n681), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n815), .A2(new_n818), .A3(new_n630), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n818), .B1(new_n815), .B2(new_n630), .ZN(new_n855));
  OAI22_X1  g669(.A1(new_n806), .A2(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n827), .B(KEYINPUT113), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(new_n756), .A3(new_n823), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n852), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n809), .A2(new_n820), .A3(new_n830), .A4(KEYINPUT117), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n821), .A2(new_n754), .A3(KEYINPUT53), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n840), .B2(new_n842), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n809), .A2(new_n820), .A3(new_n830), .A4(new_n822), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n840), .A2(new_n842), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n844), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n863), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT118), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT118), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n863), .A2(new_n867), .A3(new_n870), .A4(new_n864), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n872));
  XNOR2_X1  g686(.A(KEYINPUT119), .B(KEYINPUT50), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n763), .A2(new_n559), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n875), .A2(new_n722), .A3(new_n735), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n711), .A2(new_n566), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n874), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n875), .A2(new_n722), .A3(new_n735), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT50), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT119), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n880), .A2(new_n882), .A3(new_n877), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n728), .A2(new_n559), .A3(new_n748), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n513), .A2(new_n656), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n884), .A2(new_n707), .A3(new_n383), .A4(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n884), .A2(new_n744), .A3(new_n764), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n879), .A2(new_n883), .A3(new_n888), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n720), .A2(new_n721), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(new_n315), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n786), .A2(new_n315), .ZN(new_n893));
  INV_X1    g707(.A(new_n790), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n892), .B1(new_n895), .B2(new_n789), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n768), .A2(new_n735), .A3(new_n875), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n889), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT51), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n884), .A2(new_n764), .ZN(new_n900));
  INV_X1    g714(.A(new_n456), .ZN(new_n901));
  OAI21_X1  g715(.A(KEYINPUT48), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT48), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n884), .A2(new_n456), .A3(new_n903), .A4(new_n764), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n875), .A2(new_n625), .A3(new_n722), .A4(new_n735), .ZN(new_n906));
  INV_X1    g720(.A(new_n657), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n884), .A2(new_n707), .A3(new_n383), .A4(new_n907), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n906), .A2(new_n557), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT120), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n905), .A2(new_n909), .A3(KEYINPUT120), .ZN(new_n913));
  AOI22_X1  g727(.A1(new_n898), .A2(new_n899), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n889), .B(KEYINPUT51), .C1(new_n896), .C2(new_n897), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n872), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n892), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n897), .B1(new_n791), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n883), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n873), .B1(new_n880), .B2(new_n877), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n919), .A2(new_n920), .A3(new_n887), .A4(new_n886), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n899), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n912), .A2(new_n913), .ZN(new_n923));
  AND4_X1   g737(.A1(new_n872), .A2(new_n922), .A3(new_n915), .A4(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n916), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n851), .A2(new_n869), .A3(new_n871), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n556), .A2(new_n280), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n890), .B(KEYINPUT49), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n383), .A2(new_n315), .A3(new_n565), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n930), .A2(new_n513), .A3(new_n759), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n929), .A2(new_n707), .A3(new_n711), .A4(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(KEYINPUT122), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT122), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n928), .A2(new_n935), .A3(new_n932), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n934), .A2(new_n936), .ZN(G75));
  NOR2_X1   g751(.A1(new_n284), .A2(G952), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n300), .B1(new_n863), .B2(new_n867), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(G210), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n586), .B(new_n596), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT55), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n944), .A2(KEYINPUT56), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n939), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT56), .B1(new_n941), .B2(KEYINPUT123), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n947), .B1(KEYINPUT123), .B2(new_n941), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n946), .B1(new_n948), .B2(new_n944), .ZN(G51));
  NAND2_X1  g763(.A1(new_n863), .A2(new_n867), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(KEYINPUT54), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n868), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n776), .B(KEYINPUT57), .Z(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n321), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n940), .A2(new_n773), .A3(new_n774), .A4(new_n771), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n938), .B1(new_n955), .B2(new_n956), .ZN(G54));
  NAND3_X1  g771(.A1(new_n940), .A2(KEYINPUT58), .A3(G475), .ZN(new_n958));
  INV_X1    g772(.A(new_n506), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n958), .A2(new_n959), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n960), .A2(new_n961), .A3(new_n938), .ZN(G60));
  NAND3_X1  g776(.A1(new_n851), .A2(new_n869), .A3(new_n871), .ZN(new_n963));
  NAND2_X1  g777(.A1(G478), .A2(G902), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT59), .Z(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n758), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n952), .A2(new_n758), .A3(new_n966), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n967), .A2(new_n968), .A3(new_n938), .ZN(G63));
  INV_X1    g783(.A(KEYINPUT61), .ZN(new_n970));
  NAND2_X1  g784(.A1(G217), .A2(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT60), .Z(new_n972));
  NAND2_X1  g786(.A1(new_n950), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(KEYINPUT124), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT124), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n950), .A2(new_n975), .A3(new_n972), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n974), .A2(new_n370), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n939), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n676), .B1(new_n974), .B2(new_n976), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n970), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n979), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n981), .A2(KEYINPUT61), .A3(new_n939), .A4(new_n977), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(G66));
  INV_X1    g797(.A(new_n562), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n280), .B1(new_n984), .B2(G224), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n847), .A2(new_n821), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n985), .B1(new_n986), .B2(new_n284), .ZN(new_n987));
  INV_X1    g801(.A(G898), .ZN(new_n988));
  INV_X1    g802(.A(new_n284), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n586), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n987), .B(new_n990), .ZN(G69));
  AND3_X1   g805(.A1(new_n746), .A2(new_n696), .A3(new_n718), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n714), .A2(new_n992), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n657), .B1(new_n513), .B2(new_n799), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n456), .A2(new_n792), .A3(new_n995), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n699), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n783), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n994), .A2(new_n998), .A3(new_n794), .A4(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n284), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n409), .A2(new_n412), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(new_n502), .Z(new_n1003));
  XNOR2_X1  g817(.A(new_n1003), .B(KEYINPUT125), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT126), .ZN(new_n1006));
  INV_X1    g820(.A(G227), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n989), .B1(new_n1007), .B2(new_n691), .ZN(new_n1008));
  INV_X1    g822(.A(new_n783), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n781), .A2(new_n456), .A3(new_n698), .A4(new_n736), .ZN(new_n1010));
  AND3_X1   g824(.A1(new_n1009), .A2(new_n756), .A3(new_n1010), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n1011), .A2(new_n754), .A3(new_n794), .A4(new_n992), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n1012), .A2(new_n989), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1003), .B1(new_n691), .B2(new_n284), .ZN(new_n1014));
  OAI221_X1 g828(.A(new_n1005), .B1(new_n1006), .B2(new_n1008), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1008), .A2(new_n1006), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1015), .B(new_n1016), .ZN(G72));
  NAND2_X1  g831(.A1(G472), .A2(G902), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1018), .B(KEYINPUT63), .Z(new_n1019));
  OAI21_X1  g833(.A(new_n1019), .B1(new_n1000), .B2(new_n986), .ZN(new_n1020));
  INV_X1    g834(.A(new_n702), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1022), .B(KEYINPUT127), .Z(new_n1023));
  NOR2_X1   g837(.A1(new_n415), .A2(new_n445), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1019), .ZN(new_n1025));
  NOR3_X1   g839(.A1(new_n1021), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  OAI211_X1 g840(.A(new_n846), .B(new_n1026), .C1(new_n849), .C2(new_n850), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1019), .B1(new_n1012), .B2(new_n986), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n938), .B1(new_n1028), .B2(new_n1024), .ZN(new_n1029));
  AND3_X1   g843(.A1(new_n1023), .A2(new_n1027), .A3(new_n1029), .ZN(G57));
endmodule


