

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U552 ( .A1(n684), .A2(n757), .ZN(n686) );
  OR2_X1 U553 ( .A1(n796), .A2(n755), .ZN(n519) );
  AND2_X1 U554 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U555 ( .A(n689), .B(KEYINPUT90), .ZN(n706) );
  INV_X1 U556 ( .A(n686), .ZN(n714) );
  BUF_X1 U557 ( .A(n686), .Z(n729) );
  INV_X1 U558 ( .A(KEYINPUT84), .ZN(n524) );
  NOR2_X1 U559 ( .A1(n530), .A2(n520), .ZN(n889) );
  NOR2_X1 U560 ( .A1(G651), .A2(n634), .ZN(n648) );
  NOR2_X1 U561 ( .A1(n533), .A2(n532), .ZN(G164) );
  INV_X1 U562 ( .A(G2104), .ZN(n530) );
  INV_X1 U563 ( .A(G2105), .ZN(n520) );
  NAND2_X1 U564 ( .A1(G114), .A2(n889), .ZN(n523) );
  NOR2_X1 U565 ( .A1(n520), .A2(G2104), .ZN(n521) );
  XNOR2_X1 U566 ( .A(n521), .B(KEYINPUT64), .ZN(n537) );
  NAND2_X1 U567 ( .A1(G126), .A2(n537), .ZN(n522) );
  NAND2_X1 U568 ( .A1(n523), .A2(n522), .ZN(n525) );
  XNOR2_X1 U569 ( .A(n525), .B(n524), .ZN(n529) );
  XNOR2_X1 U570 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n527) );
  NOR2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  XNOR2_X2 U572 ( .A(n527), .B(n526), .ZN(n885) );
  NAND2_X1 U573 ( .A1(n885), .A2(G138), .ZN(n528) );
  NAND2_X1 U574 ( .A1(n529), .A2(n528), .ZN(n533) );
  NOR2_X1 U575 ( .A1(G2105), .A2(n530), .ZN(n886) );
  NAND2_X1 U576 ( .A1(G102), .A2(n886), .ZN(n531) );
  XNOR2_X1 U577 ( .A(KEYINPUT85), .B(n531), .ZN(n532) );
  NAND2_X1 U578 ( .A1(n885), .A2(G137), .ZN(n535) );
  NAND2_X1 U579 ( .A1(n889), .A2(G113), .ZN(n534) );
  NAND2_X1 U580 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U581 ( .A(n536), .B(KEYINPUT66), .ZN(n539) );
  AND2_X1 U582 ( .A1(G125), .A2(n537), .ZN(n538) );
  NOR2_X1 U583 ( .A1(n539), .A2(n538), .ZN(n682) );
  NAND2_X1 U584 ( .A1(G101), .A2(n886), .ZN(n540) );
  XOR2_X1 U585 ( .A(KEYINPUT23), .B(n540), .Z(n680) );
  AND2_X1 U586 ( .A1(n682), .A2(n680), .ZN(G160) );
  AND2_X1 U587 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U588 ( .A(G57), .ZN(G237) );
  XOR2_X1 U589 ( .A(G543), .B(KEYINPUT0), .Z(n634) );
  NAND2_X1 U590 ( .A1(n648), .A2(G51), .ZN(n541) );
  XOR2_X1 U591 ( .A(KEYINPUT75), .B(n541), .Z(n545) );
  INV_X1 U592 ( .A(G651), .ZN(n548) );
  NOR2_X1 U593 ( .A1(G543), .A2(n548), .ZN(n543) );
  XNOR2_X1 U594 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n542) );
  XNOR2_X1 U595 ( .A(n543), .B(n542), .ZN(n647) );
  NAND2_X1 U596 ( .A1(n647), .A2(G63), .ZN(n544) );
  NAND2_X1 U597 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U598 ( .A(KEYINPUT6), .B(n546), .ZN(n556) );
  NOR2_X1 U599 ( .A1(G651), .A2(G543), .ZN(n643) );
  NAND2_X1 U600 ( .A1(n643), .A2(G89), .ZN(n547) );
  XOR2_X1 U601 ( .A(KEYINPUT4), .B(n547), .Z(n551) );
  NOR2_X1 U602 ( .A1(n634), .A2(n548), .ZN(n644) );
  NAND2_X1 U603 ( .A1(n644), .A2(G76), .ZN(n549) );
  XOR2_X1 U604 ( .A(n549), .B(KEYINPUT72), .Z(n550) );
  NOR2_X1 U605 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U606 ( .A(KEYINPUT5), .B(n552), .Z(n554) );
  XNOR2_X1 U607 ( .A(KEYINPUT73), .B(KEYINPUT74), .ZN(n553) );
  XNOR2_X1 U608 ( .A(n554), .B(n553), .ZN(n555) );
  NOR2_X1 U609 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U610 ( .A(KEYINPUT7), .B(n557), .Z(G168) );
  XOR2_X1 U611 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U612 ( .A1(G7), .A2(G661), .ZN(n558) );
  XNOR2_X1 U613 ( .A(n558), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U614 ( .A(G223), .B(KEYINPUT69), .ZN(n822) );
  NAND2_X1 U615 ( .A1(n822), .A2(G567), .ZN(n559) );
  XOR2_X1 U616 ( .A(KEYINPUT11), .B(n559), .Z(G234) );
  NAND2_X1 U617 ( .A1(G56), .A2(n647), .ZN(n560) );
  XOR2_X1 U618 ( .A(KEYINPUT14), .B(n560), .Z(n566) );
  NAND2_X1 U619 ( .A1(n643), .A2(G81), .ZN(n561) );
  XNOR2_X1 U620 ( .A(n561), .B(KEYINPUT12), .ZN(n563) );
  NAND2_X1 U621 ( .A1(G68), .A2(n644), .ZN(n562) );
  NAND2_X1 U622 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U623 ( .A(KEYINPUT13), .B(n564), .Z(n565) );
  NOR2_X1 U624 ( .A1(n566), .A2(n565), .ZN(n568) );
  NAND2_X1 U625 ( .A1(n648), .A2(G43), .ZN(n567) );
  NAND2_X1 U626 ( .A1(n568), .A2(n567), .ZN(n947) );
  INV_X1 U627 ( .A(G860), .ZN(n613) );
  OR2_X1 U628 ( .A1(n947), .A2(n613), .ZN(G153) );
  NAND2_X1 U629 ( .A1(G90), .A2(n643), .ZN(n570) );
  NAND2_X1 U630 ( .A1(G77), .A2(n644), .ZN(n569) );
  NAND2_X1 U631 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U632 ( .A(KEYINPUT9), .B(n571), .ZN(n575) );
  NAND2_X1 U633 ( .A1(G64), .A2(n647), .ZN(n573) );
  NAND2_X1 U634 ( .A1(G52), .A2(n648), .ZN(n572) );
  AND2_X1 U635 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U636 ( .A1(n575), .A2(n574), .ZN(G301) );
  NAND2_X1 U637 ( .A1(G66), .A2(n647), .ZN(n577) );
  NAND2_X1 U638 ( .A1(G92), .A2(n643), .ZN(n576) );
  NAND2_X1 U639 ( .A1(n577), .A2(n576), .ZN(n582) );
  NAND2_X1 U640 ( .A1(G79), .A2(n644), .ZN(n579) );
  NAND2_X1 U641 ( .A1(G54), .A2(n648), .ZN(n578) );
  NAND2_X1 U642 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT70), .B(n580), .ZN(n581) );
  NOR2_X1 U644 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U645 ( .A(n583), .B(KEYINPUT15), .ZN(n937) );
  INV_X1 U646 ( .A(n937), .ZN(n611) );
  NOR2_X1 U647 ( .A1(n611), .A2(G868), .ZN(n584) );
  XNOR2_X1 U648 ( .A(n584), .B(KEYINPUT71), .ZN(n586) );
  NAND2_X1 U649 ( .A1(G868), .A2(G301), .ZN(n585) );
  NAND2_X1 U650 ( .A1(n586), .A2(n585), .ZN(G284) );
  NAND2_X1 U651 ( .A1(G65), .A2(n647), .ZN(n588) );
  NAND2_X1 U652 ( .A1(G91), .A2(n643), .ZN(n587) );
  NAND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U654 ( .A1(n644), .A2(G78), .ZN(n589) );
  XOR2_X1 U655 ( .A(KEYINPUT68), .B(n589), .Z(n590) );
  NOR2_X1 U656 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U657 ( .A1(n648), .A2(G53), .ZN(n592) );
  NAND2_X1 U658 ( .A1(n593), .A2(n592), .ZN(G299) );
  INV_X1 U659 ( .A(G868), .ZN(n661) );
  NOR2_X1 U660 ( .A1(G286), .A2(n661), .ZN(n595) );
  NOR2_X1 U661 ( .A1(G868), .A2(G299), .ZN(n594) );
  NOR2_X1 U662 ( .A1(n595), .A2(n594), .ZN(G297) );
  NAND2_X1 U663 ( .A1(n613), .A2(G559), .ZN(n596) );
  NAND2_X1 U664 ( .A1(n596), .A2(n611), .ZN(n597) );
  XNOR2_X1 U665 ( .A(n597), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U666 ( .A1(G868), .A2(n947), .ZN(n600) );
  NAND2_X1 U667 ( .A1(G868), .A2(n611), .ZN(n598) );
  NOR2_X1 U668 ( .A1(G559), .A2(n598), .ZN(n599) );
  NOR2_X1 U669 ( .A1(n600), .A2(n599), .ZN(G282) );
  NAND2_X1 U670 ( .A1(n885), .A2(G135), .ZN(n607) );
  NAND2_X1 U671 ( .A1(G111), .A2(n889), .ZN(n602) );
  NAND2_X1 U672 ( .A1(G99), .A2(n886), .ZN(n601) );
  NAND2_X1 U673 ( .A1(n602), .A2(n601), .ZN(n605) );
  NAND2_X1 U674 ( .A1(n537), .A2(G123), .ZN(n603) );
  XOR2_X1 U675 ( .A(KEYINPUT18), .B(n603), .Z(n604) );
  NOR2_X1 U676 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U677 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U678 ( .A(KEYINPUT76), .B(n608), .Z(n998) );
  XNOR2_X1 U679 ( .A(n998), .B(G2096), .ZN(n610) );
  INV_X1 U680 ( .A(G2100), .ZN(n609) );
  NAND2_X1 U681 ( .A1(n610), .A2(n609), .ZN(G156) );
  NAND2_X1 U682 ( .A1(G559), .A2(n611), .ZN(n612) );
  XOR2_X1 U683 ( .A(n947), .B(n612), .Z(n659) );
  NAND2_X1 U684 ( .A1(n613), .A2(n659), .ZN(n621) );
  NAND2_X1 U685 ( .A1(G67), .A2(n647), .ZN(n615) );
  NAND2_X1 U686 ( .A1(G93), .A2(n643), .ZN(n614) );
  NAND2_X1 U687 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U688 ( .A1(G80), .A2(n644), .ZN(n616) );
  XNOR2_X1 U689 ( .A(KEYINPUT77), .B(n616), .ZN(n617) );
  NOR2_X1 U690 ( .A1(n618), .A2(n617), .ZN(n620) );
  NAND2_X1 U691 ( .A1(n648), .A2(G55), .ZN(n619) );
  NAND2_X1 U692 ( .A1(n620), .A2(n619), .ZN(n662) );
  XNOR2_X1 U693 ( .A(n621), .B(n662), .ZN(G145) );
  XOR2_X1 U694 ( .A(KEYINPUT79), .B(KEYINPUT2), .Z(n623) );
  NAND2_X1 U695 ( .A1(G73), .A2(n644), .ZN(n622) );
  XNOR2_X1 U696 ( .A(n623), .B(n622), .ZN(n630) );
  NAND2_X1 U697 ( .A1(G61), .A2(n647), .ZN(n625) );
  NAND2_X1 U698 ( .A1(G48), .A2(n648), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U700 ( .A1(n643), .A2(G86), .ZN(n626) );
  XOR2_X1 U701 ( .A(KEYINPUT78), .B(n626), .Z(n627) );
  NOR2_X1 U702 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U703 ( .A1(n630), .A2(n629), .ZN(G305) );
  NAND2_X1 U704 ( .A1(G49), .A2(n648), .ZN(n632) );
  NAND2_X1 U705 ( .A1(G74), .A2(G651), .ZN(n631) );
  NAND2_X1 U706 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U707 ( .A1(n647), .A2(n633), .ZN(n636) );
  NAND2_X1 U708 ( .A1(n634), .A2(G87), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n636), .A2(n635), .ZN(G288) );
  AND2_X1 U710 ( .A1(n647), .A2(G60), .ZN(n640) );
  NAND2_X1 U711 ( .A1(G85), .A2(n643), .ZN(n638) );
  NAND2_X1 U712 ( .A1(G72), .A2(n644), .ZN(n637) );
  NAND2_X1 U713 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U714 ( .A1(n640), .A2(n639), .ZN(n642) );
  NAND2_X1 U715 ( .A1(n648), .A2(G47), .ZN(n641) );
  NAND2_X1 U716 ( .A1(n642), .A2(n641), .ZN(G290) );
  NAND2_X1 U717 ( .A1(G88), .A2(n643), .ZN(n646) );
  NAND2_X1 U718 ( .A1(G75), .A2(n644), .ZN(n645) );
  NAND2_X1 U719 ( .A1(n646), .A2(n645), .ZN(n652) );
  NAND2_X1 U720 ( .A1(G62), .A2(n647), .ZN(n650) );
  NAND2_X1 U721 ( .A1(G50), .A2(n648), .ZN(n649) );
  NAND2_X1 U722 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U723 ( .A1(n652), .A2(n651), .ZN(G166) );
  INV_X1 U724 ( .A(G166), .ZN(G303) );
  INV_X1 U725 ( .A(G299), .ZN(n940) );
  XNOR2_X1 U726 ( .A(n940), .B(G305), .ZN(n653) );
  XNOR2_X1 U727 ( .A(n653), .B(n662), .ZN(n654) );
  XNOR2_X1 U728 ( .A(KEYINPUT19), .B(n654), .ZN(n656) );
  XNOR2_X1 U729 ( .A(G288), .B(KEYINPUT80), .ZN(n655) );
  XNOR2_X1 U730 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U731 ( .A(n657), .B(G290), .ZN(n658) );
  XNOR2_X1 U732 ( .A(n658), .B(G303), .ZN(n903) );
  XOR2_X1 U733 ( .A(n903), .B(n659), .Z(n660) );
  NOR2_X1 U734 ( .A1(n661), .A2(n660), .ZN(n664) );
  NOR2_X1 U735 ( .A1(G868), .A2(n662), .ZN(n663) );
  NOR2_X1 U736 ( .A1(n664), .A2(n663), .ZN(G295) );
  NAND2_X1 U737 ( .A1(G2084), .A2(G2078), .ZN(n665) );
  XNOR2_X1 U738 ( .A(n665), .B(KEYINPUT81), .ZN(n666) );
  XNOR2_X1 U739 ( .A(n666), .B(KEYINPUT20), .ZN(n667) );
  NAND2_X1 U740 ( .A1(n667), .A2(G2090), .ZN(n668) );
  XNOR2_X1 U741 ( .A(n668), .B(KEYINPUT82), .ZN(n669) );
  XNOR2_X1 U742 ( .A(n669), .B(KEYINPUT21), .ZN(n670) );
  NAND2_X1 U743 ( .A1(n670), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U744 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U745 ( .A(KEYINPUT83), .B(KEYINPUT22), .Z(n672) );
  NAND2_X1 U746 ( .A1(G132), .A2(G82), .ZN(n671) );
  XNOR2_X1 U747 ( .A(n672), .B(n671), .ZN(n673) );
  NOR2_X1 U748 ( .A1(n673), .A2(G218), .ZN(n674) );
  NAND2_X1 U749 ( .A1(G96), .A2(n674), .ZN(n828) );
  NAND2_X1 U750 ( .A1(n828), .A2(G2106), .ZN(n678) );
  NAND2_X1 U751 ( .A1(G69), .A2(G120), .ZN(n675) );
  NOR2_X1 U752 ( .A1(G237), .A2(n675), .ZN(n676) );
  NAND2_X1 U753 ( .A1(G108), .A2(n676), .ZN(n827) );
  NAND2_X1 U754 ( .A1(n827), .A2(G567), .ZN(n677) );
  NAND2_X1 U755 ( .A1(n678), .A2(n677), .ZN(n914) );
  NAND2_X1 U756 ( .A1(G483), .A2(G661), .ZN(n679) );
  NOR2_X1 U757 ( .A1(n914), .A2(n679), .ZN(n826) );
  NAND2_X1 U758 ( .A1(n826), .A2(G36), .ZN(G176) );
  INV_X1 U759 ( .A(G301), .ZN(G171) );
  AND2_X1 U760 ( .A1(n680), .A2(G40), .ZN(n681) );
  NAND2_X1 U761 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U762 ( .A(n683), .B(KEYINPUT86), .ZN(n758) );
  INV_X1 U763 ( .A(n758), .ZN(n684) );
  NOR2_X1 U764 ( .A1(G164), .A2(G1384), .ZN(n757) );
  NAND2_X1 U765 ( .A1(G8), .A2(n686), .ZN(n796) );
  NAND2_X1 U766 ( .A1(n714), .A2(G2072), .ZN(n685) );
  XOR2_X1 U767 ( .A(KEYINPUT27), .B(n685), .Z(n688) );
  NAND2_X1 U768 ( .A1(G1956), .A2(n729), .ZN(n687) );
  NOR2_X1 U769 ( .A1(n940), .A2(n706), .ZN(n691) );
  XNOR2_X1 U770 ( .A(KEYINPUT91), .B(KEYINPUT28), .ZN(n690) );
  XNOR2_X1 U771 ( .A(n691), .B(n690), .ZN(n710) );
  XOR2_X1 U772 ( .A(KEYINPUT26), .B(KEYINPUT92), .Z(n693) );
  NAND2_X1 U773 ( .A1(n714), .A2(G1996), .ZN(n692) );
  XNOR2_X1 U774 ( .A(n693), .B(n692), .ZN(n694) );
  NOR2_X1 U775 ( .A1(n694), .A2(n947), .ZN(n696) );
  NAND2_X1 U776 ( .A1(G1341), .A2(n729), .ZN(n695) );
  NAND2_X1 U777 ( .A1(n696), .A2(n695), .ZN(n703) );
  NOR2_X1 U778 ( .A1(n937), .A2(n703), .ZN(n697) );
  XNOR2_X1 U779 ( .A(n697), .B(KEYINPUT93), .ZN(n702) );
  AND2_X1 U780 ( .A1(n714), .A2(G2067), .ZN(n698) );
  XOR2_X1 U781 ( .A(n698), .B(KEYINPUT94), .Z(n700) );
  NAND2_X1 U782 ( .A1(n729), .A2(G1348), .ZN(n699) );
  NAND2_X1 U783 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U784 ( .A1(n702), .A2(n701), .ZN(n705) );
  NAND2_X1 U785 ( .A1(n937), .A2(n703), .ZN(n704) );
  NAND2_X1 U786 ( .A1(n705), .A2(n704), .ZN(n708) );
  NAND2_X1 U787 ( .A1(n940), .A2(n706), .ZN(n707) );
  NAND2_X1 U788 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U789 ( .A1(n710), .A2(n709), .ZN(n712) );
  XNOR2_X1 U790 ( .A(KEYINPUT95), .B(KEYINPUT29), .ZN(n711) );
  XNOR2_X1 U791 ( .A(n712), .B(n711), .ZN(n718) );
  NOR2_X1 U792 ( .A1(n714), .A2(G1961), .ZN(n713) );
  XNOR2_X1 U793 ( .A(n713), .B(KEYINPUT89), .ZN(n716) );
  XNOR2_X1 U794 ( .A(KEYINPUT25), .B(G2078), .ZN(n925) );
  NAND2_X1 U795 ( .A1(n714), .A2(n925), .ZN(n715) );
  NAND2_X1 U796 ( .A1(n716), .A2(n715), .ZN(n722) );
  NAND2_X1 U797 ( .A1(n722), .A2(G171), .ZN(n717) );
  NAND2_X1 U798 ( .A1(n718), .A2(n717), .ZN(n728) );
  NOR2_X1 U799 ( .A1(G1966), .A2(n796), .ZN(n741) );
  NOR2_X1 U800 ( .A1(G2084), .A2(n729), .ZN(n740) );
  NOR2_X1 U801 ( .A1(n741), .A2(n740), .ZN(n719) );
  NAND2_X1 U802 ( .A1(G8), .A2(n719), .ZN(n720) );
  XNOR2_X1 U803 ( .A(KEYINPUT30), .B(n720), .ZN(n721) );
  NOR2_X1 U804 ( .A1(G168), .A2(n721), .ZN(n724) );
  NOR2_X1 U805 ( .A1(G171), .A2(n722), .ZN(n723) );
  NOR2_X1 U806 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U807 ( .A(n725), .B(KEYINPUT31), .Z(n726) );
  XNOR2_X1 U808 ( .A(KEYINPUT96), .B(n726), .ZN(n727) );
  NAND2_X1 U809 ( .A1(n728), .A2(n727), .ZN(n744) );
  NAND2_X1 U810 ( .A1(n744), .A2(G286), .ZN(n737) );
  INV_X1 U811 ( .A(G8), .ZN(n735) );
  NOR2_X1 U812 ( .A1(G2090), .A2(n729), .ZN(n730) );
  XNOR2_X1 U813 ( .A(KEYINPUT97), .B(n730), .ZN(n733) );
  NOR2_X1 U814 ( .A1(G1971), .A2(n796), .ZN(n731) );
  NOR2_X1 U815 ( .A1(G166), .A2(n731), .ZN(n732) );
  NAND2_X1 U816 ( .A1(n733), .A2(n732), .ZN(n734) );
  OR2_X1 U817 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U818 ( .A1(n737), .A2(n736), .ZN(n739) );
  INV_X1 U819 ( .A(KEYINPUT32), .ZN(n738) );
  XNOR2_X1 U820 ( .A(n739), .B(n738), .ZN(n788) );
  AND2_X1 U821 ( .A1(G8), .A2(n740), .ZN(n742) );
  NOR2_X1 U822 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U823 ( .A1(n744), .A2(n743), .ZN(n789) );
  NAND2_X1 U824 ( .A1(G1976), .A2(G288), .ZN(n945) );
  AND2_X1 U825 ( .A1(n789), .A2(n945), .ZN(n745) );
  NAND2_X1 U826 ( .A1(n788), .A2(n745), .ZN(n751) );
  INV_X1 U827 ( .A(n945), .ZN(n749) );
  NOR2_X1 U828 ( .A1(G1976), .A2(G288), .ZN(n944) );
  NOR2_X1 U829 ( .A1(G1971), .A2(G303), .ZN(n746) );
  XNOR2_X1 U830 ( .A(KEYINPUT98), .B(n746), .ZN(n747) );
  NOR2_X1 U831 ( .A1(n944), .A2(n747), .ZN(n748) );
  OR2_X1 U832 ( .A1(n749), .A2(n748), .ZN(n750) );
  AND2_X1 U833 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U834 ( .A1(n796), .A2(n752), .ZN(n753) );
  NOR2_X1 U835 ( .A1(KEYINPUT33), .A2(n753), .ZN(n754) );
  XNOR2_X1 U836 ( .A(KEYINPUT99), .B(n754), .ZN(n756) );
  NAND2_X1 U837 ( .A1(n944), .A2(KEYINPUT33), .ZN(n755) );
  AND2_X1 U838 ( .A1(n756), .A2(n519), .ZN(n787) );
  XOR2_X1 U839 ( .A(G1981), .B(G305), .Z(n955) );
  NOR2_X1 U840 ( .A1(n758), .A2(n757), .ZN(n816) );
  XNOR2_X1 U841 ( .A(G2067), .B(KEYINPUT37), .ZN(n801) );
  NAND2_X1 U842 ( .A1(G140), .A2(n885), .ZN(n760) );
  NAND2_X1 U843 ( .A1(G104), .A2(n886), .ZN(n759) );
  NAND2_X1 U844 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U845 ( .A(KEYINPUT34), .B(n761), .ZN(n766) );
  NAND2_X1 U846 ( .A1(G116), .A2(n889), .ZN(n763) );
  NAND2_X1 U847 ( .A1(G128), .A2(n537), .ZN(n762) );
  NAND2_X1 U848 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U849 ( .A(KEYINPUT35), .B(n764), .Z(n765) );
  NOR2_X1 U850 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U851 ( .A(KEYINPUT36), .B(n767), .ZN(n899) );
  NOR2_X1 U852 ( .A1(n801), .A2(n899), .ZN(n1003) );
  NAND2_X1 U853 ( .A1(n816), .A2(n1003), .ZN(n809) );
  NAND2_X1 U854 ( .A1(G131), .A2(n885), .ZN(n769) );
  NAND2_X1 U855 ( .A1(G107), .A2(n889), .ZN(n768) );
  NAND2_X1 U856 ( .A1(n769), .A2(n768), .ZN(n772) );
  NAND2_X1 U857 ( .A1(G95), .A2(n886), .ZN(n770) );
  XNOR2_X1 U858 ( .A(KEYINPUT87), .B(n770), .ZN(n771) );
  NOR2_X1 U859 ( .A1(n772), .A2(n771), .ZN(n774) );
  NAND2_X1 U860 ( .A1(G119), .A2(n537), .ZN(n773) );
  NAND2_X1 U861 ( .A1(n774), .A2(n773), .ZN(n881) );
  AND2_X1 U862 ( .A1(n881), .A2(G1991), .ZN(n784) );
  NAND2_X1 U863 ( .A1(G141), .A2(n885), .ZN(n776) );
  NAND2_X1 U864 ( .A1(G117), .A2(n889), .ZN(n775) );
  NAND2_X1 U865 ( .A1(n776), .A2(n775), .ZN(n779) );
  NAND2_X1 U866 ( .A1(n886), .A2(G105), .ZN(n777) );
  XOR2_X1 U867 ( .A(KEYINPUT38), .B(n777), .Z(n778) );
  NOR2_X1 U868 ( .A1(n779), .A2(n778), .ZN(n781) );
  NAND2_X1 U869 ( .A1(G129), .A2(n537), .ZN(n780) );
  NAND2_X1 U870 ( .A1(n781), .A2(n780), .ZN(n880) );
  NAND2_X1 U871 ( .A1(G1996), .A2(n880), .ZN(n782) );
  XOR2_X1 U872 ( .A(KEYINPUT88), .B(n782), .Z(n783) );
  NOR2_X1 U873 ( .A1(n784), .A2(n783), .ZN(n1000) );
  INV_X1 U874 ( .A(n1000), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n785), .A2(n816), .ZN(n802) );
  AND2_X1 U876 ( .A1(n809), .A2(n802), .ZN(n800) );
  AND2_X1 U877 ( .A1(n955), .A2(n800), .ZN(n786) );
  NAND2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n815) );
  NAND2_X1 U879 ( .A1(n789), .A2(n788), .ZN(n792) );
  NOR2_X1 U880 ( .A1(G2090), .A2(G303), .ZN(n790) );
  NAND2_X1 U881 ( .A1(G8), .A2(n790), .ZN(n791) );
  NAND2_X1 U882 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U883 ( .A1(n793), .A2(n796), .ZN(n798) );
  NOR2_X1 U884 ( .A1(G1981), .A2(G305), .ZN(n794) );
  XOR2_X1 U885 ( .A(n794), .B(KEYINPUT24), .Z(n795) );
  OR2_X1 U886 ( .A1(n796), .A2(n795), .ZN(n797) );
  NAND2_X1 U887 ( .A1(n798), .A2(n797), .ZN(n799) );
  AND2_X1 U888 ( .A1(n800), .A2(n799), .ZN(n813) );
  NAND2_X1 U889 ( .A1(n801), .A2(n899), .ZN(n1010) );
  NOR2_X1 U890 ( .A1(G1996), .A2(n880), .ZN(n994) );
  INV_X1 U891 ( .A(n802), .ZN(n805) );
  NOR2_X1 U892 ( .A1(G1986), .A2(G290), .ZN(n803) );
  NOR2_X1 U893 ( .A1(G1991), .A2(n881), .ZN(n999) );
  NOR2_X1 U894 ( .A1(n803), .A2(n999), .ZN(n804) );
  NOR2_X1 U895 ( .A1(n805), .A2(n804), .ZN(n806) );
  NOR2_X1 U896 ( .A1(n994), .A2(n806), .ZN(n807) );
  XNOR2_X1 U897 ( .A(KEYINPUT39), .B(n807), .ZN(n808) );
  XNOR2_X1 U898 ( .A(n808), .B(KEYINPUT100), .ZN(n810) );
  NAND2_X1 U899 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U900 ( .A1(n1010), .A2(n811), .ZN(n812) );
  AND2_X1 U901 ( .A1(n812), .A2(n816), .ZN(n818) );
  NOR2_X1 U902 ( .A1(n813), .A2(n818), .ZN(n814) );
  NAND2_X1 U903 ( .A1(n815), .A2(n814), .ZN(n820) );
  XNOR2_X1 U904 ( .A(G1986), .B(G290), .ZN(n939) );
  NAND2_X1 U905 ( .A1(n939), .A2(n816), .ZN(n817) );
  OR2_X1 U906 ( .A1(n818), .A2(n817), .ZN(n819) );
  AND2_X1 U907 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U908 ( .A(KEYINPUT40), .B(n821), .ZN(G329) );
  NAND2_X1 U909 ( .A1(G2106), .A2(n822), .ZN(G217) );
  NAND2_X1 U910 ( .A1(G15), .A2(G2), .ZN(n823) );
  XNOR2_X1 U911 ( .A(KEYINPUT103), .B(n823), .ZN(n824) );
  NAND2_X1 U912 ( .A1(n824), .A2(G661), .ZN(G259) );
  NAND2_X1 U913 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U914 ( .A1(n826), .A2(n825), .ZN(G188) );
  INV_X1 U916 ( .A(G132), .ZN(G219) );
  INV_X1 U917 ( .A(G120), .ZN(G236) );
  INV_X1 U918 ( .A(G96), .ZN(G221) );
  INV_X1 U919 ( .A(G82), .ZN(G220) );
  INV_X1 U920 ( .A(G69), .ZN(G235) );
  NOR2_X1 U921 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U922 ( .A(n829), .B(KEYINPUT104), .ZN(G325) );
  INV_X1 U923 ( .A(G325), .ZN(G261) );
  XOR2_X1 U924 ( .A(KEYINPUT101), .B(G2446), .Z(n831) );
  XNOR2_X1 U925 ( .A(G2435), .B(G2438), .ZN(n830) );
  XNOR2_X1 U926 ( .A(n831), .B(n830), .ZN(n838) );
  XOR2_X1 U927 ( .A(G2451), .B(G2430), .Z(n833) );
  XNOR2_X1 U928 ( .A(G2454), .B(G2427), .ZN(n832) );
  XNOR2_X1 U929 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U930 ( .A(n834), .B(G2443), .Z(n836) );
  XNOR2_X1 U931 ( .A(G1348), .B(G1341), .ZN(n835) );
  XNOR2_X1 U932 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U933 ( .A(n838), .B(n837), .ZN(n839) );
  NAND2_X1 U934 ( .A1(n839), .A2(G14), .ZN(n840) );
  XOR2_X1 U935 ( .A(KEYINPUT102), .B(n840), .Z(G401) );
  XOR2_X1 U936 ( .A(KEYINPUT109), .B(G1981), .Z(n842) );
  XNOR2_X1 U937 ( .A(G1996), .B(G1991), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U939 ( .A(n843), .B(KEYINPUT41), .Z(n845) );
  XNOR2_X1 U940 ( .A(G1956), .B(G1976), .ZN(n844) );
  XNOR2_X1 U941 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U942 ( .A(G1971), .B(G1961), .Z(n847) );
  XNOR2_X1 U943 ( .A(G1986), .B(G1966), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U945 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U946 ( .A(KEYINPUT110), .B(G2474), .ZN(n850) );
  XNOR2_X1 U947 ( .A(n851), .B(n850), .ZN(G229) );
  XOR2_X1 U948 ( .A(G2678), .B(G2090), .Z(n853) );
  XNOR2_X1 U949 ( .A(G2067), .B(G2072), .ZN(n852) );
  XNOR2_X1 U950 ( .A(n853), .B(n852), .ZN(n863) );
  XOR2_X1 U951 ( .A(KEYINPUT42), .B(KEYINPUT43), .Z(n855) );
  XNOR2_X1 U952 ( .A(G2100), .B(KEYINPUT106), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U954 ( .A(KEYINPUT105), .B(KEYINPUT107), .Z(n857) );
  XNOR2_X1 U955 ( .A(KEYINPUT108), .B(G2096), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U957 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U958 ( .A(G2084), .B(G2078), .ZN(n860) );
  XNOR2_X1 U959 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U960 ( .A(n863), .B(n862), .Z(G227) );
  NAND2_X1 U961 ( .A1(G112), .A2(n889), .ZN(n865) );
  NAND2_X1 U962 ( .A1(G100), .A2(n886), .ZN(n864) );
  NAND2_X1 U963 ( .A1(n865), .A2(n864), .ZN(n870) );
  NAND2_X1 U964 ( .A1(n537), .A2(G124), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n866), .B(KEYINPUT44), .ZN(n868) );
  NAND2_X1 U966 ( .A1(n885), .A2(G136), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n869) );
  NOR2_X1 U968 ( .A1(n870), .A2(n869), .ZN(G162) );
  XNOR2_X1 U969 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n872) );
  XNOR2_X1 U970 ( .A(n998), .B(KEYINPUT111), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n898) );
  NAND2_X1 U972 ( .A1(G118), .A2(n889), .ZN(n874) );
  NAND2_X1 U973 ( .A1(G130), .A2(n537), .ZN(n873) );
  NAND2_X1 U974 ( .A1(n874), .A2(n873), .ZN(n879) );
  NAND2_X1 U975 ( .A1(G142), .A2(n885), .ZN(n876) );
  NAND2_X1 U976 ( .A1(G106), .A2(n886), .ZN(n875) );
  NAND2_X1 U977 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U978 ( .A(KEYINPUT45), .B(n877), .Z(n878) );
  NOR2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n884) );
  XNOR2_X1 U980 ( .A(G160), .B(n880), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U982 ( .A(n884), .B(n883), .Z(n896) );
  NAND2_X1 U983 ( .A1(G139), .A2(n885), .ZN(n888) );
  NAND2_X1 U984 ( .A1(G103), .A2(n886), .ZN(n887) );
  NAND2_X1 U985 ( .A1(n888), .A2(n887), .ZN(n894) );
  NAND2_X1 U986 ( .A1(G115), .A2(n889), .ZN(n891) );
  NAND2_X1 U987 ( .A1(G127), .A2(n537), .ZN(n890) );
  NAND2_X1 U988 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U989 ( .A(KEYINPUT47), .B(n892), .Z(n893) );
  NOR2_X1 U990 ( .A1(n894), .A2(n893), .ZN(n1012) );
  XNOR2_X1 U991 ( .A(G164), .B(n1012), .ZN(n895) );
  XNOR2_X1 U992 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(n901) );
  XNOR2_X1 U994 ( .A(n899), .B(G162), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U996 ( .A1(G37), .A2(n902), .ZN(G395) );
  XOR2_X1 U997 ( .A(KEYINPUT112), .B(n903), .Z(n905) );
  XNOR2_X1 U998 ( .A(G171), .B(G286), .ZN(n904) );
  XNOR2_X1 U999 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1000 ( .A(n906), .B(n937), .Z(n907) );
  XNOR2_X1 U1001 ( .A(n947), .B(n907), .ZN(n908) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n908), .ZN(G397) );
  OR2_X1 U1003 ( .A1(n914), .A2(G401), .ZN(n911) );
  NOR2_X1 U1004 ( .A1(G229), .A2(G227), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n909), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(n911), .A2(n910), .ZN(n913) );
  NOR2_X1 U1007 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1008 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1009 ( .A(G225), .ZN(G308) );
  INV_X1 U1010 ( .A(n914), .ZN(G319) );
  INV_X1 U1011 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1012 ( .A(KEYINPUT54), .B(G34), .ZN(n915) );
  XNOR2_X1 U1013 ( .A(n915), .B(KEYINPUT120), .ZN(n916) );
  XNOR2_X1 U1014 ( .A(G2084), .B(n916), .ZN(n933) );
  XNOR2_X1 U1015 ( .A(G2090), .B(G35), .ZN(n930) );
  XNOR2_X1 U1016 ( .A(G2067), .B(G26), .ZN(n918) );
  XNOR2_X1 U1017 ( .A(G32), .B(G1996), .ZN(n917) );
  NOR2_X1 U1018 ( .A1(n918), .A2(n917), .ZN(n924) );
  XOR2_X1 U1019 ( .A(G25), .B(G1991), .Z(n919) );
  NAND2_X1 U1020 ( .A1(n919), .A2(G28), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(KEYINPUT118), .B(G2072), .ZN(n920) );
  XNOR2_X1 U1022 ( .A(G33), .B(n920), .ZN(n921) );
  NOR2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n927) );
  XOR2_X1 U1025 ( .A(G27), .B(n925), .Z(n926) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1027 ( .A(KEYINPUT53), .B(n928), .ZN(n929) );
  NOR2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(KEYINPUT119), .B(n931), .ZN(n932) );
  NOR2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1031 ( .A(KEYINPUT55), .B(n934), .Z(n935) );
  NOR2_X1 U1032 ( .A1(G29), .A2(n935), .ZN(n936) );
  XOR2_X1 U1033 ( .A(KEYINPUT121), .B(n936), .Z(n991) );
  XNOR2_X1 U1034 ( .A(G16), .B(KEYINPUT56), .ZN(n961) );
  XNOR2_X1 U1035 ( .A(G1348), .B(n937), .ZN(n953) );
  XNOR2_X1 U1036 ( .A(G1971), .B(G303), .ZN(n938) );
  NOR2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n951) );
  XNOR2_X1 U1038 ( .A(n940), .B(G1956), .ZN(n942) );
  XNOR2_X1 U1039 ( .A(G171), .B(G1961), .ZN(n941) );
  NAND2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n946) );
  NAND2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(G1341), .B(n947), .ZN(n948) );
  NOR2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(KEYINPUT122), .B(n954), .ZN(n959) );
  XNOR2_X1 U1048 ( .A(G1966), .B(G168), .ZN(n956) );
  NAND2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(KEYINPUT57), .B(n957), .ZN(n958) );
  NAND2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1052 ( .A1(n961), .A2(n960), .ZN(n987) );
  INV_X1 U1053 ( .A(G16), .ZN(n985) );
  XOR2_X1 U1054 ( .A(G1976), .B(G23), .Z(n963) );
  XOR2_X1 U1055 ( .A(G1971), .B(G22), .Z(n962) );
  NAND2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n965) );
  XNOR2_X1 U1057 ( .A(G24), .B(G1986), .ZN(n964) );
  NOR2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1059 ( .A(KEYINPUT58), .B(n966), .Z(n982) );
  XOR2_X1 U1060 ( .A(G1961), .B(G5), .Z(n977) );
  XOR2_X1 U1061 ( .A(KEYINPUT123), .B(G4), .Z(n968) );
  XNOR2_X1 U1062 ( .A(G1348), .B(KEYINPUT59), .ZN(n967) );
  XNOR2_X1 U1063 ( .A(n968), .B(n967), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(G1341), .B(G19), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(G1981), .B(G6), .ZN(n969) );
  NOR2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(G20), .B(G1956), .ZN(n973) );
  NOR2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1070 ( .A(KEYINPUT60), .B(n975), .ZN(n976) );
  NAND2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(G21), .B(G1966), .ZN(n978) );
  NOR2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1074 ( .A(KEYINPUT124), .B(n980), .Z(n981) );
  NOR2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(KEYINPUT61), .B(n983), .ZN(n984) );
  NAND2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1079 ( .A(KEYINPUT125), .B(n988), .ZN(n989) );
  NAND2_X1 U1080 ( .A1(n989), .A2(G11), .ZN(n990) );
  NOR2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(n992), .B(KEYINPUT126), .ZN(n1023) );
  XNOR2_X1 U1083 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n997) );
  XOR2_X1 U1084 ( .A(G2090), .B(G162), .Z(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1086 ( .A(KEYINPUT51), .B(n995), .Z(n996) );
  XNOR2_X1 U1087 ( .A(n997), .B(n996), .ZN(n1008) );
  NOR2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1005) );
  XNOR2_X1 U1089 ( .A(G160), .B(G2084), .ZN(n1001) );
  NAND2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1093 ( .A(KEYINPUT113), .B(n1006), .Z(n1007) );
  NOR2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1095 ( .A(n1009), .B(KEYINPUT116), .ZN(n1011) );
  NAND2_X1 U1096 ( .A1(n1011), .A2(n1010), .ZN(n1017) );
  XOR2_X1 U1097 ( .A(G2072), .B(n1012), .Z(n1014) );
  XOR2_X1 U1098 ( .A(G164), .B(G2078), .Z(n1013) );
  NOR2_X1 U1099 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1100 ( .A(KEYINPUT50), .B(n1015), .Z(n1016) );
  NOR2_X1 U1101 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1102 ( .A(KEYINPUT52), .B(n1018), .Z(n1019) );
  NOR2_X1 U1103 ( .A1(KEYINPUT55), .A2(n1019), .ZN(n1020) );
  XNOR2_X1 U1104 ( .A(KEYINPUT117), .B(n1020), .ZN(n1021) );
  NAND2_X1 U1105 ( .A1(n1021), .A2(G29), .ZN(n1022) );
  NAND2_X1 U1106 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1024), .Z(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

