//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1189,
    new_n1190, new_n1191, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  OAI21_X1  g0010(.A(G50), .B1(G58), .B2(G68), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  INV_X1    g0024(.A(G107), .ZN(new_n225));
  INV_X1    g0025(.A(G264), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n223), .B1(new_n202), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n207), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n210), .B(new_n216), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT64), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n234), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT65), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  XNOR2_X1  g0047(.A(KEYINPUT3), .B(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n248), .A2(G223), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G87), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n248), .A2(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(G226), .ZN(new_n253));
  OAI211_X1 g0053(.A(new_n250), .B(new_n251), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G274), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(G41), .B2(G45), .ZN(new_n259));
  NOR3_X1   g0059(.A1(new_n255), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n259), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n255), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n260), .B1(G232), .B2(new_n262), .ZN(new_n263));
  AND3_X1   g0063(.A1(new_n256), .A2(G190), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G200), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n265), .B1(new_n256), .B2(new_n263), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT7), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n248), .A2(new_n268), .A3(G20), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(KEYINPUT7), .B1(new_n274), .B2(new_n214), .ZN(new_n275));
  OAI21_X1  g0075(.A(G68), .B1(new_n269), .B2(new_n275), .ZN(new_n276));
  AND2_X1   g0076(.A1(G58), .A2(G68), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G58), .A2(G68), .ZN(new_n278));
  OAI211_X1 g0078(.A(KEYINPUT73), .B(G20), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G159), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(G58), .B(G68), .ZN(new_n283));
  AOI21_X1  g0083(.A(KEYINPUT73), .B1(new_n283), .B2(G20), .ZN(new_n284));
  OAI21_X1  g0084(.A(KEYINPUT74), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(G20), .B1(new_n277), .B2(new_n278), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT73), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT74), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n288), .A2(new_n289), .A3(new_n281), .A4(new_n279), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n276), .A2(new_n285), .A3(KEYINPUT16), .A4(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n213), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT16), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n268), .B1(new_n248), .B2(G20), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n274), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n218), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n288), .A2(new_n281), .A3(new_n279), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n294), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n291), .A2(new_n293), .A3(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT8), .ZN(new_n301));
  INV_X1    g0101(.A(G58), .ZN(new_n302));
  OR3_X1    g0102(.A1(new_n301), .A2(new_n302), .A3(KEYINPUT67), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n301), .B1(new_n302), .B2(KEYINPUT67), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G13), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n306), .A2(G1), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G20), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n293), .B1(new_n258), .B2(G20), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n309), .B1(new_n310), .B2(new_n305), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n267), .A2(new_n300), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT17), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT17), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(KEYINPUT77), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT77), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n312), .A2(new_n315), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n300), .A2(new_n311), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT17), .B1(new_n321), .B2(new_n267), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n318), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n317), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT76), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT18), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT75), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n300), .A2(new_n327), .A3(new_n311), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n327), .B1(new_n300), .B2(new_n311), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G169), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(new_n256), .B2(new_n263), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n256), .A2(new_n263), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n332), .B1(G179), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n326), .B1(new_n330), .B2(new_n335), .ZN(new_n336));
  NOR4_X1   g0136(.A1(new_n328), .A2(new_n329), .A3(KEYINPUT18), .A4(new_n334), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n325), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n330), .A2(new_n326), .A3(new_n335), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n320), .A2(KEYINPUT75), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n300), .A2(new_n327), .A3(new_n311), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(new_n341), .A3(new_n335), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT18), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n339), .A2(new_n343), .A3(KEYINPUT76), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n324), .B1(new_n338), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n214), .A2(G33), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n305), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G150), .ZN(new_n348));
  INV_X1    g0148(.A(new_n280), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n348), .A2(new_n349), .B1(new_n201), .B2(new_n214), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n293), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n310), .A2(G50), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n351), .B(new_n352), .C1(G50), .C2(new_n308), .ZN(new_n353));
  OR2_X1    g0153(.A1(new_n353), .A2(KEYINPUT9), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(KEYINPUT9), .ZN(new_n355));
  INV_X1    g0155(.A(new_n255), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n259), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(new_n253), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n274), .A2(G1698), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G222), .ZN(new_n360));
  XNOR2_X1  g0160(.A(KEYINPUT66), .B(G223), .ZN(new_n361));
  OAI221_X1 g0161(.A(new_n360), .B1(new_n202), .B2(new_n248), .C1(new_n252), .C2(new_n361), .ZN(new_n362));
  AOI211_X1 g0162(.A(new_n260), .B(new_n358), .C1(new_n362), .C2(new_n255), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n354), .A2(new_n355), .B1(G190), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT10), .B1(new_n364), .B2(KEYINPUT69), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n364), .B1(new_n265), .B2(new_n363), .ZN(new_n366));
  XOR2_X1   g0166(.A(new_n365), .B(new_n366), .Z(new_n367));
  INV_X1    g0167(.A(G179), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n369), .B(new_n353), .C1(G169), .C2(new_n363), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n248), .A2(G232), .A3(new_n249), .ZN(new_n372));
  OAI221_X1 g0172(.A(new_n372), .B1(new_n225), .B2(new_n248), .C1(new_n252), .C2(new_n219), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n255), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n260), .B1(G244), .B2(new_n262), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n331), .ZN(new_n377));
  INV_X1    g0177(.A(new_n293), .ZN(new_n378));
  XNOR2_X1  g0178(.A(KEYINPUT15), .B(G87), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n379), .A2(KEYINPUT68), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(KEYINPUT68), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OR2_X1    g0182(.A1(new_n382), .A2(new_n346), .ZN(new_n383));
  XNOR2_X1  g0183(.A(KEYINPUT8), .B(G58), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n385), .A2(new_n280), .B1(G20), .B2(G77), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n378), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n310), .A2(G77), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(G77), .B2(new_n308), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n377), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n376), .A2(G179), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n387), .A2(new_n389), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n376), .A2(G200), .ZN(new_n395));
  INV_X1    g0195(.A(G190), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n394), .B(new_n395), .C1(new_n396), .C2(new_n376), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n371), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT71), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n219), .B1(new_n357), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n262), .A2(KEYINPUT71), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n260), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n359), .A2(KEYINPUT70), .A3(G226), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT70), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n248), .A2(new_n249), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n405), .B1(new_n406), .B2(new_n253), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n248), .A2(G232), .A3(G1698), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G97), .ZN(new_n409));
  AND4_X1   g0209(.A1(new_n404), .A2(new_n407), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n403), .B1(new_n410), .B2(new_n356), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT13), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n411), .B(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT14), .B1(new_n413), .B2(new_n331), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(G179), .ZN(new_n415));
  XNOR2_X1  g0215(.A(new_n411), .B(KEYINPUT13), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT14), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n416), .A2(new_n417), .A3(G169), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n414), .A2(new_n415), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n310), .A2(G68), .ZN(new_n420));
  XOR2_X1   g0220(.A(new_n420), .B(KEYINPUT72), .Z(new_n421));
  INV_X1    g0221(.A(G50), .ZN(new_n422));
  OAI22_X1  g0222(.A1(new_n349), .A2(new_n422), .B1(new_n214), .B2(G68), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n346), .A2(new_n202), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n293), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT11), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n308), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n218), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT12), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n425), .A2(new_n426), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n421), .A2(new_n427), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n419), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n416), .A2(G200), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n413), .A2(G190), .ZN(new_n435));
  INV_X1    g0235(.A(new_n432), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  AND4_X1   g0237(.A1(new_n345), .A2(new_n399), .A3(new_n433), .A4(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G33), .A2(G116), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(new_n252), .B2(new_n224), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n406), .A2(new_n219), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n255), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G45), .ZN(new_n443));
  OAI21_X1  g0243(.A(G250), .B1(new_n443), .B2(G1), .ZN(new_n444));
  OR3_X1    g0244(.A1(new_n255), .A2(new_n444), .A3(KEYINPUT82), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT82), .B1(new_n255), .B2(new_n444), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n255), .A2(new_n257), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n443), .A2(G1), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n445), .A2(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n442), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n368), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n331), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n258), .A2(G33), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n378), .A2(new_n308), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT78), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT78), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n378), .A2(new_n308), .A3(new_n458), .A4(new_n455), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n382), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n248), .A2(new_n214), .A3(G68), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT19), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n214), .B1(new_n409), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(G87), .B2(new_n205), .ZN(new_n466));
  INV_X1    g0266(.A(G97), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n464), .B1(new_n346), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n463), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n428), .A2(new_n382), .B1(new_n469), .B2(new_n293), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n462), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(KEYINPUT83), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT83), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n473), .B1(new_n462), .B2(new_n470), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n454), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n248), .A2(G257), .A3(G1698), .ZN(new_n476));
  XNOR2_X1  g0276(.A(KEYINPUT85), .B(G294), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G33), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n476), .B(new_n478), .C1(new_n406), .C2(new_n221), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n255), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT5), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G41), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n448), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT80), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n448), .A2(KEYINPUT80), .A3(new_n482), .ZN(new_n486));
  INV_X1    g0286(.A(G41), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT5), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n485), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n489), .A2(G264), .A3(new_n356), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n480), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n485), .A2(new_n486), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT81), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n485), .A2(KEYINPUT81), .A3(new_n486), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n494), .A2(new_n447), .A3(new_n495), .A4(new_n488), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G200), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n248), .A2(new_n214), .A3(G87), .ZN(new_n499));
  XNOR2_X1  g0299(.A(new_n499), .B(KEYINPUT22), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT24), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT23), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n214), .B2(G107), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n225), .A2(KEYINPUT23), .A3(G20), .ZN(new_n504));
  INV_X1    g0304(.A(new_n439), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n503), .A2(new_n504), .B1(new_n505), .B2(new_n214), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n500), .A2(new_n501), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n501), .B1(new_n500), .B2(new_n506), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n293), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n460), .A2(G107), .ZN(new_n511));
  XOR2_X1   g0311(.A(KEYINPUT84), .B(KEYINPUT25), .Z(new_n512));
  INV_X1    g0312(.A(KEYINPUT84), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT25), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n307), .A2(G20), .A3(new_n225), .ZN(new_n515));
  MUX2_X1   g0315(.A(new_n512), .B(new_n514), .S(new_n515), .Z(new_n516));
  NAND2_X1  g0316(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n491), .A2(G190), .A3(new_n496), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n498), .A2(new_n510), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n497), .A2(new_n331), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n491), .A2(new_n368), .A3(new_n496), .ZN(new_n522));
  INV_X1    g0322(.A(new_n509), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n378), .B1(new_n523), .B2(new_n507), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n521), .B(new_n522), .C1(new_n524), .C2(new_n517), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n451), .A2(new_n265), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n457), .A2(new_n459), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n470), .B1(new_n220), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n451), .A2(G190), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n475), .A2(new_n520), .A3(new_n525), .A4(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n248), .A2(G257), .A3(new_n249), .ZN(new_n533));
  INV_X1    g0333(.A(G303), .ZN(new_n534));
  OAI221_X1 g0334(.A(new_n533), .B1(new_n534), .B2(new_n248), .C1(new_n252), .C2(new_n226), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n255), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n489), .A2(G270), .A3(new_n356), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n496), .A2(new_n536), .A3(G179), .A4(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(G116), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n428), .A2(new_n540), .ZN(new_n541));
  OR2_X1    g0341(.A1(new_n456), .A2(new_n540), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G283), .ZN(new_n543));
  XNOR2_X1  g0343(.A(new_n543), .B(KEYINPUT79), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n544), .B(new_n214), .C1(G33), .C2(new_n467), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n378), .B1(G20), .B2(new_n540), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n545), .A2(KEYINPUT20), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT20), .B1(new_n545), .B2(new_n546), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n541), .B(new_n542), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n539), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n496), .A2(new_n536), .A3(new_n537), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n549), .A2(new_n551), .A3(KEYINPUT21), .A4(G169), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n549), .A2(new_n551), .A3(G169), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT21), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n551), .A2(G200), .ZN(new_n557));
  INV_X1    g0357(.A(new_n549), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n496), .A2(new_n536), .A3(G190), .A4(new_n537), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n553), .A2(new_n556), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n225), .A2(KEYINPUT6), .A3(G97), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n467), .A2(new_n225), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n563), .A2(new_n204), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n562), .B1(new_n564), .B2(KEYINPUT6), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n565), .A2(G20), .B1(G77), .B2(new_n280), .ZN(new_n566));
  OAI21_X1  g0366(.A(G107), .B1(new_n269), .B2(new_n275), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n378), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n428), .A2(new_n467), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n527), .B2(new_n467), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n248), .A2(G250), .A3(G1698), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n248), .A2(G244), .A3(new_n249), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT4), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n544), .B(new_n573), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT4), .B1(new_n359), .B2(G244), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n255), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n489), .A2(G257), .A3(new_n356), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n496), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n331), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n572), .B(new_n581), .C1(G179), .C2(new_n580), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(G200), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n583), .B(new_n571), .C1(new_n396), .C2(new_n580), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n532), .A2(new_n561), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n438), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g0387(.A(new_n587), .B(KEYINPUT86), .ZN(G372));
  NAND2_X1  g0388(.A1(new_n529), .A2(KEYINPUT87), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT87), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(new_n526), .B2(new_n528), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n591), .A3(new_n530), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n592), .A2(new_n475), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n582), .A2(new_n584), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n553), .A2(new_n525), .A3(new_n556), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n520), .A4(new_n595), .ZN(new_n596));
  XNOR2_X1  g0396(.A(new_n471), .B(KEYINPUT83), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n597), .A2(new_n454), .B1(new_n530), .B2(new_n529), .ZN(new_n598));
  INV_X1    g0398(.A(new_n582), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n600), .A2(KEYINPUT88), .A3(KEYINPUT26), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n596), .A2(new_n475), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(KEYINPUT26), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT88), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n592), .A2(new_n599), .A3(new_n475), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT26), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n603), .A2(new_n604), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n602), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n438), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n437), .ZN(new_n611));
  AOI211_X1 g0411(.A(new_n611), .B(new_n324), .C1(new_n433), .C2(new_n393), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n321), .A2(new_n334), .ZN(new_n613));
  XNOR2_X1  g0413(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n614));
  XNOR2_X1  g0414(.A(new_n613), .B(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n367), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n616), .A2(new_n370), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n610), .A2(new_n617), .ZN(G369));
  NAND2_X1  g0418(.A1(new_n553), .A2(new_n556), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n307), .A2(new_n214), .ZN(new_n620));
  OR2_X1    g0420(.A1(new_n620), .A2(KEYINPUT27), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(KEYINPUT27), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n621), .A2(G213), .A3(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(G343), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n558), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n619), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n628), .B1(new_n561), .B2(new_n627), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n629), .A2(G330), .ZN(new_n630));
  INV_X1    g0430(.A(new_n520), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n626), .B1(new_n510), .B2(new_n518), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n525), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n525), .A2(new_n625), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g0437(.A(new_n637), .B(KEYINPUT90), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n625), .B1(new_n553), .B2(new_n556), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n635), .B1(new_n633), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n639), .A2(new_n641), .ZN(G399));
  INV_X1    g0442(.A(new_n208), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n643), .A2(G41), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(G1), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(new_n211), .B2(new_n645), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n648), .B(KEYINPUT28), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT29), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n609), .A2(new_n650), .A3(new_n626), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n605), .A2(KEYINPUT26), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n600), .A2(new_n606), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n596), .A2(new_n475), .A3(new_n652), .A4(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n650), .B1(new_n654), .B2(new_n626), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n538), .A2(new_n580), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n442), .A2(new_n480), .A3(new_n449), .A4(new_n490), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT91), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n658), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT30), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT92), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n450), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n442), .A2(new_n449), .A3(KEYINPUT92), .ZN(new_n667));
  AND4_X1   g0467(.A1(new_n551), .A2(new_n666), .A3(new_n580), .A4(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(G179), .B1(new_n491), .B2(new_n496), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n663), .A2(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n658), .B(KEYINPUT30), .C1(new_n661), .C2(new_n662), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n672), .A2(KEYINPUT31), .A3(new_n625), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT93), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT93), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n626), .B1(new_n670), .B2(new_n671), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT31), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n674), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(KEYINPUT94), .B1(new_n586), .B2(new_n626), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n525), .A2(new_n520), .ZN(new_n680));
  AND4_X1   g0480(.A1(new_n556), .A2(new_n560), .A3(new_n550), .A4(new_n552), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n680), .A2(new_n594), .A3(new_n681), .A4(new_n598), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT94), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n682), .A2(new_n683), .A3(new_n625), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(G330), .B1(new_n678), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT95), .B1(new_n657), .B2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n625), .B1(new_n602), .B2(new_n608), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n655), .B1(new_n689), .B2(new_n650), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT95), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(new_n691), .A3(new_n686), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n649), .B1(new_n693), .B2(G1), .ZN(G364));
  NOR2_X1   g0494(.A1(new_n629), .A2(G330), .ZN(new_n695));
  XOR2_X1   g0495(.A(new_n695), .B(KEYINPUT96), .Z(new_n696));
  NOR2_X1   g0496(.A1(new_n306), .A2(G20), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n258), .B1(new_n697), .B2(G45), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OR3_X1    g0499(.A1(new_n644), .A2(new_n699), .A3(KEYINPUT97), .ZN(new_n700));
  OAI21_X1  g0500(.A(KEYINPUT97), .B1(new_n644), .B2(new_n699), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n630), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n696), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n213), .B1(G20), .B2(new_n331), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n396), .A2(G179), .A3(G200), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(new_n214), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n214), .A2(new_n368), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(G200), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n396), .ZN(new_n713));
  XNOR2_X1  g0513(.A(KEYINPUT99), .B(G326), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n477), .A2(new_n710), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT100), .ZN(new_n717));
  NOR2_X1   g0517(.A1(G190), .A2(G200), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n711), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(G311), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n214), .A2(G179), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n718), .ZN(new_n722));
  INV_X1    g0522(.A(G329), .ZN(new_n723));
  OAI22_X1  g0523(.A1(new_n719), .A2(new_n720), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n711), .A2(G190), .A3(new_n265), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI211_X1 g0526(.A(new_n248), .B(new_n724), .C1(G322), .C2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n712), .A2(G190), .ZN(new_n728));
  INV_X1    g0528(.A(G317), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT33), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n729), .A2(KEYINPUT33), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n728), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n721), .A2(G190), .A3(G200), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n721), .A2(new_n396), .A3(G200), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n734), .A2(G303), .B1(new_n736), .B2(G283), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n717), .A2(new_n727), .A3(new_n732), .A4(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n722), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G159), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(KEYINPUT32), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n728), .A2(G68), .B1(new_n736), .B2(G107), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n710), .A2(G97), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n733), .A2(new_n220), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n740), .A2(KEYINPUT32), .ZN(new_n747));
  INV_X1    g0547(.A(new_n713), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n747), .B1(new_n422), .B2(new_n748), .ZN(new_n749));
  OAI221_X1 g0549(.A(new_n248), .B1(new_n719), .B2(new_n202), .C1(new_n302), .C2(new_n725), .ZN(new_n750));
  OR4_X1    g0550(.A1(new_n741), .A2(new_n746), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n707), .B1(new_n738), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G13), .A2(G33), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n706), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n643), .A2(new_n274), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT98), .ZN(new_n758));
  INV_X1    g0558(.A(G355), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n758), .A2(new_n759), .B1(G116), .B2(new_n208), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n643), .A2(new_n248), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(G45), .B2(new_n211), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n762), .B1(new_n246), .B2(G45), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n702), .B(new_n752), .C1(new_n756), .C2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n755), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n765), .B1(new_n629), .B2(new_n766), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n705), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(G396));
  OAI21_X1  g0569(.A(new_n397), .B1(new_n394), .B2(new_n626), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(new_n393), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n392), .A2(new_n626), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n689), .B(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n703), .B1(new_n775), .B2(new_n686), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(new_n686), .B2(new_n775), .ZN(new_n777));
  INV_X1    g0577(.A(G283), .ZN(new_n778));
  INV_X1    g0578(.A(new_n728), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n778), .A2(new_n779), .B1(new_n748), .B2(new_n534), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(G107), .B2(new_n734), .ZN(new_n781));
  INV_X1    g0581(.A(G294), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n725), .A2(new_n782), .B1(new_n722), .B2(new_n720), .ZN(new_n783));
  INV_X1    g0583(.A(new_n719), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n248), .B(new_n783), .C1(G116), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n736), .A2(G87), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n781), .A2(new_n743), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n726), .A2(G143), .B1(new_n784), .B2(G159), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n713), .A2(G137), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n788), .B(new_n789), .C1(new_n348), .C2(new_n779), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT34), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n736), .A2(G68), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n274), .B1(new_n739), .B2(G132), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n710), .A2(G58), .B1(new_n734), .B2(G50), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n792), .A2(new_n793), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n790), .A2(new_n791), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n787), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n706), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n706), .A2(new_n753), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n702), .B1(new_n202), .B2(new_n800), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT101), .Z(new_n802));
  OAI211_X1 g0602(.A(new_n799), .B(new_n802), .C1(new_n774), .C2(new_n754), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n777), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(G384));
  OR2_X1    g0605(.A1(new_n565), .A2(KEYINPUT35), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n565), .A2(KEYINPUT35), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n806), .A2(G116), .A3(new_n215), .A4(new_n807), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT36), .Z(new_n809));
  OAI211_X1 g0609(.A(new_n212), .B(G77), .C1(new_n302), .C2(new_n218), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n422), .A2(G68), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n258), .B(G13), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT38), .ZN(new_n814));
  INV_X1    g0614(.A(new_n311), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n291), .A2(new_n293), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n276), .A2(new_n285), .A3(new_n290), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n294), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n815), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(new_n623), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n338), .A2(new_n344), .ZN(new_n822));
  INV_X1    g0622(.A(new_n324), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n312), .B1(new_n819), .B2(new_n623), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n819), .A2(new_n334), .ZN(new_n826));
  OAI21_X1  g0626(.A(KEYINPUT37), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  XOR2_X1   g0627(.A(KEYINPUT102), .B(KEYINPUT37), .Z(new_n828));
  AND2_X1   g0628(.A1(new_n312), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n623), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n340), .A2(new_n341), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n829), .A2(new_n342), .A3(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT103), .ZN(new_n833));
  AND3_X1   g0633(.A1(new_n827), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n833), .B1(new_n827), .B2(new_n832), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n814), .B1(new_n824), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT104), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n827), .A2(new_n832), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(KEYINPUT103), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n827), .A2(new_n832), .A3(new_n833), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n842), .B(KEYINPUT38), .C1(new_n345), .C2(new_n821), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n837), .A2(new_n838), .A3(new_n843), .ZN(new_n844));
  OAI211_X1 g0644(.A(KEYINPUT104), .B(new_n814), .C1(new_n824), .C2(new_n836), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n433), .B(new_n437), .C1(new_n436), .C2(new_n626), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n432), .B(new_n625), .C1(new_n611), .C2(new_n419), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n608), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n596), .A2(new_n475), .A3(new_n601), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n626), .B(new_n774), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n850), .B1(new_n853), .B2(new_n772), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n846), .A2(new_n854), .B1(new_n615), .B2(new_n623), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n844), .A2(KEYINPUT39), .A3(new_n845), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT105), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n844), .A2(KEYINPUT105), .A3(KEYINPUT39), .A4(new_n845), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT107), .ZN(new_n860));
  NOR3_X1   g0660(.A1(new_n615), .A2(new_n322), .A3(new_n319), .ZN(new_n861));
  INV_X1    g0661(.A(new_n832), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n613), .A2(new_n313), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n828), .B1(new_n863), .B2(new_n831), .ZN(new_n864));
  OAI22_X1  g0664(.A1(new_n861), .A2(new_n831), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  XNOR2_X1  g0665(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n843), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n860), .B1(new_n868), .B2(KEYINPUT39), .ZN(new_n869));
  INV_X1    g0669(.A(new_n868), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT39), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n870), .A2(KEYINPUT107), .A3(new_n871), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n858), .A2(new_n859), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n419), .A2(new_n432), .A3(new_n626), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n855), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n657), .A2(new_n438), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n617), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n875), .B(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(G330), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n673), .B(new_n677), .C1(new_n679), .C2(new_n684), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n773), .B1(new_n847), .B2(new_n848), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n880), .A2(new_n881), .A3(KEYINPUT40), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT108), .B1(new_n870), .B2(new_n882), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n880), .A2(new_n881), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT108), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n884), .A2(new_n885), .A3(KEYINPUT40), .A4(new_n868), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n884), .A2(new_n845), .A3(new_n844), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT40), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n438), .A2(new_n880), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n879), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n892), .B2(new_n891), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n878), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n258), .B2(new_n697), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n878), .A2(new_n894), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n813), .B1(new_n896), .B2(new_n897), .ZN(G367));
  INV_X1    g0698(.A(new_n693), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n636), .B(new_n640), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(new_n630), .ZN(new_n901));
  INV_X1    g0701(.A(new_n692), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n691), .B1(new_n690), .B2(new_n686), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT110), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT110), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n693), .A2(new_n906), .A3(new_n901), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT44), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n594), .B1(new_n571), .B2(new_n626), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n599), .A2(new_n625), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n908), .B1(new_n641), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n641), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(new_n911), .A3(KEYINPUT44), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n641), .A2(KEYINPUT45), .A3(new_n912), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT45), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n914), .B2(new_n911), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n639), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n639), .A2(new_n921), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n905), .A2(new_n907), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(KEYINPUT111), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT111), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n905), .A2(new_n907), .A3(new_n927), .A4(new_n924), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n899), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n644), .B(KEYINPUT41), .Z(new_n930));
  OAI21_X1  g0730(.A(new_n698), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n912), .A2(new_n636), .A3(new_n640), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT42), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n582), .B1(new_n909), .B2(new_n525), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n933), .B1(new_n626), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n528), .A2(new_n625), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n593), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n475), .B2(new_n936), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n935), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT109), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n935), .A2(new_n939), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n941), .A2(new_n942), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n639), .A2(new_n911), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n946), .B(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n931), .A2(new_n948), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n938), .A2(new_n766), .ZN(new_n950));
  INV_X1    g0750(.A(new_n756), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(new_n233), .B2(new_n761), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n208), .B2(new_n382), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n703), .A2(new_n953), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n728), .A2(G159), .B1(new_n734), .B2(G58), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n218), .B2(new_n709), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n713), .A2(G143), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n202), .B2(new_n735), .ZN(new_n958));
  XOR2_X1   g0758(.A(KEYINPUT113), .B(G137), .Z(new_n959));
  OAI21_X1  g0759(.A(new_n248), .B1(new_n959), .B2(new_n722), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n725), .A2(new_n348), .B1(new_n719), .B2(new_n422), .ZN(new_n961));
  NOR4_X1   g0761(.A1(new_n956), .A2(new_n958), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n728), .A2(new_n477), .B1(new_n736), .B2(G97), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n963), .B1(new_n225), .B2(new_n709), .C1(new_n720), .C2(new_n748), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n274), .B1(new_n719), .B2(new_n778), .ZN(new_n965));
  XNOR2_X1  g0765(.A(KEYINPUT112), .B(G317), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n725), .A2(new_n534), .B1(new_n722), .B2(new_n966), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n734), .A2(G116), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT46), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n962), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT47), .Z(new_n972));
  AOI21_X1  g0772(.A(new_n954), .B1(new_n972), .B2(new_n706), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n950), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n949), .A2(new_n974), .ZN(G387));
  NAND2_X1  g0775(.A1(new_n905), .A2(new_n907), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n976), .B(new_n644), .C1(new_n693), .C2(new_n901), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n901), .A2(new_n699), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT114), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n761), .B1(new_n238), .B2(new_n443), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n646), .B2(new_n758), .ZN(new_n981));
  OR3_X1    g0781(.A1(new_n384), .A2(KEYINPUT50), .A3(G50), .ZN(new_n982));
  OAI21_X1  g0782(.A(KEYINPUT50), .B1(new_n384), .B2(G50), .ZN(new_n983));
  AOI21_X1  g0783(.A(G45), .B1(G68), .B2(G77), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n982), .A2(new_n646), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n981), .A2(new_n985), .B1(new_n225), .B2(new_n643), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n703), .B1(new_n986), .B2(new_n951), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n636), .A2(new_n766), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n725), .A2(new_n422), .B1(new_n722), .B2(new_n348), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n274), .B(new_n989), .C1(G68), .C2(new_n784), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n734), .A2(G77), .B1(new_n736), .B2(G97), .ZN(new_n991));
  INV_X1    g0791(.A(new_n305), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n992), .A2(new_n728), .B1(new_n713), .B2(G159), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n382), .A2(new_n709), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n990), .A2(new_n991), .A3(new_n993), .A4(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n966), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n726), .A2(new_n997), .B1(new_n784), .B2(G303), .ZN(new_n998));
  INV_X1    g0798(.A(G322), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n998), .B1(new_n779), .B2(new_n720), .C1(new_n999), .C2(new_n748), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT48), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n710), .A2(G283), .B1(new_n734), .B2(new_n477), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT49), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(KEYINPUT115), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n248), .B1(new_n739), .B2(new_n715), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1007), .B(new_n1008), .C1(new_n540), .C2(new_n735), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1006), .A2(KEYINPUT115), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n996), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n987), .B(new_n988), .C1(new_n1011), .C2(new_n706), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n979), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n977), .A2(new_n1013), .ZN(G393));
  OR2_X1    g0814(.A1(new_n924), .A2(KEYINPUT116), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n924), .A2(KEYINPUT116), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1015), .A2(new_n1016), .A3(new_n699), .ZN(new_n1017));
  NOR3_X1   g0817(.A1(new_n243), .A2(new_n643), .A3(new_n248), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n756), .B1(new_n467), .B2(new_n208), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n703), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G317), .A2(new_n713), .B1(new_n726), .B2(G311), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT52), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n274), .B1(new_n722), .B2(new_n999), .C1(new_n782), .C2(new_n719), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n779), .A2(new_n534), .B1(new_n735), .B2(new_n225), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n709), .A2(new_n540), .B1(new_n733), .B2(new_n778), .ZN(new_n1025));
  OR4_X1    g0825(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G150), .A2(new_n713), .B1(new_n726), .B2(G159), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT117), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT51), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n274), .B1(new_n739), .B2(G143), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1030), .B(new_n786), .C1(new_n218), .C2(new_n733), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT118), .Z(new_n1032));
  NOR2_X1   g0832(.A1(new_n719), .A2(new_n384), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n709), .A2(new_n202), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n1033), .B(new_n1034), .C1(G50), .C2(new_n728), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1026), .B1(new_n1029), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1020), .B1(new_n1037), .B2(new_n706), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n912), .B2(new_n766), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1017), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n926), .A2(new_n928), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n924), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n645), .B1(new_n976), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1040), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(G390));
  INV_X1    g0845(.A(new_n874), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n654), .A2(new_n626), .A3(new_n771), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n772), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1046), .B1(new_n1048), .B2(new_n849), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n868), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  NOR3_X1   g0851(.A1(new_n686), .A2(new_n773), .A3(new_n850), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n854), .A2(new_n1046), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1051), .B(new_n1052), .C1(new_n873), .C2(new_n1053), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n880), .A2(G330), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n881), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n858), .A2(new_n859), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n872), .A2(new_n869), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1057), .A2(new_n1058), .A3(new_n1053), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1056), .B1(new_n1059), .B2(new_n1050), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1054), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n873), .A2(new_n753), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n734), .A2(G150), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT53), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G159), .A2(new_n710), .B1(new_n713), .B2(G128), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n422), .B2(new_n735), .C1(new_n779), .C2(new_n959), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n274), .B1(new_n739), .B2(G125), .ZN(new_n1067));
  INV_X1    g0867(.A(G132), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(KEYINPUT54), .B(G143), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1067), .B1(new_n1068), .B2(new_n725), .C1(new_n719), .C2(new_n1069), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1064), .A2(new_n1066), .A3(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n779), .A2(new_n225), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1034), .B(new_n1072), .C1(G283), .C2(new_n713), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n719), .A2(new_n467), .B1(new_n722), .B2(new_n782), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n248), .B(new_n1074), .C1(G116), .C2(new_n726), .ZN(new_n1075));
  AND3_X1   g0875(.A1(new_n1075), .A2(new_n745), .A3(new_n793), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1071), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1077), .A2(new_n707), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n702), .B(new_n1078), .C1(new_n305), .C2(new_n800), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1061), .A2(new_n699), .B1(new_n1062), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT120), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1055), .A2(new_n774), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1048), .B1(new_n1082), .B2(new_n850), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1052), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n850), .B1(new_n686), .B2(new_n773), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n1056), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n853), .A2(new_n772), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1083), .A2(new_n1084), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n438), .A2(new_n1055), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n876), .A2(new_n617), .A3(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(KEYINPUT119), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n645), .B1(new_n1061), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1088), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1090), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g0895(.A(KEYINPUT119), .B(new_n1095), .C1(new_n1054), .C2(new_n1060), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1081), .B1(new_n1092), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1059), .A2(new_n1050), .A3(new_n1084), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1051), .B1(new_n873), .B2(new_n1053), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1091), .B(new_n1098), .C1(new_n1099), .C2(new_n1056), .ZN(new_n1100));
  AND4_X1   g0900(.A1(new_n1081), .A2(new_n1096), .A3(new_n644), .A4(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1080), .B1(new_n1097), .B2(new_n1101), .ZN(G378));
  NAND3_X1  g0902(.A1(new_n887), .A2(new_n890), .A3(G330), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n353), .A2(new_n830), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n371), .B(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1105), .B(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1103), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n887), .A2(new_n1107), .A3(new_n890), .A4(G330), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n875), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n1046), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1114), .A2(new_n1109), .A3(new_n855), .A4(new_n1110), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1108), .A2(new_n753), .ZN(new_n1117));
  AOI211_X1 g0917(.A(G41), .B(new_n248), .C1(new_n739), .C2(G283), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1118), .B1(new_n302), .B2(new_n735), .C1(new_n202), .C2(new_n733), .ZN(new_n1119));
  XOR2_X1   g0919(.A(new_n1119), .B(KEYINPUT121), .Z(new_n1120));
  OAI22_X1  g0920(.A1(new_n709), .A2(new_n218), .B1(new_n725), .B2(new_n225), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n467), .A2(new_n779), .B1(new_n748), .B2(new_n540), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n1121), .B(new_n1122), .C1(new_n461), .C2(new_n784), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT58), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(G33), .A2(G41), .ZN(new_n1126));
  AOI211_X1 g0926(.A(G50), .B(new_n1126), .C1(new_n274), .C2(new_n487), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n713), .A2(G125), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n779), .B2(new_n1068), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(G150), .B2(new_n710), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n726), .A2(G128), .B1(new_n784), .B2(G137), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1130), .B(new_n1131), .C1(new_n733), .C2(new_n1069), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n1132), .A2(KEYINPUT59), .ZN(new_n1133));
  INV_X1    g0933(.A(G124), .ZN(new_n1134));
  INV_X1    g0934(.A(G159), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1126), .B1(new_n722), .B2(new_n1134), .C1(new_n1135), .C2(new_n735), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n1132), .B2(KEYINPUT59), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1127), .B1(new_n1133), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n707), .B1(new_n1125), .B2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT122), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n702), .B(new_n1140), .C1(new_n422), .C2(new_n800), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1116), .A2(new_n699), .B1(new_n1117), .B2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1098), .B(new_n1093), .C1(new_n1099), .C2(new_n1056), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n1094), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1144), .A2(KEYINPUT57), .A3(new_n1116), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n644), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1143), .A2(new_n1094), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1147), .A2(KEYINPUT57), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1142), .B1(new_n1146), .B2(new_n1148), .ZN(G375));
  INV_X1    g0949(.A(new_n930), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1095), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n850), .A2(new_n753), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT123), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(G50), .A2(new_n710), .B1(new_n713), .B2(G132), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n1135), .B2(new_n733), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n248), .B1(new_n725), .B2(new_n959), .ZN(new_n1157));
  INV_X1    g0957(.A(G128), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n719), .A2(new_n348), .B1(new_n722), .B2(new_n1158), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n779), .A2(new_n1069), .B1(new_n302), .B2(new_n735), .ZN(new_n1160));
  NOR4_X1   g0960(.A1(new_n1156), .A2(new_n1157), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n248), .B1(new_n739), .B2(G303), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1162), .B1(new_n225), .B2(new_n719), .C1(new_n778), .C2(new_n725), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n540), .A2(new_n779), .B1(new_n748), .B2(new_n782), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n202), .A2(new_n735), .B1(new_n733), .B2(new_n467), .ZN(new_n1165));
  NOR4_X1   g0965(.A1(new_n1163), .A2(new_n1164), .A3(new_n994), .A4(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n706), .B1(new_n1161), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n702), .B1(new_n218), .B2(new_n800), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1154), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n1088), .B2(new_n698), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1152), .A2(new_n1171), .ZN(G381));
  NOR3_X1   g0972(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT124), .ZN(new_n1174));
  NOR3_X1   g0974(.A1(new_n1174), .A2(G390), .A3(G381), .ZN(new_n1175));
  INV_X1    g0975(.A(G387), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1117), .A2(new_n1141), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1116), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1177), .B1(new_n1178), .B2(new_n698), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n645), .B1(new_n1147), .B2(KEYINPUT57), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1144), .A2(new_n1116), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT57), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1179), .B1(new_n1180), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1096), .A2(new_n644), .A3(new_n1100), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n1080), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1175), .A2(new_n1176), .A3(new_n1184), .A4(new_n1187), .ZN(G407));
  NAND2_X1  g0988(.A1(new_n624), .A2(G213), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1184), .A2(new_n1187), .A3(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(G407), .A2(G213), .A3(new_n1191), .ZN(G409));
  NAND2_X1  g0992(.A1(G387), .A2(new_n1044), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(G393), .B(new_n768), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n949), .A2(new_n974), .A3(G390), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1194), .ZN(new_n1197));
  AOI21_X1  g0997(.A(G390), .B1(new_n949), .B2(new_n974), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n974), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1199), .B(new_n1044), .C1(new_n931), .C2(new_n948), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1197), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1196), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1088), .A2(KEYINPUT60), .A3(new_n1090), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n644), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1095), .A2(KEYINPUT60), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1204), .B1(new_n1205), .B2(new_n1151), .ZN(new_n1206));
  OR3_X1    g1006(.A1(new_n1206), .A2(new_n804), .A3(new_n1170), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n804), .B1(new_n1206), .B2(new_n1170), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1190), .A2(G2897), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1209), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1142), .B1(new_n1181), .B2(new_n930), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1184), .A2(G378), .B1(new_n1187), .B2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1212), .B1(new_n1214), .B2(new_n1190), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1213), .A2(new_n1187), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1080), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1185), .A2(KEYINPUT120), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1092), .A2(new_n1081), .A3(new_n1096), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1217), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1216), .B1(G375), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT62), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1221), .A2(new_n1222), .A3(new_n1224), .A4(new_n1189), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT61), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1215), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  XOR2_X1   g1027(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n1228));
  NOR2_X1   g1028(.A1(new_n1214), .A2(new_n1190), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1228), .B1(new_n1229), .B2(new_n1224), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1202), .B1(new_n1227), .B2(new_n1230), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n1196), .A2(new_n1201), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1229), .A2(KEYINPUT63), .A3(new_n1224), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT63), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1221), .A2(new_n1189), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1234), .B1(new_n1235), .B2(new_n1223), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT61), .B1(new_n1235), .B2(new_n1212), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1232), .A2(new_n1233), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1231), .A2(new_n1238), .ZN(G405));
  NOR2_X1   g1039(.A1(G375), .A2(new_n1220), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1186), .B1(new_n1241), .B2(new_n1142), .ZN(new_n1242));
  OAI21_X1  g1042(.A(KEYINPUT126), .B1(new_n1240), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(G375), .A2(new_n1187), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1184), .A2(G378), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT126), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1243), .A2(new_n1223), .A3(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1223), .B1(new_n1243), .B2(new_n1247), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1202), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1247), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1246), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1224), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1243), .A2(new_n1223), .A3(new_n1247), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1253), .A2(new_n1232), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1250), .A2(new_n1255), .ZN(G402));
endmodule


