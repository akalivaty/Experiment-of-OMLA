

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581;

  NOR2_X1 U321 ( .A1(n578), .A2(n486), .ZN(n457) );
  OR2_X1 U322 ( .A1(n479), .A2(n533), .ZN(n480) );
  XNOR2_X1 U323 ( .A(G50GAT), .B(G29GAT), .ZN(n438) );
  XNOR2_X1 U324 ( .A(n289), .B(KEYINPUT55), .ZN(n479) );
  NOR2_X1 U325 ( .A1(n565), .A2(n478), .ZN(n289) );
  XNOR2_X1 U326 ( .A(n290), .B(n314), .ZN(n322) );
  XNOR2_X1 U327 ( .A(n313), .B(KEYINPUT9), .ZN(n290) );
  XNOR2_X1 U328 ( .A(n457), .B(KEYINPUT45), .ZN(n458) );
  AND2_X1 U329 ( .A1(n459), .A2(n291), .ZN(n460) );
  XNOR2_X1 U330 ( .A(n391), .B(KEYINPUT25), .ZN(n392) );
  XNOR2_X1 U331 ( .A(n423), .B(n294), .ZN(n431) );
  XNOR2_X1 U332 ( .A(n330), .B(n329), .ZN(n554) );
  XNOR2_X1 U333 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U334 ( .A(KEYINPUT79), .B(n554), .Z(n560) );
  XOR2_X1 U335 ( .A(n478), .B(KEYINPUT28), .Z(n528) );
  XOR2_X1 U336 ( .A(KEYINPUT92), .B(n402), .Z(n521) );
  NOR2_X1 U337 ( .A1(n571), .A2(n567), .ZN(n291) );
  XOR2_X1 U338 ( .A(KEYINPUT104), .B(KEYINPUT36), .Z(n292) );
  XOR2_X1 U339 ( .A(G134GAT), .B(G162GAT), .Z(n293) );
  XOR2_X1 U340 ( .A(n422), .B(n421), .Z(n294) );
  NOR2_X1 U341 ( .A1(n461), .A2(n507), .ZN(n463) );
  INV_X1 U342 ( .A(KEYINPUT98), .ZN(n391) );
  XNOR2_X1 U343 ( .A(n393), .B(n392), .ZN(n398) );
  NOR2_X1 U344 ( .A1(n554), .A2(n466), .ZN(n467) );
  INV_X1 U345 ( .A(KEYINPUT99), .ZN(n400) );
  XNOR2_X1 U346 ( .A(n377), .B(n312), .ZN(n313) );
  XNOR2_X1 U347 ( .A(n357), .B(n293), .ZN(n358) );
  XNOR2_X1 U348 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U349 ( .A(G43GAT), .B(G134GAT), .Z(n377) );
  XNOR2_X1 U350 ( .A(n560), .B(n292), .ZN(n578) );
  XNOR2_X1 U351 ( .A(n431), .B(n430), .ZN(n571) );
  INV_X1 U352 ( .A(G43GAT), .ZN(n454) );
  AND2_X1 U353 ( .A1(n560), .A2(n559), .ZN(n564) );
  XNOR2_X1 U354 ( .A(n451), .B(G50GAT), .ZN(n452) );
  XNOR2_X1 U355 ( .A(n454), .B(KEYINPUT40), .ZN(n455) );
  XNOR2_X1 U356 ( .A(n485), .B(n484), .ZN(G1349GAT) );
  XNOR2_X1 U357 ( .A(n453), .B(n452), .ZN(G1331GAT) );
  XOR2_X1 U358 ( .A(G148GAT), .B(KEYINPUT89), .Z(n296) );
  NAND2_X1 U359 ( .A1(G228GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U360 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U361 ( .A(n297), .B(KEYINPUT23), .Z(n305) );
  XOR2_X1 U362 ( .A(KEYINPUT3), .B(KEYINPUT88), .Z(n299) );
  XNOR2_X1 U363 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n298) );
  XNOR2_X1 U364 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U365 ( .A(G141GAT), .B(n300), .ZN(n362) );
  XOR2_X1 U366 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n302) );
  XNOR2_X1 U367 ( .A(G218GAT), .B(G106GAT), .ZN(n301) );
  XNOR2_X1 U368 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U369 ( .A(n362), .B(n303), .Z(n304) );
  XNOR2_X1 U370 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U371 ( .A(G22GAT), .B(G78GAT), .Z(n337) );
  XOR2_X1 U372 ( .A(n306), .B(n337), .Z(n310) );
  XOR2_X1 U373 ( .A(G50GAT), .B(G162GAT), .Z(n311) );
  XOR2_X1 U374 ( .A(G204GAT), .B(G211GAT), .Z(n308) );
  XNOR2_X1 U375 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n307) );
  XNOR2_X1 U376 ( .A(n308), .B(n307), .ZN(n381) );
  XNOR2_X1 U377 ( .A(n311), .B(n381), .ZN(n309) );
  XNOR2_X1 U378 ( .A(n310), .B(n309), .ZN(n478) );
  XOR2_X1 U379 ( .A(G29GAT), .B(G85GAT), .Z(n354) );
  XNOR2_X1 U380 ( .A(n311), .B(n354), .ZN(n314) );
  AND2_X1 U381 ( .A1(G232GAT), .A2(G233GAT), .ZN(n312) );
  XOR2_X1 U382 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n316) );
  XNOR2_X1 U383 ( .A(KEYINPUT10), .B(KEYINPUT74), .ZN(n315) );
  XNOR2_X1 U384 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U385 ( .A(KEYINPUT66), .B(KEYINPUT77), .Z(n318) );
  XNOR2_X1 U386 ( .A(KEYINPUT11), .B(KEYINPUT78), .ZN(n317) );
  XNOR2_X1 U387 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U388 ( .A(n320), .B(n319), .Z(n321) );
  XNOR2_X1 U389 ( .A(n322), .B(n321), .ZN(n330) );
  XNOR2_X1 U390 ( .A(G99GAT), .B(G106GAT), .ZN(n323) );
  XNOR2_X1 U391 ( .A(n323), .B(KEYINPUT73), .ZN(n427) );
  XOR2_X1 U392 ( .A(n427), .B(KEYINPUT67), .Z(n328) );
  XNOR2_X1 U393 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n324) );
  XNOR2_X1 U394 ( .A(n324), .B(KEYINPUT69), .ZN(n445) );
  XOR2_X1 U395 ( .A(G92GAT), .B(G218GAT), .Z(n326) );
  XNOR2_X1 U396 ( .A(G36GAT), .B(G190GAT), .ZN(n325) );
  XNOR2_X1 U397 ( .A(n326), .B(n325), .ZN(n380) );
  XNOR2_X1 U398 ( .A(n445), .B(n380), .ZN(n327) );
  XOR2_X1 U399 ( .A(KEYINPUT13), .B(KEYINPUT71), .Z(n416) );
  XOR2_X1 U400 ( .A(G8GAT), .B(G64GAT), .Z(n385) );
  XOR2_X1 U401 ( .A(n416), .B(n385), .Z(n332) );
  XNOR2_X1 U402 ( .A(G155GAT), .B(G211GAT), .ZN(n331) );
  XNOR2_X1 U403 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U404 ( .A(KEYINPUT15), .B(KEYINPUT80), .Z(n334) );
  NAND2_X1 U405 ( .A1(G231GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U406 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U407 ( .A(n336), .B(n335), .Z(n339) );
  XOR2_X1 U408 ( .A(G15GAT), .B(G1GAT), .Z(n441) );
  XNOR2_X1 U409 ( .A(n441), .B(n337), .ZN(n338) );
  XNOR2_X1 U410 ( .A(n339), .B(n338), .ZN(n347) );
  XOR2_X1 U411 ( .A(G57GAT), .B(G71GAT), .Z(n341) );
  XNOR2_X1 U412 ( .A(G183GAT), .B(G127GAT), .ZN(n340) );
  XNOR2_X1 U413 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U414 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n343) );
  XNOR2_X1 U415 ( .A(KEYINPUT81), .B(KEYINPUT82), .ZN(n342) );
  XNOR2_X1 U416 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U417 ( .A(n345), .B(n344), .Z(n346) );
  XOR2_X1 U418 ( .A(n347), .B(n346), .Z(n574) );
  XOR2_X1 U419 ( .A(KEYINPUT90), .B(KEYINPUT4), .Z(n349) );
  XNOR2_X1 U420 ( .A(KEYINPUT5), .B(KEYINPUT91), .ZN(n348) );
  XNOR2_X1 U421 ( .A(n349), .B(n348), .ZN(n361) );
  XOR2_X1 U422 ( .A(G120GAT), .B(G127GAT), .Z(n351) );
  XNOR2_X1 U423 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n350) );
  XNOR2_X1 U424 ( .A(n351), .B(n350), .ZN(n376) );
  XOR2_X1 U425 ( .A(n376), .B(G1GAT), .Z(n353) );
  NAND2_X1 U426 ( .A1(G225GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U427 ( .A(n353), .B(n352), .ZN(n359) );
  XOR2_X1 U428 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n356) );
  XOR2_X1 U429 ( .A(G148GAT), .B(G57GAT), .Z(n415) );
  XNOR2_X1 U430 ( .A(n354), .B(n415), .ZN(n355) );
  XNOR2_X1 U431 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U432 ( .A(n361), .B(n360), .ZN(n363) );
  XOR2_X1 U433 ( .A(n363), .B(n362), .Z(n402) );
  XOR2_X1 U434 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n365) );
  NAND2_X1 U435 ( .A1(G227GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U436 ( .A(n365), .B(n364), .ZN(n369) );
  XOR2_X1 U437 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n367) );
  XNOR2_X1 U438 ( .A(G99GAT), .B(G190GAT), .ZN(n366) );
  XNOR2_X1 U439 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U440 ( .A(n369), .B(n368), .Z(n374) );
  XOR2_X1 U441 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n371) );
  XNOR2_X1 U442 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n370) );
  XNOR2_X1 U443 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U444 ( .A(G169GAT), .B(n372), .Z(n389) );
  XNOR2_X1 U445 ( .A(G15GAT), .B(n389), .ZN(n373) );
  XNOR2_X1 U446 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U447 ( .A(G176GAT), .B(G71GAT), .Z(n422) );
  XOR2_X1 U448 ( .A(n375), .B(n422), .Z(n379) );
  XNOR2_X1 U449 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U450 ( .A(n379), .B(n378), .ZN(n533) );
  XOR2_X1 U451 ( .A(KEYINPUT93), .B(n380), .Z(n383) );
  XNOR2_X1 U452 ( .A(G176GAT), .B(n381), .ZN(n382) );
  XNOR2_X1 U453 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U454 ( .A(n385), .B(n384), .Z(n387) );
  NAND2_X1 U455 ( .A1(G226GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U456 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X2 U457 ( .A(n389), .B(n388), .Z(n523) );
  NOR2_X1 U458 ( .A1(n533), .A2(n523), .ZN(n390) );
  NOR2_X1 U459 ( .A1(n478), .A2(n390), .ZN(n393) );
  XOR2_X1 U460 ( .A(KEYINPUT26), .B(KEYINPUT97), .Z(n395) );
  NAND2_X1 U461 ( .A1(n478), .A2(n533), .ZN(n394) );
  XNOR2_X1 U462 ( .A(n395), .B(n394), .ZN(n566) );
  XOR2_X1 U463 ( .A(KEYINPUT27), .B(KEYINPUT94), .Z(n396) );
  XOR2_X1 U464 ( .A(n523), .B(n396), .Z(n403) );
  NOR2_X1 U465 ( .A1(n566), .A2(n403), .ZN(n397) );
  NOR2_X1 U466 ( .A1(n398), .A2(n397), .ZN(n399) );
  NOR2_X1 U467 ( .A1(n402), .A2(n399), .ZN(n401) );
  XNOR2_X1 U468 ( .A(n401), .B(n400), .ZN(n409) );
  INV_X1 U469 ( .A(n528), .ZN(n536) );
  NOR2_X1 U470 ( .A1(n521), .A2(n403), .ZN(n404) );
  XOR2_X1 U471 ( .A(KEYINPUT95), .B(n404), .Z(n532) );
  XOR2_X1 U472 ( .A(n533), .B(KEYINPUT87), .Z(n405) );
  NAND2_X1 U473 ( .A1(n532), .A2(n405), .ZN(n406) );
  NOR2_X1 U474 ( .A1(n536), .A2(n406), .ZN(n407) );
  XNOR2_X1 U475 ( .A(KEYINPUT96), .B(n407), .ZN(n408) );
  NOR2_X1 U476 ( .A1(n409), .A2(n408), .ZN(n489) );
  NOR2_X1 U477 ( .A1(n574), .A2(n489), .ZN(n410) );
  XNOR2_X1 U478 ( .A(n410), .B(KEYINPUT105), .ZN(n411) );
  NOR2_X1 U479 ( .A1(n578), .A2(n411), .ZN(n414) );
  XNOR2_X1 U480 ( .A(KEYINPUT37), .B(KEYINPUT106), .ZN(n412) );
  XNOR2_X1 U481 ( .A(n412), .B(KEYINPUT107), .ZN(n413) );
  XNOR2_X1 U482 ( .A(n414), .B(n413), .ZN(n519) );
  XOR2_X1 U483 ( .A(n416), .B(n415), .Z(n418) );
  NAND2_X1 U484 ( .A1(G230GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U485 ( .A(n418), .B(n417), .ZN(n423) );
  XOR2_X1 U486 ( .A(G92GAT), .B(G85GAT), .Z(n420) );
  XNOR2_X1 U487 ( .A(G204GAT), .B(G78GAT), .ZN(n419) );
  XNOR2_X1 U488 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U489 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n429) );
  XOR2_X1 U490 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n425) );
  XNOR2_X1 U491 ( .A(G120GAT), .B(G64GAT), .ZN(n424) );
  XNOR2_X1 U492 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U493 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U494 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U495 ( .A(G22GAT), .B(G197GAT), .Z(n433) );
  XNOR2_X1 U496 ( .A(G169GAT), .B(G141GAT), .ZN(n432) );
  XNOR2_X1 U497 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U498 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n435) );
  XNOR2_X1 U499 ( .A(G113GAT), .B(G8GAT), .ZN(n434) );
  XNOR2_X1 U500 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U501 ( .A(n437), .B(n436), .ZN(n449) );
  XOR2_X1 U502 ( .A(G43GAT), .B(G36GAT), .Z(n439) );
  XNOR2_X1 U503 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U504 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U505 ( .A1(G229GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U506 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U507 ( .A(n444), .B(KEYINPUT29), .Z(n447) );
  XNOR2_X1 U508 ( .A(n445), .B(KEYINPUT70), .ZN(n446) );
  XNOR2_X1 U509 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U510 ( .A(n449), .B(n448), .Z(n461) );
  NOR2_X1 U511 ( .A1(n571), .A2(n461), .ZN(n492) );
  NAND2_X1 U512 ( .A1(n519), .A2(n492), .ZN(n450) );
  XNOR2_X1 U513 ( .A(n450), .B(KEYINPUT38), .ZN(n505) );
  NOR2_X1 U514 ( .A1(n528), .A2(n505), .ZN(n453) );
  XNOR2_X1 U515 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n451) );
  NOR2_X1 U516 ( .A1(n533), .A2(n505), .ZN(n456) );
  XNOR2_X1 U517 ( .A(n456), .B(n455), .ZN(G1330GAT) );
  INV_X1 U518 ( .A(n574), .ZN(n486) );
  XNOR2_X1 U519 ( .A(n458), .B(KEYINPUT116), .ZN(n459) );
  INV_X1 U520 ( .A(n461), .ZN(n567) );
  XNOR2_X1 U521 ( .A(n460), .B(KEYINPUT117), .ZN(n469) );
  XOR2_X1 U522 ( .A(n571), .B(KEYINPUT41), .Z(n550) );
  INV_X1 U523 ( .A(n550), .ZN(n507) );
  XNOR2_X1 U524 ( .A(KEYINPUT46), .B(KEYINPUT114), .ZN(n462) );
  XNOR2_X1 U525 ( .A(n463), .B(n462), .ZN(n464) );
  NOR2_X1 U526 ( .A1(n574), .A2(n464), .ZN(n465) );
  XNOR2_X1 U527 ( .A(n465), .B(KEYINPUT115), .ZN(n466) );
  XNOR2_X1 U528 ( .A(KEYINPUT47), .B(n467), .ZN(n468) );
  NAND2_X1 U529 ( .A1(n469), .A2(n468), .ZN(n471) );
  XNOR2_X1 U530 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n470) );
  XNOR2_X1 U531 ( .A(n471), .B(n470), .ZN(n531) );
  INV_X1 U532 ( .A(n523), .ZN(n472) );
  NAND2_X1 U533 ( .A1(n531), .A2(n472), .ZN(n474) );
  XOR2_X1 U534 ( .A(KEYINPUT122), .B(KEYINPUT54), .Z(n473) );
  XNOR2_X1 U535 ( .A(n474), .B(n473), .ZN(n475) );
  NAND2_X1 U536 ( .A1(n475), .A2(n521), .ZN(n477) );
  INV_X1 U537 ( .A(KEYINPUT65), .ZN(n476) );
  XNOR2_X1 U538 ( .A(n477), .B(n476), .ZN(n565) );
  XNOR2_X2 U539 ( .A(n480), .B(KEYINPUT123), .ZN(n559) );
  NAND2_X1 U540 ( .A1(n559), .A2(n567), .ZN(n482) );
  XNOR2_X1 U541 ( .A(G169GAT), .B(KEYINPUT124), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n482), .B(n481), .ZN(G1348GAT) );
  NAND2_X1 U543 ( .A1(n559), .A2(n550), .ZN(n485) );
  XOR2_X1 U544 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n483) );
  XNOR2_X1 U545 ( .A(n483), .B(G176GAT), .ZN(n484) );
  XOR2_X1 U546 ( .A(KEYINPUT16), .B(KEYINPUT83), .Z(n488) );
  OR2_X1 U547 ( .A1(n486), .A2(n560), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(n490) );
  NOR2_X1 U549 ( .A1(n490), .A2(n489), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n491), .B(KEYINPUT100), .ZN(n508) );
  NAND2_X1 U551 ( .A1(n492), .A2(n508), .ZN(n500) );
  NOR2_X1 U552 ( .A1(n521), .A2(n500), .ZN(n494) );
  XNOR2_X1 U553 ( .A(KEYINPUT34), .B(KEYINPUT101), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U555 ( .A(G1GAT), .B(n495), .ZN(G1324GAT) );
  NOR2_X1 U556 ( .A1(n523), .A2(n500), .ZN(n496) );
  XOR2_X1 U557 ( .A(G8GAT), .B(n496), .Z(G1325GAT) );
  NOR2_X1 U558 ( .A1(n533), .A2(n500), .ZN(n498) );
  XNOR2_X1 U559 ( .A(KEYINPUT35), .B(KEYINPUT102), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U561 ( .A(G15GAT), .B(n499), .ZN(G1326GAT) );
  NOR2_X1 U562 ( .A1(n528), .A2(n500), .ZN(n502) );
  XNOR2_X1 U563 ( .A(G22GAT), .B(KEYINPUT103), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(G1327GAT) );
  NOR2_X1 U565 ( .A1(n505), .A2(n521), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n503), .B(KEYINPUT39), .ZN(n504) );
  XNOR2_X1 U567 ( .A(G29GAT), .B(n504), .ZN(G1328GAT) );
  NOR2_X1 U568 ( .A1(n523), .A2(n505), .ZN(n506) );
  XOR2_X1 U569 ( .A(G36GAT), .B(n506), .Z(G1329GAT) );
  NOR2_X1 U570 ( .A1(n567), .A2(n507), .ZN(n520) );
  NAND2_X1 U571 ( .A1(n520), .A2(n508), .ZN(n516) );
  NOR2_X1 U572 ( .A1(n521), .A2(n516), .ZN(n510) );
  XNOR2_X1 U573 ( .A(KEYINPUT42), .B(KEYINPUT110), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U575 ( .A(G57GAT), .B(n511), .Z(G1332GAT) );
  NOR2_X1 U576 ( .A1(n523), .A2(n516), .ZN(n513) );
  XNOR2_X1 U577 ( .A(G64GAT), .B(KEYINPUT111), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(G1333GAT) );
  NOR2_X1 U579 ( .A1(n533), .A2(n516), .ZN(n514) );
  XOR2_X1 U580 ( .A(KEYINPUT112), .B(n514), .Z(n515) );
  XNOR2_X1 U581 ( .A(G71GAT), .B(n515), .ZN(G1334GAT) );
  NOR2_X1 U582 ( .A1(n528), .A2(n516), .ZN(n518) );
  XNOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n518), .B(n517), .ZN(G1335GAT) );
  NAND2_X1 U585 ( .A1(n520), .A2(n519), .ZN(n527) );
  NOR2_X1 U586 ( .A1(n521), .A2(n527), .ZN(n522) );
  XOR2_X1 U587 ( .A(G85GAT), .B(n522), .Z(G1336GAT) );
  NOR2_X1 U588 ( .A1(n523), .A2(n527), .ZN(n524) );
  XOR2_X1 U589 ( .A(G92GAT), .B(n524), .Z(G1337GAT) );
  NOR2_X1 U590 ( .A1(n533), .A2(n527), .ZN(n526) );
  XNOR2_X1 U591 ( .A(G99GAT), .B(KEYINPUT113), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(G1338GAT) );
  NOR2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U594 ( .A(KEYINPUT44), .B(n529), .Z(n530) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n530), .ZN(G1339GAT) );
  NAND2_X1 U596 ( .A1(n532), .A2(n531), .ZN(n545) );
  NOR2_X1 U597 ( .A1(n533), .A2(n545), .ZN(n534) );
  XOR2_X1 U598 ( .A(KEYINPUT118), .B(n534), .Z(n535) );
  NOR2_X1 U599 ( .A1(n536), .A2(n535), .ZN(n542) );
  NAND2_X1 U600 ( .A1(n542), .A2(n567), .ZN(n537) );
  XNOR2_X1 U601 ( .A(n537), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U602 ( .A(G120GAT), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U603 ( .A1(n542), .A2(n550), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  NAND2_X1 U605 ( .A1(n542), .A2(n574), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n540), .B(KEYINPUT50), .ZN(n541) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n541), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U609 ( .A1(n542), .A2(n560), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NOR2_X1 U611 ( .A1(n566), .A2(n545), .ZN(n555) );
  NAND2_X1 U612 ( .A1(n567), .A2(n555), .ZN(n546) );
  XNOR2_X1 U613 ( .A(G141GAT), .B(n546), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n548) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U617 ( .A(KEYINPUT119), .B(n549), .Z(n552) );
  NAND2_X1 U618 ( .A1(n555), .A2(n550), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(G1345GAT) );
  NAND2_X1 U620 ( .A1(n555), .A2(n574), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n553), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U622 ( .A(G162GAT), .B(KEYINPUT121), .Z(n557) );
  NAND2_X1 U623 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1347GAT) );
  NAND2_X1 U625 ( .A1(n559), .A2(n574), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n558), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U627 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(KEYINPUT125), .ZN(n562) );
  XNOR2_X1 U629 ( .A(KEYINPUT126), .B(n562), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1351GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n569) );
  NOR2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n576) );
  NAND2_X1 U633 ( .A1(n576), .A2(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(G204GAT), .B(KEYINPUT61), .Z(n573) );
  NAND2_X1 U637 ( .A1(n576), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  NAND2_X1 U639 ( .A1(n576), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U641 ( .A(n576), .ZN(n577) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

