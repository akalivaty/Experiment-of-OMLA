//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n562, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XNOR2_X1  g016(.A(KEYINPUT64), .B(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  XOR2_X1   g032(.A(G325), .B(KEYINPUT67), .Z(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT68), .Z(new_n460));
  NAND2_X1  g035(.A1(new_n456), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n466), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n469), .B1(new_n466), .B2(new_n468), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  XOR2_X1   g048(.A(new_n473), .B(KEYINPUT70), .Z(new_n474));
  AOI21_X1  g049(.A(new_n464), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G101), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n466), .A2(new_n468), .ZN(new_n477));
  INV_X1    g052(.A(G137), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(new_n464), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n475), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT71), .ZN(G160));
  NOR2_X1   g058(.A1(new_n477), .A2(new_n464), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n466), .A2(new_n468), .A3(new_n464), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  NOR2_X1   g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(new_n464), .B2(G112), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n485), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  NOR2_X1   g067(.A1(new_n467), .A2(G2104), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT69), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n466), .A2(new_n468), .A3(new_n469), .ZN(new_n496));
  AOI21_X1  g071(.A(G2105), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(KEYINPUT4), .B1(new_n497), .B2(G138), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(new_n464), .B2(G114), .ZN(new_n499));
  NOR2_X1   g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT72), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n500), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n502), .A2(new_n504), .A3(new_n505), .A4(G2104), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT4), .A2(G138), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n466), .A2(new_n468), .A3(new_n508), .A4(new_n464), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n466), .A2(new_n468), .A3(G126), .A4(G2105), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n507), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n498), .A2(new_n511), .ZN(G164));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n515), .B(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT74), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n518), .B1(new_n519), .B2(G651), .ZN(new_n520));
  NOR3_X1   g095(.A1(new_n514), .A2(KEYINPUT74), .A3(KEYINPUT6), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n517), .A2(G543), .A3(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT5), .ZN(new_n524));
  OAI21_X1  g099(.A(KEYINPUT75), .B1(new_n524), .B2(G543), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT75), .ZN(new_n526));
  INV_X1    g101(.A(G543), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n526), .A2(new_n527), .A3(KEYINPUT5), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n525), .A2(new_n528), .B1(new_n524), .B2(G543), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n517), .A2(new_n529), .A3(new_n522), .ZN(new_n530));
  INV_X1    g105(.A(G88), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n513), .A2(new_n523), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n529), .A2(G62), .ZN(new_n533));
  NAND2_X1  g108(.A1(G75), .A2(G543), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT76), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n514), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n532), .A2(new_n536), .ZN(G303));
  INV_X1    g112(.A(G303), .ZN(G166));
  NAND3_X1  g113(.A1(new_n517), .A2(G89), .A3(new_n522), .ZN(new_n539));
  INV_X1    g114(.A(G63), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n540), .B2(new_n514), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(new_n529), .ZN(new_n542));
  INV_X1    g117(.A(new_n523), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G51), .ZN(new_n544));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT7), .ZN(new_n546));
  AND3_X1   g121(.A1(new_n542), .A2(new_n544), .A3(new_n546), .ZN(G168));
  INV_X1    g122(.A(G52), .ZN(new_n548));
  INV_X1    g123(.A(G90), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n548), .A2(new_n523), .B1(new_n530), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n529), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n514), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n550), .A2(new_n552), .ZN(G171));
  NAND2_X1  g128(.A1(new_n543), .A2(G43), .ZN(new_n554));
  INV_X1    g129(.A(new_n530), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G81), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n529), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(new_n514), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n554), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(G188));
  XNOR2_X1  g141(.A(KEYINPUT78), .B(G65), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n529), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n514), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(G53), .ZN(new_n571));
  OR3_X1    g146(.A1(new_n523), .A2(KEYINPUT9), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT9), .B1(new_n523), .B2(new_n571), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n570), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT77), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n530), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n517), .A2(KEYINPUT77), .A3(new_n529), .A4(new_n522), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G91), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n574), .A2(new_n579), .ZN(G299));
  INV_X1    g155(.A(G171), .ZN(G301));
  NOR2_X1   g156(.A1(G168), .A2(KEYINPUT79), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n542), .A2(new_n544), .A3(new_n546), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G286));
  NAND2_X1  g162(.A1(new_n578), .A2(G87), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n529), .B2(G74), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT80), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n543), .A2(G49), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(G288));
  INV_X1    g167(.A(G48), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n529), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n593), .A2(new_n523), .B1(new_n594), .B2(new_n514), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(new_n578), .B2(G86), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT81), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G305));
  AOI22_X1  g174(.A1(new_n529), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(new_n514), .ZN(new_n601));
  XOR2_X1   g176(.A(new_n601), .B(KEYINPUT82), .Z(new_n602));
  NAND2_X1  g177(.A1(new_n555), .A2(G85), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n543), .A2(G47), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n543), .A2(G54), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n529), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n608), .A2(new_n514), .ZN(new_n609));
  AOI21_X1  g184(.A(KEYINPUT10), .B1(new_n578), .B2(G92), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  AOI211_X1 g187(.A(new_n611), .B(new_n612), .C1(new_n576), .C2(new_n577), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n607), .B(new_n609), .C1(new_n610), .C2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n606), .B1(new_n615), .B2(G868), .ZN(G321));
  XOR2_X1   g191(.A(G321), .B(KEYINPUT83), .Z(G284));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(G299), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(new_n586), .B2(new_n618), .ZN(G297));
  OAI21_X1  g195(.A(new_n619), .B1(new_n586), .B2(new_n618), .ZN(G280));
  XNOR2_X1  g196(.A(KEYINPUT84), .B(G559), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n615), .B1(G860), .B2(new_n623), .ZN(G148));
  NAND2_X1  g199(.A1(new_n559), .A2(new_n618), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n614), .A2(new_n622), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(new_n618), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n495), .A2(new_n496), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n629), .A2(G2104), .A3(new_n464), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2100), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n464), .A2(G111), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n465), .B1(new_n634), .B2(KEYINPUT85), .ZN(new_n635));
  OAI221_X1 g210(.A(new_n635), .B1(KEYINPUT85), .B2(new_n634), .C1(G99), .C2(G2105), .ZN(new_n636));
  AOI22_X1  g211(.A1(G123), .A2(new_n484), .B1(new_n487), .B2(G135), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(G2096), .Z(new_n639));
  NAND2_X1  g214(.A1(new_n633), .A2(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XOR2_X1   g217(.A(KEYINPUT15), .B(G2435), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT14), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n645), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT87), .B(KEYINPUT88), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G1341), .B(G1348), .Z(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n651), .B(new_n654), .Z(new_n655));
  AND2_X1   g230(.A1(new_n655), .A2(G14), .ZN(G401));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2072), .B(G2078), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT17), .ZN(new_n659));
  XOR2_X1   g234(.A(G2067), .B(G2678), .Z(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n657), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n661), .B2(new_n658), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT89), .Z(new_n664));
  NAND3_X1  g239(.A1(new_n661), .A2(new_n657), .A3(new_n658), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT18), .Z(new_n666));
  INV_X1    g241(.A(new_n659), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n667), .A2(new_n657), .A3(new_n660), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n664), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2096), .B(G2100), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G227));
  XNOR2_X1  g247(.A(G1961), .B(G1966), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT91), .ZN(new_n674));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT92), .Z(new_n681));
  AND2_X1   g256(.A1(new_n674), .A2(new_n675), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(new_n679), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT20), .ZN(new_n684));
  OR3_X1    g259(.A1(new_n682), .A2(new_n676), .A3(new_n679), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n681), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1981), .B(G1986), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT95), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G1991), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n689), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G229));
  INV_X1    g271(.A(G29), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G33), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n487), .A2(G139), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT25), .Z(new_n701));
  AOI22_X1  g276(.A1(new_n629), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n699), .B(new_n701), .C1(new_n702), .C2(new_n464), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n703), .A2(KEYINPUT99), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(KEYINPUT99), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n698), .B1(new_n706), .B2(new_n697), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G2072), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n560), .A2(G16), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G16), .B2(G19), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT98), .B(G1341), .Z(new_n711));
  NAND2_X1  g286(.A1(new_n697), .A2(G26), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n484), .A2(G128), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n487), .A2(G140), .ZN(new_n714));
  OR2_X1    g289(.A1(G104), .A2(G2105), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n715), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n713), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n712), .B1(new_n718), .B2(new_n697), .ZN(new_n719));
  MUX2_X1   g294(.A(new_n712), .B(new_n719), .S(KEYINPUT28), .Z(new_n720));
  AOI22_X1  g295(.A1(new_n710), .A2(new_n711), .B1(new_n720), .B2(G2067), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n697), .A2(G27), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G164), .B2(new_n697), .ZN(new_n723));
  INV_X1    g298(.A(G2078), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n721), .B(new_n725), .C1(G2067), .C2(new_n720), .ZN(new_n726));
  INV_X1    g301(.A(G1961), .ZN(new_n727));
  NAND2_X1  g302(.A1(G171), .A2(G16), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G5), .B2(G16), .ZN(new_n729));
  OAI22_X1  g304(.A1(new_n710), .A2(new_n711), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  AOI22_X1  g305(.A1(G129), .A2(new_n484), .B1(new_n487), .B2(G141), .ZN(new_n731));
  NAND3_X1  g306(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT26), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT101), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G29), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G29), .B2(G32), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT27), .B(G1996), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n697), .A2(G35), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G162), .B2(new_n697), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT29), .B(G2090), .Z(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n739), .A2(new_n740), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT30), .B(G28), .Z(new_n747));
  MUX2_X1   g322(.A(new_n747), .B(new_n638), .S(G29), .Z(new_n748));
  NAND4_X1  g323(.A1(new_n741), .A2(new_n745), .A3(new_n746), .A4(new_n748), .ZN(new_n749));
  NOR3_X1   g324(.A1(new_n726), .A2(new_n730), .A3(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G16), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G4), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n615), .B2(new_n751), .ZN(new_n753));
  INV_X1    g328(.A(G1348), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT31), .B(G11), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT100), .ZN(new_n757));
  NOR2_X1   g332(.A1(KEYINPUT24), .A2(G34), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(KEYINPUT24), .A2(G34), .ZN(new_n760));
  AOI21_X1  g335(.A(G29), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  AOI22_X1  g336(.A1(G160), .A2(G29), .B1(new_n757), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n757), .B2(new_n761), .ZN(new_n763));
  INV_X1    g338(.A(G2084), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n763), .A2(new_n764), .B1(new_n727), .B2(new_n729), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n750), .A2(new_n755), .A3(new_n756), .A4(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(G16), .A2(G21), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G168), .B2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1966), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n763), .A2(new_n764), .ZN(new_n771));
  INV_X1    g346(.A(G1956), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n751), .A2(G20), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT23), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n574), .A2(new_n579), .ZN(new_n776));
  OAI21_X1  g351(.A(KEYINPUT23), .B1(new_n776), .B2(new_n751), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n775), .B1(new_n777), .B2(new_n773), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n771), .B1(new_n772), .B2(new_n778), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n770), .B(new_n779), .C1(new_n772), .C2(new_n778), .ZN(new_n780));
  NOR2_X1   g355(.A1(G6), .A2(G16), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n598), .B2(G16), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT32), .ZN(new_n783));
  INV_X1    g358(.A(G1981), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n751), .A2(G22), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G166), .B2(new_n751), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(G1971), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n751), .A2(G23), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G288), .B2(G16), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT33), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n791), .A2(G1976), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n791), .A2(G1976), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n787), .A2(G1971), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n785), .A2(new_n788), .A3(new_n795), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n796), .A2(KEYINPUT34), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n484), .A2(G119), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n487), .A2(G131), .ZN(new_n799));
  OR2_X1    g374(.A1(G95), .A2(G2105), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n800), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n798), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  MUX2_X1   g377(.A(G25), .B(new_n802), .S(G29), .Z(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT35), .B(G1991), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT96), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n803), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n751), .A2(G24), .ZN(new_n807));
  INV_X1    g382(.A(G290), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(new_n751), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT97), .B(G1986), .Z(new_n810));
  XOR2_X1   g385(.A(new_n809), .B(new_n810), .Z(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n796), .B2(KEYINPUT34), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n797), .A2(new_n806), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(KEYINPUT36), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT36), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n797), .A2(new_n812), .A3(new_n815), .A4(new_n806), .ZN(new_n816));
  AOI211_X1 g391(.A(new_n708), .B(new_n780), .C1(new_n814), .C2(new_n816), .ZN(G311));
  AOI21_X1  g392(.A(new_n780), .B1(new_n814), .B2(new_n816), .ZN(new_n818));
  INV_X1    g393(.A(new_n708), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(G150));
  AOI22_X1  g395(.A1(G55), .A2(new_n543), .B1(new_n555), .B2(G93), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n529), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n514), .B2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT105), .B(G860), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT37), .Z(new_n826));
  NAND2_X1  g401(.A1(new_n615), .A2(G559), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT103), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n823), .B(new_n559), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n828), .B(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT39), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT104), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n824), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n836), .B2(new_n835), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n833), .A2(new_n834), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n826), .B1(new_n838), .B2(new_n839), .ZN(G145));
  INV_X1    g415(.A(new_n737), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n704), .A2(new_n705), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n842), .A2(KEYINPUT107), .A3(new_n717), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n717), .B1(new_n842), .B2(KEYINPUT107), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT106), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n498), .A2(new_n846), .A3(new_n511), .ZN(new_n847));
  AND3_X1   g422(.A1(new_n507), .A2(new_n509), .A3(new_n510), .ZN(new_n848));
  OAI211_X1 g423(.A(G138), .B(new_n464), .C1(new_n470), .C2(new_n471), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT4), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(KEYINPUT106), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n847), .A2(new_n852), .ZN(new_n853));
  NOR3_X1   g428(.A1(new_n844), .A2(new_n845), .A3(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n853), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT107), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n718), .B1(new_n706), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n855), .B1(new_n857), .B2(new_n843), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n841), .B1(new_n854), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n853), .B1(new_n844), .B2(new_n845), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n857), .A2(new_n843), .A3(new_n855), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n860), .A2(new_n861), .A3(new_n737), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n484), .A2(G130), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n487), .A2(G142), .ZN(new_n865));
  NOR2_X1   g440(.A1(G106), .A2(G2105), .ZN(new_n866));
  OAI21_X1  g441(.A(G2104), .B1(new_n464), .B2(G118), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n864), .B(new_n865), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n631), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n802), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n863), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT108), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n859), .A2(new_n870), .A3(new_n862), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(G160), .B(new_n638), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(G162), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n874), .A2(new_n873), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n875), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(G37), .ZN(new_n880));
  INV_X1    g455(.A(new_n877), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n872), .A2(new_n874), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g459(.A(KEYINPUT109), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(new_n614), .B2(new_n776), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n614), .A2(new_n776), .A3(new_n885), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n615), .A2(G299), .ZN(new_n889));
  AND4_X1   g464(.A1(KEYINPUT41), .A2(new_n887), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(KEYINPUT110), .A3(new_n888), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT110), .ZN(new_n892));
  INV_X1    g467(.A(new_n888), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n892), .B1(new_n893), .B2(new_n886), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(new_n894), .A3(new_n889), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n890), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n829), .B(new_n626), .Z(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n893), .A2(new_n886), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n889), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  OR3_X1    g477(.A1(new_n899), .A2(KEYINPUT42), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(G288), .B(G303), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n904), .A2(new_n598), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n598), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n906), .A2(new_n808), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n808), .B1(new_n906), .B2(new_n907), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT42), .B1(new_n899), .B2(new_n902), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n903), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n910), .B1(new_n903), .B2(new_n911), .ZN(new_n913));
  OAI21_X1  g488(.A(G868), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n823), .A2(new_n618), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(G295));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n915), .ZN(G331));
  OAI21_X1  g492(.A(G171), .B1(new_n582), .B2(new_n585), .ZN(new_n918));
  NAND2_X1  g493(.A1(G168), .A2(G301), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n829), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n830), .A2(new_n918), .A3(new_n919), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n897), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n923), .A2(new_n901), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(G37), .B1(new_n927), .B2(new_n910), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n925), .B1(new_n897), .B2(new_n923), .ZN(new_n929));
  INV_X1    g504(.A(new_n910), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT43), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n880), .B1(new_n929), .B2(new_n930), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n921), .A2(new_n922), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n900), .B(new_n889), .C1(new_n935), .C2(new_n896), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n923), .A2(new_n895), .A3(KEYINPUT41), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n930), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n933), .A2(new_n934), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT44), .B1(new_n932), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n931), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT43), .B1(new_n941), .B2(new_n933), .ZN(new_n942));
  INV_X1    g517(.A(new_n938), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n928), .A2(new_n943), .A3(new_n934), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n940), .B1(new_n946), .B2(KEYINPUT44), .ZN(G397));
  NOR2_X1   g522(.A1(G290), .A2(G1986), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n737), .B(G1996), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n802), .A2(new_n804), .ZN(new_n950));
  OR2_X1    g525(.A1(new_n802), .A2(new_n804), .ZN(new_n951));
  INV_X1    g526(.A(G2067), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n717), .B(new_n952), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n949), .A2(new_n950), .A3(new_n951), .A4(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n948), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G1986), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n955), .B1(new_n956), .B2(new_n808), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n958));
  XOR2_X1   g533(.A(KEYINPUT111), .B(G1384), .Z(new_n959));
  OAI21_X1  g534(.A(new_n958), .B1(new_n853), .B2(new_n959), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n472), .A2(new_n474), .ZN(new_n961));
  OAI211_X1 g536(.A(G40), .B(new_n480), .C1(new_n961), .C2(new_n464), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n957), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G40), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n475), .A2(new_n965), .A3(new_n481), .ZN(new_n966));
  AOI21_X1  g541(.A(G1384), .B1(new_n848), .B2(new_n851), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n966), .B1(new_n967), .B2(KEYINPUT45), .ZN(new_n968));
  INV_X1    g543(.A(new_n959), .ZN(new_n969));
  OAI211_X1 g544(.A(KEYINPUT45), .B(new_n969), .C1(new_n847), .C2(new_n852), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT112), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n846), .B1(new_n498), .B2(new_n511), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n848), .A2(new_n851), .A3(KEYINPUT106), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n959), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT112), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n974), .A2(new_n975), .A3(KEYINPUT45), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n968), .B1(new_n971), .B2(new_n976), .ZN(new_n977));
  OR2_X1    g552(.A1(new_n977), .A2(G1971), .ZN(new_n978));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n498), .B2(new_n511), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n966), .B1(new_n980), .B2(KEYINPUT50), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT113), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n983), .B1(new_n980), .B2(KEYINPUT50), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT50), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n967), .A2(KEYINPUT113), .A3(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n982), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT114), .B1(new_n987), .B2(G2090), .ZN(new_n988));
  OR3_X1    g563(.A1(new_n987), .A2(KEYINPUT114), .A3(G2090), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n978), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n990), .A2(G8), .ZN(new_n991));
  NAND2_X1  g566(.A1(G303), .A2(G8), .ZN(new_n992));
  NAND2_X1  g567(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n993));
  OR2_X1    g568(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n995), .B1(new_n992), .B2(new_n993), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n991), .A2(new_n997), .ZN(new_n998));
  OR2_X1    g573(.A1(new_n998), .A2(KEYINPUT116), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(KEYINPUT116), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n966), .A2(new_n967), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G8), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT49), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n555), .A2(G86), .ZN(new_n1007));
  OAI21_X1  g582(.A(G1981), .B1(new_n1007), .B2(new_n595), .ZN(new_n1008));
  OR2_X1    g583(.A1(new_n1008), .A2(KEYINPUT117), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n596), .A2(new_n784), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1008), .A2(KEYINPUT117), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n1012), .A2(KEYINPUT118), .A3(new_n1006), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT118), .B1(new_n1012), .B2(new_n1006), .ZN(new_n1014));
  OAI221_X1 g589(.A(new_n1005), .B1(new_n1006), .B2(new_n1012), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G1976), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1005), .B1(new_n1016), .B2(G288), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT52), .ZN(new_n1018));
  INV_X1    g593(.A(G288), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1019), .A2(G1976), .ZN(new_n1020));
  OR3_X1    g595(.A1(new_n1017), .A2(KEYINPUT52), .A3(new_n1020), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n1015), .A2(new_n1018), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n978), .ZN(new_n1023));
  INV_X1    g598(.A(G2090), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n967), .A2(new_n985), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n981), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1023), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n996), .B1(new_n1027), .B2(new_n1004), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1001), .A2(new_n1022), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT119), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1026), .A2(G1956), .ZN(new_n1031));
  XNOR2_X1  g606(.A(KEYINPUT56), .B(G2072), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1031), .B1(new_n977), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT57), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G299), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n574), .A2(KEYINPUT57), .A3(new_n579), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1030), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n968), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n970), .A2(KEYINPUT112), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n975), .B1(new_n974), .B2(KEYINPUT45), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1039), .B(new_n1032), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1031), .ZN(new_n1043));
  AND4_X1   g618(.A1(new_n1030), .A2(new_n1042), .A3(new_n1037), .A4(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1038), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1037), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT121), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT121), .ZN(new_n1049));
  AOI211_X1 g624(.A(new_n1049), .B(new_n1037), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n1002), .A2(KEYINPUT120), .A3(G2067), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n987), .B2(new_n754), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT120), .B1(new_n1002), .B2(G2067), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n614), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1045), .B1(new_n1051), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1053), .A2(KEYINPUT60), .A3(new_n1054), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT60), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1057), .B1(new_n1058), .B2(new_n614), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1053), .A2(KEYINPUT60), .A3(new_n615), .A4(new_n1054), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT61), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1062), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT59), .ZN(new_n1065));
  INV_X1    g640(.A(G1996), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n977), .A2(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT58), .B(G1341), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1003), .A2(new_n1068), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1065), .B(new_n560), .C1(new_n1067), .C2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1069), .B1(new_n977), .B2(new_n1066), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT59), .B1(new_n1071), .B2(new_n559), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1061), .A2(new_n1064), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT122), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1076));
  AOI211_X1 g651(.A(KEYINPUT122), .B(new_n1037), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT61), .B1(new_n1078), .B2(new_n1045), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1056), .B1(new_n1074), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT123), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n977), .A2(new_n724), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1084), .A2(new_n1085), .B1(new_n727), .B2(new_n987), .ZN(new_n1086));
  XOR2_X1   g661(.A(new_n480), .B(KEYINPUT125), .Z(new_n1087));
  NOR2_X1   g662(.A1(new_n475), .A2(new_n965), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI211_X1 g664(.A(KEYINPUT53), .B(new_n724), .C1(new_n1089), .C2(KEYINPUT126), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(KEYINPUT126), .B2(new_n1089), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1091), .B(new_n960), .C1(new_n1041), .C2(new_n1040), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1086), .A2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1093), .A2(G171), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n980), .A2(new_n958), .ZN(new_n1095));
  OR4_X1    g670(.A1(new_n1085), .A2(new_n968), .A3(new_n1095), .A4(G2078), .ZN(new_n1096));
  AOI21_X1  g671(.A(G301), .B1(new_n1086), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1083), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n982), .B(new_n764), .C1(new_n984), .C2(new_n986), .ZN(new_n1099));
  INV_X1    g674(.A(G1966), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1100), .B1(new_n968), .B2(new_n1095), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1099), .A2(KEYINPUT124), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT124), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1103));
  NOR3_X1   g678(.A1(new_n1102), .A2(new_n1103), .A3(new_n583), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT51), .B1(new_n1104), .B2(new_n1004), .ZN(new_n1105));
  OAI211_X1 g680(.A(G8), .B(new_n583), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1107));
  OAI21_X1  g682(.A(G8), .B1(new_n1107), .B2(new_n583), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1105), .B(new_n1106), .C1(KEYINPUT51), .C2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1093), .A2(G171), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1086), .A2(G301), .A3(new_n1096), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(KEYINPUT54), .A3(new_n1111), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1098), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1113));
  OAI211_X1 g688(.A(KEYINPUT123), .B(new_n1056), .C1(new_n1074), .C2(new_n1079), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1082), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1109), .A2(KEYINPUT62), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1109), .A2(KEYINPUT62), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(new_n1097), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1029), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1015), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1010), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n1005), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1022), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1107), .A2(G8), .A3(new_n586), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n991), .B2(new_n997), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT63), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1124), .A2(KEYINPUT63), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n999), .A2(new_n1000), .B1(new_n1028), .B2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1122), .B(new_n1127), .C1(new_n1129), .C2(new_n1123), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n964), .B1(new_n1119), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n948), .A2(new_n963), .ZN(new_n1132));
  XOR2_X1   g707(.A(new_n1132), .B(KEYINPUT48), .Z(new_n1133));
  AOI21_X1  g708(.A(new_n1133), .B1(new_n963), .B2(new_n954), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n960), .A2(G1996), .A3(new_n962), .ZN(new_n1135));
  OR2_X1    g710(.A1(new_n1135), .A2(KEYINPUT46), .ZN(new_n1136));
  INV_X1    g711(.A(new_n953), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n963), .B1(new_n841), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1135), .A2(KEYINPUT46), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1136), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  XOR2_X1   g715(.A(new_n1140), .B(KEYINPUT47), .Z(new_n1141));
  NAND2_X1  g716(.A1(new_n949), .A2(new_n953), .ZN(new_n1142));
  OAI22_X1  g717(.A1(new_n1142), .A2(new_n951), .B1(G2067), .B2(new_n717), .ZN(new_n1143));
  AOI211_X1 g718(.A(new_n1134), .B(new_n1141), .C1(new_n963), .C2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1131), .A2(new_n1144), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g720(.A(new_n934), .B1(new_n928), .B2(new_n931), .ZN(new_n1147));
  NOR3_X1   g721(.A1(new_n933), .A2(KEYINPUT43), .A3(new_n938), .ZN(new_n1148));
  OAI21_X1  g722(.A(new_n695), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g723(.A1(G401), .A2(new_n462), .ZN(new_n1150));
  NAND3_X1  g724(.A1(new_n883), .A2(new_n671), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g725(.A(KEYINPUT127), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  AND3_X1   g726(.A1(new_n883), .A2(new_n671), .A3(new_n1150), .ZN(new_n1153));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n1154));
  NAND4_X1  g728(.A1(new_n1153), .A2(new_n1154), .A3(new_n695), .A4(new_n945), .ZN(new_n1155));
  NAND2_X1  g729(.A1(new_n1152), .A2(new_n1155), .ZN(G308));
  NAND3_X1  g730(.A1(new_n1153), .A2(new_n695), .A3(new_n945), .ZN(G225));
endmodule


