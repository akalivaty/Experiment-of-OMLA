

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584;

  NOR2_X2 U323 ( .A1(n386), .A2(n385), .ZN(n387) );
  XOR2_X1 U324 ( .A(n301), .B(n300), .Z(n291) );
  XOR2_X1 U325 ( .A(n432), .B(n391), .Z(n292) );
  XNOR2_X1 U326 ( .A(n333), .B(KEYINPUT72), .ZN(n334) );
  XNOR2_X1 U327 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U328 ( .A(n337), .B(n303), .Z(n482) );
  XNOR2_X1 U329 ( .A(n388), .B(KEYINPUT48), .ZN(n544) );
  XNOR2_X1 U330 ( .A(n448), .B(n447), .ZN(n560) );
  XNOR2_X1 U331 ( .A(n449), .B(G183GAT), .ZN(n450) );
  XNOR2_X1 U332 ( .A(n451), .B(n450), .ZN(G1350GAT) );
  XOR2_X1 U333 ( .A(G64GAT), .B(KEYINPUT13), .Z(n294) );
  XNOR2_X1 U334 ( .A(G71GAT), .B(G78GAT), .ZN(n293) );
  XNOR2_X1 U335 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U336 ( .A(G57GAT), .B(n295), .Z(n337) );
  XOR2_X1 U337 ( .A(G22GAT), .B(G155GAT), .Z(n432) );
  XNOR2_X1 U338 ( .A(G8GAT), .B(G183GAT), .ZN(n296) );
  XNOR2_X1 U339 ( .A(n296), .B(G211GAT), .ZN(n391) );
  NAND2_X1 U340 ( .A1(G231GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U341 ( .A(n292), .B(n297), .ZN(n301) );
  XOR2_X1 U342 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n299) );
  XNOR2_X1 U343 ( .A(KEYINPUT15), .B(KEYINPUT80), .ZN(n298) );
  XNOR2_X1 U344 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U345 ( .A(G1GAT), .B(KEYINPUT70), .Z(n348) );
  XOR2_X1 U346 ( .A(G15GAT), .B(G127GAT), .Z(n306) );
  XNOR2_X1 U347 ( .A(n348), .B(n306), .ZN(n302) );
  XNOR2_X1 U348 ( .A(n291), .B(n302), .ZN(n303) );
  XOR2_X1 U349 ( .A(KEYINPUT111), .B(n482), .Z(n533) );
  XOR2_X1 U350 ( .A(G183GAT), .B(KEYINPUT20), .Z(n305) );
  XNOR2_X1 U351 ( .A(KEYINPUT83), .B(KEYINPUT65), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n318) );
  XOR2_X1 U353 ( .A(KEYINPUT84), .B(G99GAT), .Z(n308) );
  XOR2_X1 U354 ( .A(G176GAT), .B(G120GAT), .Z(n332) );
  XNOR2_X1 U355 ( .A(n332), .B(n306), .ZN(n307) );
  XNOR2_X1 U356 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U357 ( .A(n309), .B(G190GAT), .Z(n316) );
  XOR2_X1 U358 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n311) );
  XNOR2_X1 U359 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n310) );
  XNOR2_X1 U360 ( .A(n311), .B(n310), .ZN(n399) );
  XOR2_X1 U361 ( .A(n399), .B(G71GAT), .Z(n313) );
  NAND2_X1 U362 ( .A1(G227GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U364 ( .A(G43GAT), .B(n314), .ZN(n315) );
  XNOR2_X1 U365 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U366 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U367 ( .A(KEYINPUT81), .B(G134GAT), .Z(n320) );
  XNOR2_X1 U368 ( .A(KEYINPUT82), .B(KEYINPUT0), .ZN(n319) );
  XNOR2_X1 U369 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U370 ( .A(G113GAT), .B(n321), .ZN(n408) );
  XOR2_X1 U371 ( .A(n322), .B(n408), .Z(n520) );
  INV_X1 U372 ( .A(n520), .ZN(n526) );
  INV_X1 U373 ( .A(KEYINPUT41), .ZN(n338) );
  XOR2_X1 U374 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n324) );
  NAND2_X1 U375 ( .A1(G230GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U377 ( .A(n325), .B(KEYINPUT31), .Z(n331) );
  XOR2_X1 U378 ( .A(G148GAT), .B(G204GAT), .Z(n327) );
  XNOR2_X1 U379 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n437) );
  XOR2_X1 U381 ( .A(G92GAT), .B(KEYINPUT74), .Z(n329) );
  XNOR2_X1 U382 ( .A(G99GAT), .B(G85GAT), .ZN(n328) );
  XNOR2_X1 U383 ( .A(n329), .B(n328), .ZN(n367) );
  XNOR2_X1 U384 ( .A(n437), .B(n367), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n331), .B(n330), .ZN(n335) );
  XNOR2_X1 U386 ( .A(n332), .B(KEYINPUT32), .ZN(n333) );
  XNOR2_X1 U387 ( .A(n337), .B(n336), .ZN(n574) );
  XNOR2_X1 U388 ( .A(n338), .B(n574), .ZN(n498) );
  XOR2_X1 U389 ( .A(G15GAT), .B(G113GAT), .Z(n340) );
  XNOR2_X1 U390 ( .A(G169GAT), .B(G197GAT), .ZN(n339) );
  XNOR2_X1 U391 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U392 ( .A(KEYINPUT69), .B(KEYINPUT29), .Z(n342) );
  XNOR2_X1 U393 ( .A(G8GAT), .B(KEYINPUT30), .ZN(n341) );
  XNOR2_X1 U394 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U395 ( .A(n344), .B(n343), .ZN(n357) );
  XOR2_X1 U396 ( .A(G141GAT), .B(G22GAT), .Z(n346) );
  XNOR2_X1 U397 ( .A(G50GAT), .B(G36GAT), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U399 ( .A(n348), .B(n347), .Z(n350) );
  NAND2_X1 U400 ( .A1(G229GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U401 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U402 ( .A(n351), .B(KEYINPUT71), .Z(n355) );
  XOR2_X1 U403 ( .A(G29GAT), .B(G43GAT), .Z(n353) );
  XNOR2_X1 U404 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n352) );
  XNOR2_X1 U405 ( .A(n353), .B(n352), .ZN(n368) );
  XNOR2_X1 U406 ( .A(n368), .B(KEYINPUT68), .ZN(n354) );
  XNOR2_X1 U407 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U408 ( .A(n357), .B(n356), .Z(n570) );
  NOR2_X1 U409 ( .A1(n498), .A2(n570), .ZN(n358) );
  XNOR2_X1 U410 ( .A(n358), .B(KEYINPUT46), .ZN(n359) );
  NOR2_X1 U411 ( .A1(n359), .A2(n533), .ZN(n360) );
  XNOR2_X1 U412 ( .A(n360), .B(KEYINPUT112), .ZN(n378) );
  XOR2_X1 U413 ( .A(KEYINPUT67), .B(KEYINPUT77), .Z(n362) );
  XNOR2_X1 U414 ( .A(KEYINPUT9), .B(KEYINPUT10), .ZN(n361) );
  XNOR2_X1 U415 ( .A(n362), .B(n361), .ZN(n377) );
  XOR2_X1 U416 ( .A(KEYINPUT78), .B(KEYINPUT11), .Z(n364) );
  NAND2_X1 U417 ( .A1(G232GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U418 ( .A(n364), .B(n363), .ZN(n366) );
  XNOR2_X1 U419 ( .A(G36GAT), .B(G190GAT), .ZN(n365) );
  XNOR2_X1 U420 ( .A(n365), .B(KEYINPUT79), .ZN(n398) );
  XOR2_X1 U421 ( .A(n366), .B(n398), .Z(n370) );
  XNOR2_X1 U422 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U423 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U424 ( .A(n371), .B(G106GAT), .Z(n375) );
  XOR2_X1 U425 ( .A(G162GAT), .B(KEYINPUT76), .Z(n373) );
  XNOR2_X1 U426 ( .A(G50GAT), .B(G218GAT), .ZN(n372) );
  XNOR2_X1 U427 ( .A(n373), .B(n372), .ZN(n438) );
  XNOR2_X1 U428 ( .A(G134GAT), .B(n438), .ZN(n374) );
  XNOR2_X1 U429 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U430 ( .A(n377), .B(n376), .ZN(n538) );
  INV_X1 U431 ( .A(n538), .ZN(n555) );
  NAND2_X1 U432 ( .A1(n378), .A2(n555), .ZN(n379) );
  XNOR2_X1 U433 ( .A(n379), .B(KEYINPUT47), .ZN(n386) );
  XOR2_X1 U434 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n382) );
  XOR2_X1 U435 ( .A(KEYINPUT36), .B(KEYINPUT100), .Z(n380) );
  XOR2_X1 U436 ( .A(n538), .B(n380), .Z(n582) );
  NAND2_X1 U437 ( .A1(n482), .A2(n582), .ZN(n381) );
  XNOR2_X1 U438 ( .A(n382), .B(n381), .ZN(n383) );
  NAND2_X1 U439 ( .A1(n574), .A2(n383), .ZN(n384) );
  INV_X1 U440 ( .A(n570), .ZN(n558) );
  NOR2_X1 U441 ( .A1(n384), .A2(n558), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n387), .B(KEYINPUT64), .ZN(n388) );
  XOR2_X1 U443 ( .A(G92GAT), .B(G204GAT), .Z(n390) );
  XNOR2_X1 U444 ( .A(G176GAT), .B(G218GAT), .ZN(n389) );
  XNOR2_X1 U445 ( .A(n390), .B(n389), .ZN(n403) );
  XOR2_X1 U446 ( .A(G197GAT), .B(KEYINPUT21), .Z(n428) );
  XOR2_X1 U447 ( .A(n391), .B(n428), .Z(n393) );
  NAND2_X1 U448 ( .A1(G226GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U449 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U450 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n395) );
  XNOR2_X1 U451 ( .A(G64GAT), .B(KEYINPUT93), .ZN(n394) );
  XNOR2_X1 U452 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U453 ( .A(n397), .B(n396), .Z(n401) );
  XNOR2_X1 U454 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U456 ( .A(n403), .B(n402), .Z(n505) );
  INV_X1 U457 ( .A(n505), .ZN(n518) );
  NOR2_X1 U458 ( .A1(n544), .A2(n518), .ZN(n404) );
  XNOR2_X1 U459 ( .A(KEYINPUT54), .B(n404), .ZN(n566) );
  XOR2_X1 U460 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n406) );
  XNOR2_X1 U461 ( .A(KEYINPUT90), .B(KEYINPUT6), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U463 ( .A(n408), .B(n407), .Z(n422) );
  XOR2_X1 U464 ( .A(G85GAT), .B(G155GAT), .Z(n410) );
  XNOR2_X1 U465 ( .A(G120GAT), .B(G148GAT), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n414) );
  XOR2_X1 U467 ( .A(G57GAT), .B(KEYINPUT1), .Z(n412) );
  XNOR2_X1 U468 ( .A(G1GAT), .B(G127GAT), .ZN(n411) );
  XNOR2_X1 U469 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U470 ( .A(n414), .B(n413), .Z(n420) );
  XNOR2_X1 U471 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n415), .B(KEYINPUT2), .ZN(n431) );
  XOR2_X1 U473 ( .A(n431), .B(G162GAT), .Z(n417) );
  NAND2_X1 U474 ( .A1(G225GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U476 ( .A(G29GAT), .B(n418), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U478 ( .A(n422), .B(n421), .Z(n567) );
  XOR2_X1 U479 ( .A(KEYINPUT89), .B(KEYINPUT22), .Z(n424) );
  XNOR2_X1 U480 ( .A(KEYINPUT88), .B(KEYINPUT85), .ZN(n423) );
  XNOR2_X1 U481 ( .A(n424), .B(n423), .ZN(n442) );
  XOR2_X1 U482 ( .A(KEYINPUT24), .B(G78GAT), .Z(n426) );
  XNOR2_X1 U483 ( .A(G211GAT), .B(KEYINPUT87), .ZN(n425) );
  XNOR2_X1 U484 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U485 ( .A(n427), .B(KEYINPUT23), .Z(n430) );
  XNOR2_X1 U486 ( .A(n428), .B(KEYINPUT86), .ZN(n429) );
  XNOR2_X1 U487 ( .A(n430), .B(n429), .ZN(n436) );
  XOR2_X1 U488 ( .A(n432), .B(n431), .Z(n434) );
  NAND2_X1 U489 ( .A1(G228GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U490 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U491 ( .A(n436), .B(n435), .Z(n440) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U493 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U494 ( .A(n442), .B(n441), .ZN(n461) );
  AND2_X1 U495 ( .A1(n567), .A2(n461), .ZN(n443) );
  NAND2_X1 U496 ( .A1(n566), .A2(n443), .ZN(n445) );
  XOR2_X1 U497 ( .A(KEYINPUT55), .B(KEYINPUT121), .Z(n444) );
  XNOR2_X1 U498 ( .A(n445), .B(n444), .ZN(n446) );
  NAND2_X1 U499 ( .A1(n526), .A2(n446), .ZN(n448) );
  INV_X1 U500 ( .A(KEYINPUT122), .ZN(n447) );
  NAND2_X1 U501 ( .A1(n533), .A2(n560), .ZN(n451) );
  XOR2_X1 U502 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n449) );
  INV_X1 U503 ( .A(G190GAT), .ZN(n455) );
  NAND2_X1 U504 ( .A1(n560), .A2(n538), .ZN(n453) );
  XOR2_X1 U505 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n452) );
  XNOR2_X1 U506 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n455), .B(n454), .ZN(G1351GAT) );
  AND2_X1 U508 ( .A1(n558), .A2(n574), .ZN(n485) );
  INV_X1 U509 ( .A(n482), .ZN(n578) );
  NOR2_X1 U510 ( .A1(n538), .A2(n578), .ZN(n456) );
  XNOR2_X1 U511 ( .A(KEYINPUT16), .B(n456), .ZN(n468) );
  XNOR2_X1 U512 ( .A(KEYINPUT27), .B(n505), .ZN(n459) );
  INV_X1 U513 ( .A(n567), .ZN(n502) );
  NAND2_X1 U514 ( .A1(n459), .A2(n502), .ZN(n457) );
  XNOR2_X1 U515 ( .A(n457), .B(KEYINPUT94), .ZN(n543) );
  XNOR2_X1 U516 ( .A(KEYINPUT28), .B(n461), .ZN(n523) );
  INV_X1 U517 ( .A(n523), .ZN(n509) );
  NOR2_X1 U518 ( .A1(n543), .A2(n509), .ZN(n527) );
  NAND2_X1 U519 ( .A1(n520), .A2(n527), .ZN(n467) );
  NOR2_X1 U520 ( .A1(n461), .A2(n526), .ZN(n458) );
  XNOR2_X1 U521 ( .A(n458), .B(KEYINPUT26), .ZN(n568) );
  NAND2_X1 U522 ( .A1(n459), .A2(n568), .ZN(n464) );
  NAND2_X1 U523 ( .A1(n505), .A2(n526), .ZN(n460) );
  NAND2_X1 U524 ( .A1(n461), .A2(n460), .ZN(n462) );
  XOR2_X1 U525 ( .A(KEYINPUT25), .B(n462), .Z(n463) );
  NAND2_X1 U526 ( .A1(n464), .A2(n463), .ZN(n465) );
  NAND2_X1 U527 ( .A1(n465), .A2(n567), .ZN(n466) );
  NAND2_X1 U528 ( .A1(n467), .A2(n466), .ZN(n480) );
  NAND2_X1 U529 ( .A1(n468), .A2(n480), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n469), .B(KEYINPUT95), .ZN(n500) );
  NAND2_X1 U531 ( .A1(n485), .A2(n500), .ZN(n477) );
  NOR2_X1 U532 ( .A1(n567), .A2(n477), .ZN(n471) );
  XNOR2_X1 U533 ( .A(KEYINPUT96), .B(KEYINPUT34), .ZN(n470) );
  XNOR2_X1 U534 ( .A(n471), .B(n470), .ZN(n472) );
  XOR2_X1 U535 ( .A(G1GAT), .B(n472), .Z(G1324GAT) );
  NOR2_X1 U536 ( .A1(n518), .A2(n477), .ZN(n474) );
  XNOR2_X1 U537 ( .A(G8GAT), .B(KEYINPUT97), .ZN(n473) );
  XNOR2_X1 U538 ( .A(n474), .B(n473), .ZN(G1325GAT) );
  NOR2_X1 U539 ( .A1(n520), .A2(n477), .ZN(n476) );
  XNOR2_X1 U540 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n475) );
  XNOR2_X1 U541 ( .A(n476), .B(n475), .ZN(G1326GAT) );
  NOR2_X1 U542 ( .A1(n523), .A2(n477), .ZN(n478) );
  XOR2_X1 U543 ( .A(G22GAT), .B(n478), .Z(n479) );
  XNOR2_X1 U544 ( .A(KEYINPUT98), .B(n479), .ZN(G1327GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT99), .B(KEYINPUT39), .Z(n488) );
  NAND2_X1 U546 ( .A1(n582), .A2(n480), .ZN(n481) );
  NOR2_X1 U547 ( .A1(n482), .A2(n481), .ZN(n484) );
  XNOR2_X1 U548 ( .A(KEYINPUT101), .B(KEYINPUT37), .ZN(n483) );
  XNOR2_X1 U549 ( .A(n484), .B(n483), .ZN(n515) );
  NAND2_X1 U550 ( .A1(n485), .A2(n515), .ZN(n486) );
  XOR2_X1 U551 ( .A(KEYINPUT38), .B(n486), .Z(n494) );
  NAND2_X1 U552 ( .A1(n502), .A2(n494), .ZN(n487) );
  XNOR2_X1 U553 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U554 ( .A(G29GAT), .B(n489), .Z(G1328GAT) );
  NAND2_X1 U555 ( .A1(n494), .A2(n505), .ZN(n490) );
  XNOR2_X1 U556 ( .A(n490), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT40), .B(KEYINPUT102), .Z(n492) );
  NAND2_X1 U558 ( .A1(n494), .A2(n526), .ZN(n491) );
  XNOR2_X1 U559 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U560 ( .A(G43GAT), .B(n493), .Z(G1330GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n496) );
  NAND2_X1 U562 ( .A1(n494), .A2(n509), .ZN(n495) );
  XNOR2_X1 U563 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U564 ( .A(G50GAT), .B(n497), .ZN(G1331GAT) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n498), .B(KEYINPUT105), .ZN(n561) );
  NAND2_X1 U567 ( .A1(n561), .A2(n570), .ZN(n499) );
  XOR2_X1 U568 ( .A(KEYINPUT106), .B(n499), .Z(n514) );
  NAND2_X1 U569 ( .A1(n500), .A2(n514), .ZN(n501) );
  XNOR2_X1 U570 ( .A(KEYINPUT107), .B(n501), .ZN(n510) );
  NAND2_X1 U571 ( .A1(n502), .A2(n510), .ZN(n503) );
  XNOR2_X1 U572 ( .A(n504), .B(n503), .ZN(G1332GAT) );
  NAND2_X1 U573 ( .A1(n510), .A2(n505), .ZN(n506) );
  XNOR2_X1 U574 ( .A(n506), .B(KEYINPUT108), .ZN(n507) );
  XNOR2_X1 U575 ( .A(G64GAT), .B(n507), .ZN(G1333GAT) );
  NAND2_X1 U576 ( .A1(n526), .A2(n510), .ZN(n508) );
  XNOR2_X1 U577 ( .A(n508), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n512) );
  NAND2_X1 U579 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U580 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U581 ( .A(G78GAT), .B(n513), .Z(G1335GAT) );
  NAND2_X1 U582 ( .A1(n515), .A2(n514), .ZN(n522) );
  NOR2_X1 U583 ( .A1(n567), .A2(n522), .ZN(n516) );
  XOR2_X1 U584 ( .A(G85GAT), .B(n516), .Z(n517) );
  XNOR2_X1 U585 ( .A(KEYINPUT110), .B(n517), .ZN(G1336GAT) );
  NOR2_X1 U586 ( .A1(n518), .A2(n522), .ZN(n519) );
  XOR2_X1 U587 ( .A(G92GAT), .B(n519), .Z(G1337GAT) );
  NOR2_X1 U588 ( .A1(n520), .A2(n522), .ZN(n521) );
  XOR2_X1 U589 ( .A(G99GAT), .B(n521), .Z(G1338GAT) );
  NOR2_X1 U590 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U591 ( .A(KEYINPUT44), .B(n524), .Z(n525) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n525), .ZN(G1339GAT) );
  NAND2_X1 U593 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U594 ( .A1(n544), .A2(n528), .ZN(n539) );
  NAND2_X1 U595 ( .A1(n539), .A2(n558), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n529), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT49), .B(KEYINPUT113), .Z(n531) );
  NAND2_X1 U598 ( .A1(n539), .A2(n561), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U600 ( .A(G120GAT), .B(n532), .Z(G1341GAT) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(KEYINPUT114), .ZN(n537) );
  XOR2_X1 U602 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n535) );
  NAND2_X1 U603 ( .A1(n539), .A2(n533), .ZN(n534) );
  XNOR2_X1 U604 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n537), .B(n536), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U607 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U609 ( .A(G134GAT), .B(n542), .ZN(G1343GAT) );
  NOR2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U611 ( .A1(n545), .A2(n568), .ZN(n554) );
  NOR2_X1 U612 ( .A1(n570), .A2(n554), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n549) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n548) );
  XNOR2_X1 U617 ( .A(n549), .B(n548), .ZN(n551) );
  NOR2_X1 U618 ( .A1(n498), .A2(n554), .ZN(n550) );
  XOR2_X1 U619 ( .A(n551), .B(n550), .Z(G1345GAT) );
  NOR2_X1 U620 ( .A1(n578), .A2(n554), .ZN(n553) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n552) );
  XNOR2_X1 U622 ( .A(n553), .B(n552), .ZN(G1346GAT) );
  NOR2_X1 U623 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U624 ( .A(KEYINPUT120), .B(n556), .Z(n557) );
  XNOR2_X1 U625 ( .A(G162GAT), .B(n557), .ZN(G1347GAT) );
  NAND2_X1 U626 ( .A1(n558), .A2(n560), .ZN(n559) );
  XNOR2_X1 U627 ( .A(G169GAT), .B(n559), .ZN(G1348GAT) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n563) );
  XOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT57), .Z(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n565) );
  XOR2_X1 U631 ( .A(KEYINPUT123), .B(KEYINPUT56), .Z(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  AND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n569) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n580) );
  NOR2_X1 U635 ( .A1(n570), .A2(n580), .ZN(n572) );
  XNOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(n573), .ZN(G1352GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n580), .ZN(n576) );
  XNOR2_X1 U640 ( .A(KEYINPUT61), .B(KEYINPUT127), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U642 ( .A(G204GAT), .B(n577), .Z(G1353GAT) );
  NOR2_X1 U643 ( .A1(n578), .A2(n580), .ZN(n579) );
  XOR2_X1 U644 ( .A(G211GAT), .B(n579), .Z(G1354GAT) );
  INV_X1 U645 ( .A(n580), .ZN(n581) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n583), .B(KEYINPUT62), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

