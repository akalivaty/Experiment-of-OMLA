//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AND2_X1   g0006(.A1(G116), .A2(G270), .ZN(new_n207));
  INV_X1    g0007(.A(G77), .ZN(new_n208));
  INV_X1    g0008(.A(G244), .ZN(new_n209));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  OAI22_X1  g0011(.A1(new_n208), .A2(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI211_X1 g0012(.A(new_n207), .B(new_n212), .C1(G87), .C2(G250), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G58), .A2(G232), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G107), .A2(G264), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G50), .A2(G226), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n206), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT1), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n206), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT0), .ZN(new_n225));
  OR2_X1    g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n224), .A2(new_n225), .ZN(new_n227));
  NAND3_X1  g0027(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n228));
  INV_X1    g0028(.A(new_n201), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n226), .B(new_n227), .C1(new_n228), .C2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT64), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n222), .A2(new_n232), .ZN(G361));
  XOR2_X1   g0033(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G226), .B(G232), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  INV_X1    g0043(.A(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(KEYINPUT66), .B(G107), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XOR2_X1   g0048(.A(G50), .B(G58), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G20), .ZN(new_n252));
  OAI21_X1  g0052(.A(KEYINPUT23), .B1(new_n252), .B2(G107), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT23), .ZN(new_n254));
  INV_X1    g0054(.A(G107), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(new_n255), .A3(G20), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n252), .A2(G33), .A3(G116), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n253), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT78), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n253), .A2(new_n256), .A3(new_n257), .A4(KEYINPUT78), .ZN(new_n261));
  AND2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n252), .B(G87), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT22), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OR2_X1    g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n270), .A2(KEYINPUT22), .A3(new_n252), .A4(G87), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(KEYINPUT79), .B1(new_n262), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n260), .A2(new_n261), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT79), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n274), .A2(new_n275), .A3(new_n267), .A4(new_n271), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n273), .A2(KEYINPUT24), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G1), .A2(G13), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT24), .ZN(new_n281));
  OAI211_X1 g0081(.A(KEYINPUT79), .B(new_n281), .C1(new_n262), .C2(new_n272), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n277), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT25), .ZN(new_n284));
  INV_X1    g0084(.A(G13), .ZN(new_n285));
  NOR3_X1   g0085(.A1(new_n285), .A2(new_n252), .A3(G1), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n284), .B1(new_n287), .B2(G107), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(KEYINPUT25), .A3(new_n255), .ZN(new_n289));
  INV_X1    g0089(.A(G33), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(G1), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n286), .A2(new_n280), .A3(new_n291), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n288), .A2(new_n289), .B1(new_n292), .B2(G107), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n283), .A2(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(G257), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT80), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n270), .A2(KEYINPUT80), .A3(G257), .A4(G1698), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G294), .ZN(new_n299));
  INV_X1    g0099(.A(G1698), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n270), .A2(G250), .A3(new_n300), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n297), .A2(new_n298), .A3(new_n299), .A4(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G33), .A2(G41), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n303), .A2(G1), .A3(G13), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G1), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT5), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n307), .B(G45), .C1(new_n308), .C2(G41), .ZN(new_n309));
  INV_X1    g0109(.A(G41), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n310), .A2(KEYINPUT5), .ZN(new_n311));
  OAI211_X1 g0111(.A(G264), .B(new_n304), .C1(new_n309), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n307), .A2(G45), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n308), .A2(G41), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n310), .A2(KEYINPUT5), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n314), .A2(new_n315), .A3(new_n316), .A4(G274), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n306), .A2(new_n312), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G169), .ZN(new_n319));
  INV_X1    g0119(.A(new_n312), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(new_n302), .B2(new_n305), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n321), .A2(G179), .A3(new_n317), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n294), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT81), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT81), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n294), .A2(new_n326), .A3(new_n323), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  OAI211_X1 g0128(.A(G226), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT75), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT75), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n270), .A2(new_n331), .A3(G226), .A4(G1698), .ZN(new_n332));
  NAND2_X1  g0132(.A1(G33), .A2(G87), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n270), .A2(G223), .A3(new_n300), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n330), .A2(new_n332), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n305), .ZN(new_n336));
  INV_X1    g0136(.A(G190), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n307), .B1(G41), .B2(G45), .ZN(new_n338));
  INV_X1    g0138(.A(G274), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n304), .A2(new_n338), .ZN(new_n342));
  INV_X1    g0142(.A(G232), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n336), .A2(new_n337), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT76), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n336), .A2(new_n345), .ZN(new_n348));
  INV_X1    g0148(.A(G200), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT76), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n336), .A2(new_n351), .A3(new_n337), .A4(new_n345), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n347), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT16), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT7), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(new_n270), .B2(G20), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n263), .A2(new_n264), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n357), .A2(KEYINPUT7), .A3(new_n252), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n218), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G58), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n360), .A2(new_n218), .ZN(new_n361));
  OAI21_X1  g0161(.A(G20), .B1(new_n361), .B2(new_n201), .ZN(new_n362));
  NOR2_X1   g0162(.A1(G20), .A2(G33), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G159), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n354), .B1(new_n359), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(KEYINPUT7), .B1(new_n357), .B2(new_n252), .ZN(new_n367));
  NOR4_X1   g0167(.A1(new_n263), .A2(new_n264), .A3(new_n355), .A4(G20), .ZN(new_n368));
  OAI21_X1  g0168(.A(G68), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n365), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n369), .A2(KEYINPUT16), .A3(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n366), .A2(new_n280), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n280), .B1(new_n307), .B2(G20), .ZN(new_n373));
  XNOR2_X1  g0173(.A(KEYINPUT8), .B(G58), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(new_n286), .ZN(new_n377));
  AND3_X1   g0177(.A1(new_n372), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  AND3_X1   g0178(.A1(new_n353), .A2(new_n378), .A3(KEYINPUT17), .ZN(new_n379));
  AOI21_X1  g0179(.A(KEYINPUT17), .B1(new_n353), .B2(new_n378), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n372), .A2(new_n376), .A3(new_n377), .ZN(new_n382));
  AOI21_X1  g0182(.A(G169), .B1(new_n336), .B2(new_n345), .ZN(new_n383));
  AOI211_X1 g0183(.A(G179), .B(new_n344), .C1(new_n335), .C2(new_n305), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT18), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n382), .A2(new_n385), .A3(KEYINPUT18), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n381), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n373), .A2(G77), .ZN(new_n391));
  XOR2_X1   g0191(.A(new_n391), .B(KEYINPUT73), .Z(new_n392));
  AOI22_X1  g0192(.A1(new_n375), .A2(new_n363), .B1(G20), .B2(G77), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n252), .A2(G33), .ZN(new_n394));
  XOR2_X1   g0194(.A(KEYINPUT15), .B(G87), .Z(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n393), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n397), .A2(new_n280), .B1(new_n208), .B2(new_n286), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n392), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n270), .A2(G238), .A3(G1698), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n270), .A2(G232), .A3(new_n300), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n400), .B(new_n401), .C1(new_n255), .C2(new_n270), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n305), .ZN(new_n403));
  INV_X1    g0203(.A(G179), .ZN(new_n404));
  INV_X1    g0204(.A(new_n342), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(G244), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n403), .A2(new_n404), .A3(new_n341), .A4(new_n406), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n403), .A2(new_n341), .A3(new_n406), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n399), .B(new_n407), .C1(new_n408), .C2(G169), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(G190), .ZN(new_n410));
  XOR2_X1   g0210(.A(KEYINPUT74), .B(G200), .Z(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n410), .B1(new_n412), .B2(new_n408), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n409), .B1(new_n413), .B2(new_n399), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n390), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n373), .A2(G50), .ZN(new_n416));
  INV_X1    g0216(.A(G150), .ZN(new_n417));
  INV_X1    g0217(.A(new_n363), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n374), .A2(new_n394), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(G20), .B2(new_n203), .ZN(new_n420));
  INV_X1    g0220(.A(new_n280), .ZN(new_n421));
  OAI221_X1 g0221(.A(new_n416), .B1(G50), .B2(new_n287), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n422), .B(KEYINPUT9), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  OR2_X1    g0224(.A1(G222), .A2(G1698), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT68), .B(G223), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n425), .B1(new_n426), .B2(new_n300), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n270), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n357), .A2(new_n208), .ZN(new_n429));
  AND3_X1   g0229(.A1(new_n428), .A2(KEYINPUT69), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT69), .B1(new_n428), .B2(new_n429), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n305), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT67), .ZN(new_n433));
  OR2_X1    g0233(.A1(new_n433), .A2(G226), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(G226), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n405), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n432), .A2(new_n341), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT70), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n432), .A2(KEYINPUT70), .A3(new_n341), .A4(new_n436), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n424), .B1(new_n441), .B2(G190), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n439), .A2(new_n411), .A3(new_n440), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT10), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT10), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n442), .A2(new_n446), .A3(new_n443), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G169), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n439), .A2(new_n449), .A3(new_n440), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n422), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT71), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n450), .A2(KEYINPUT71), .A3(new_n422), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT72), .ZN(new_n456));
  INV_X1    g0256(.A(new_n441), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n456), .B1(new_n457), .B2(G179), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n441), .A2(KEYINPUT72), .A3(new_n404), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n270), .A2(G226), .A3(new_n300), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n270), .A2(G232), .A3(G1698), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n462), .B(new_n463), .C1(new_n290), .C2(new_n210), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n340), .B1(new_n464), .B2(new_n305), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT13), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n405), .A2(G238), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n466), .B1(new_n465), .B2(new_n467), .ZN(new_n470));
  OAI21_X1  g0270(.A(G169), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT14), .ZN(new_n472));
  INV_X1    g0272(.A(new_n470), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(G179), .A3(new_n468), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT14), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n475), .B(G169), .C1(new_n469), .C2(new_n470), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n472), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  OAI22_X1  g0277(.A1(new_n418), .A2(new_n202), .B1(new_n252), .B2(G68), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n394), .A2(new_n208), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n280), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  XOR2_X1   g0280(.A(new_n480), .B(KEYINPUT11), .Z(new_n481));
  AND2_X1   g0281(.A1(new_n373), .A2(G68), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n286), .A2(new_n218), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT12), .ZN(new_n484));
  XNOR2_X1  g0284(.A(new_n483), .B(new_n484), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n481), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n477), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(G200), .B1(new_n469), .B2(new_n470), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n473), .A2(G190), .A3(new_n468), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n489), .A2(new_n490), .A3(new_n486), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  AND4_X1   g0292(.A1(new_n415), .A2(new_n448), .A3(new_n461), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G283), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n494), .B(new_n252), .C1(G33), .C2(new_n210), .ZN(new_n495));
  OR2_X1    g0295(.A1(KEYINPUT77), .A2(KEYINPUT20), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n244), .A2(G20), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n495), .A2(new_n280), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(KEYINPUT77), .A2(KEYINPUT20), .ZN(new_n499));
  XNOR2_X1  g0299(.A(new_n498), .B(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n292), .A2(G116), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n500), .B(new_n501), .C1(G116), .C2(new_n287), .ZN(new_n502));
  OAI211_X1 g0302(.A(G257), .B(new_n300), .C1(new_n263), .C2(new_n264), .ZN(new_n503));
  OAI211_X1 g0303(.A(G264), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n504));
  INV_X1    g0304(.A(G303), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n503), .B(new_n504), .C1(new_n505), .C2(new_n270), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n305), .ZN(new_n507));
  OAI211_X1 g0307(.A(G270), .B(new_n304), .C1(new_n309), .C2(new_n311), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n508), .A2(new_n317), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n502), .A2(G169), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT21), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n502), .A2(G179), .A3(new_n507), .A4(new_n509), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n502), .A2(KEYINPUT21), .A3(G169), .A4(new_n510), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n502), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n510), .A2(new_n337), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n518), .B1(G200), .B2(new_n510), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n516), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n219), .A2(new_n300), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n209), .A2(G1698), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n521), .B(new_n522), .C1(new_n263), .C2(new_n264), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G116), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n304), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n313), .A2(new_n339), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n304), .A2(G250), .A3(new_n313), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NOR3_X1   g0328(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n529), .A2(new_n412), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n287), .A2(new_n395), .ZN(new_n531));
  NAND3_X1  g0331(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n252), .ZN(new_n533));
  NOR2_X1   g0333(.A1(G97), .A2(G107), .ZN(new_n534));
  INV_X1    g0334(.A(G87), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n252), .A2(G33), .A3(G97), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT19), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n533), .A2(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n270), .A2(new_n252), .A3(G68), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n531), .B1(new_n541), .B2(new_n280), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n292), .A2(G87), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n530), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n529), .A2(G190), .ZN(new_n546));
  INV_X1    g0346(.A(new_n526), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n523), .A2(new_n524), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n547), .B(new_n527), .C1(new_n548), .C2(new_n304), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n292), .A2(new_n395), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n449), .A2(new_n549), .B1(new_n542), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n529), .A2(new_n404), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n545), .A2(new_n546), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT6), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n554), .A2(new_n210), .A3(G107), .ZN(new_n555));
  XNOR2_X1  g0355(.A(G97), .B(G107), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n555), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  OAI22_X1  g0357(.A1(new_n557), .A2(new_n252), .B1(new_n208), .B2(new_n418), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n255), .B1(new_n356), .B2(new_n358), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n280), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n292), .A2(G97), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n286), .A2(new_n210), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(G244), .B(new_n300), .C1(new_n263), .C2(new_n264), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT4), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n270), .A2(KEYINPUT4), .A3(G244), .A4(new_n300), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n270), .A2(G250), .A3(G1698), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n494), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n305), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n304), .B1(new_n309), .B2(new_n311), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n317), .B1(new_n571), .B2(new_n211), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(G200), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n572), .B1(new_n569), .B2(new_n305), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G190), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n563), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n574), .A2(new_n449), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n576), .A2(new_n404), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n553), .A2(new_n578), .A3(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n306), .A2(new_n337), .A3(new_n312), .A4(new_n317), .ZN(new_n584));
  INV_X1    g0384(.A(new_n317), .ZN(new_n585));
  AOI211_X1 g0385(.A(new_n320), .B(new_n585), .C1(new_n302), .C2(new_n305), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n584), .B1(new_n586), .B2(G200), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n283), .A2(new_n293), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT82), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n283), .A2(new_n587), .A3(KEYINPUT82), .A4(new_n293), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n583), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AND4_X1   g0392(.A1(new_n328), .A2(new_n493), .A3(new_n520), .A4(new_n592), .ZN(new_n593));
  XNOR2_X1  g0393(.A(new_n593), .B(KEYINPUT83), .ZN(G372));
  INV_X1    g0394(.A(new_n447), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n446), .B1(new_n442), .B2(new_n443), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n388), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n598), .A2(new_n386), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT84), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n409), .A2(new_n600), .ZN(new_n601));
  OR2_X1    g0401(.A1(new_n408), .A2(G169), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n602), .A2(KEYINPUT84), .A3(new_n399), .A4(new_n407), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n491), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n488), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n599), .B1(new_n606), .B2(new_n381), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n461), .B1(new_n597), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(KEYINPUT85), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT85), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n610), .B(new_n461), .C1(new_n597), .C2(new_n607), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n582), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n613), .A2(KEYINPUT26), .A3(new_n553), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT26), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n542), .A2(new_n550), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n616), .B(new_n552), .C1(G169), .C2(new_n529), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n549), .A2(new_n411), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n618), .A2(new_n546), .A3(new_n542), .A4(new_n543), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n615), .B1(new_n620), .B2(new_n582), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n614), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n617), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n516), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n324), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n592), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n493), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n612), .A2(new_n629), .ZN(G369));
  INV_X1    g0430(.A(G330), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n285), .A2(G20), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  OR3_X1    g0433(.A1(new_n633), .A2(KEYINPUT27), .A3(G1), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT27), .B1(new_n633), .B2(G1), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(G213), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(G343), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n517), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n516), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n519), .A2(new_n517), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n625), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n644), .B(KEYINPUT86), .ZN(new_n645));
  AOI211_X1 g0445(.A(new_n631), .B(new_n642), .C1(new_n645), .C2(new_n641), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n294), .A2(new_n323), .A3(new_n638), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT87), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n294), .A2(KEYINPUT87), .A3(new_n323), .A4(new_n638), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n294), .A2(new_n638), .ZN(new_n652));
  AOI221_X4 g0452(.A(KEYINPUT81), .B1(new_n319), .B2(new_n322), .C1(new_n283), .C2(new_n293), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n326), .B1(new_n294), .B2(new_n323), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n590), .A2(new_n591), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n651), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n646), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n324), .A2(new_n638), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n625), .A2(new_n638), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n660), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n659), .A2(new_n662), .ZN(G399));
  NAND3_X1  g0463(.A1(new_n534), .A2(new_n535), .A3(new_n244), .ZN(new_n664));
  XOR2_X1   g0464(.A(new_n664), .B(KEYINPUT88), .Z(new_n665));
  INV_X1    g0465(.A(new_n223), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(G41), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n665), .A2(new_n307), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n230), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n668), .B1(new_n669), .B2(new_n667), .ZN(new_n670));
  XNOR2_X1  g0470(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n321), .A2(new_n576), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n529), .A2(G179), .A3(new_n507), .A4(new_n509), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT30), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n507), .A2(new_n509), .A3(G179), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(new_n549), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT30), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n677), .A2(new_n678), .A3(new_n321), .A4(new_n576), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n576), .A2(G179), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n681), .A2(new_n318), .A3(new_n510), .A4(new_n549), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n683), .A2(KEYINPUT31), .A3(new_n638), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n680), .A2(KEYINPUT90), .A3(new_n682), .ZN(new_n685));
  AOI21_X1  g0485(.A(KEYINPUT90), .B1(new_n680), .B2(new_n682), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n685), .A2(new_n686), .A3(new_n639), .ZN(new_n687));
  OAI211_X1 g0487(.A(KEYINPUT91), .B(new_n684), .C1(new_n687), .C2(KEYINPUT31), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n328), .A2(new_n592), .A3(new_n520), .A4(new_n639), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT90), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n683), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n680), .A2(KEYINPUT90), .A3(new_n682), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(new_n638), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT31), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(KEYINPUT91), .B1(new_n696), .B2(new_n684), .ZN(new_n697));
  OAI21_X1  g0497(.A(G330), .B1(new_n690), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n625), .B1(new_n653), .B2(new_n654), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n578), .A2(new_n582), .A3(new_n619), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n700), .B1(new_n590), .B2(new_n591), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n624), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n639), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT29), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n638), .B1(new_n624), .B2(new_n627), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n698), .B(new_n705), .C1(KEYINPUT29), .C2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n672), .B1(new_n709), .B2(G1), .ZN(G364));
  AOI21_X1  g0510(.A(new_n307), .B1(new_n632), .B2(G45), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n667), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n279), .B1(G20), .B2(new_n449), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n252), .A2(G190), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n411), .A2(new_n404), .A3(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(G179), .A2(G200), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI22_X1  g0522(.A1(new_n719), .A2(G283), .B1(G329), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT93), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n270), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n252), .A2(new_n337), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n404), .A2(G200), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G322), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n411), .A2(new_n404), .A3(new_n726), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT92), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G303), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n404), .A2(new_n349), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n726), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n252), .B1(new_n720), .B2(G190), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n737), .A2(G326), .B1(new_n739), .B2(G294), .ZN(new_n740));
  INV_X1    g0540(.A(G311), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n727), .A2(new_n717), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n735), .A2(new_n717), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  XNOR2_X1  g0545(.A(KEYINPUT94), .B(KEYINPUT33), .ZN(new_n746));
  INV_X1    g0546(.A(G317), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n746), .B(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n743), .B1(new_n745), .B2(new_n748), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n725), .A2(new_n730), .A3(new_n734), .A4(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n731), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n751), .A2(G87), .B1(G97), .B2(new_n739), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n270), .B1(new_n736), .B2(new_n202), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n753), .B1(new_n719), .B2(G107), .ZN(new_n754));
  INV_X1    g0554(.A(G159), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n721), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT32), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n728), .A2(new_n360), .B1(new_n742), .B2(new_n208), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(G68), .B2(new_n745), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n752), .A2(new_n754), .A3(new_n757), .A4(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n716), .B1(new_n750), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n715), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n666), .A2(new_n270), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(new_n250), .B2(G45), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(G45), .B2(new_n230), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n270), .A2(G355), .A3(new_n223), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n769), .B(new_n770), .C1(G116), .C2(new_n223), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n714), .B(new_n761), .C1(new_n765), .C2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n642), .B1(new_n645), .B2(new_n641), .ZN(new_n773));
  INV_X1    g0573(.A(new_n764), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n775), .A2(KEYINPUT95), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(KEYINPUT95), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n773), .A2(G330), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n773), .A2(G330), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n714), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n776), .A2(new_n777), .B1(new_n778), .B2(new_n780), .ZN(G396));
  NAND4_X1  g0581(.A1(new_n601), .A2(new_n603), .A3(new_n399), .A4(new_n638), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n399), .A2(new_n638), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n414), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n706), .B(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(new_n698), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n714), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT96), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n716), .A2(new_n763), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n713), .B1(new_n790), .B2(G77), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n785), .A2(new_n762), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n357), .B1(new_n732), .B2(new_n255), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT98), .Z(new_n794));
  XNOR2_X1  g0594(.A(KEYINPUT97), .B(G283), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n718), .A2(new_n535), .B1(new_n744), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n742), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G116), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n722), .A2(G311), .ZN(new_n801));
  INV_X1    g0601(.A(G294), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n728), .A2(new_n802), .B1(new_n738), .B2(new_n210), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT99), .Z(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(G303), .B2(new_n737), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n798), .A2(new_n800), .A3(new_n801), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n739), .A2(G58), .ZN(new_n807));
  INV_X1    g0607(.A(G132), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G143), .A2(new_n729), .B1(new_n799), .B2(G159), .ZN(new_n809));
  INV_X1    g0609(.A(G137), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n809), .B1(new_n810), .B2(new_n736), .C1(new_n417), .C2(new_n744), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT34), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n807), .B1(new_n808), .B2(new_n721), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n719), .A2(G68), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n733), .A2(G50), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n357), .B1(new_n811), .B2(new_n812), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n814), .A2(new_n815), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n806), .A2(new_n818), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n792), .B1(new_n789), .B2(new_n791), .C1(new_n819), .C2(new_n716), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n788), .A2(new_n820), .ZN(G384));
  NAND4_X1  g0621(.A1(new_n692), .A2(KEYINPUT31), .A3(new_n638), .A4(new_n693), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n689), .A2(new_n696), .A3(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n785), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n487), .A2(new_n638), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n488), .A2(new_n491), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n477), .A2(new_n487), .A3(new_n638), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n823), .A2(new_n824), .A3(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT103), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OR2_X1    g0631(.A1(KEYINPUT103), .A2(KEYINPUT40), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n823), .A2(new_n824), .A3(new_n828), .A4(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n378), .A2(new_n636), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n353), .A2(new_n378), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT17), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n353), .A2(new_n378), .A3(KEYINPUT17), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n834), .B1(new_n839), .B2(new_n599), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT37), .ZN(new_n841));
  INV_X1    g0641(.A(new_n636), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n382), .B1(new_n385), .B2(new_n842), .ZN(new_n843));
  AOI211_X1 g0643(.A(KEYINPUT100), .B(new_n841), .C1(new_n835), .C2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n835), .A2(new_n843), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(KEYINPUT37), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n835), .A2(new_n841), .A3(new_n843), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n847), .A2(KEYINPUT100), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n840), .A2(new_n845), .A3(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT38), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n840), .A2(new_n849), .A3(KEYINPUT38), .A4(new_n845), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n831), .A2(new_n833), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n847), .A2(KEYINPUT101), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n848), .A2(KEYINPUT102), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT102), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n835), .A2(new_n843), .A3(new_n858), .A4(new_n841), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT101), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n846), .A2(new_n860), .A3(KEYINPUT37), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n856), .A2(new_n857), .A3(new_n859), .A4(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT38), .B1(new_n862), .B2(new_n840), .ZN(new_n863));
  INV_X1    g0663(.A(new_n853), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT40), .B1(new_n865), .B2(new_n833), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n855), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n493), .A2(new_n823), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(G330), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n867), .B2(new_n869), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n599), .A2(new_n636), .ZN(new_n872));
  INV_X1    g0672(.A(new_n854), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n409), .A2(new_n638), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(new_n706), .B2(new_n824), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n828), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n844), .B1(new_n390), .B2(new_n834), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT38), .B1(new_n878), .B2(new_n849), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT39), .B1(new_n879), .B2(new_n864), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT39), .ZN(new_n881));
  INV_X1    g0681(.A(new_n834), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n381), .B2(new_n389), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n857), .A2(new_n859), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n860), .B1(new_n846), .B2(KEYINPUT37), .ZN(new_n885));
  AOI211_X1 g0685(.A(KEYINPUT101), .B(new_n841), .C1(new_n835), .C2(new_n843), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n883), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n881), .B(new_n853), .C1(new_n888), .C2(KEYINPUT38), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n880), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n477), .A2(new_n487), .A3(new_n639), .ZN(new_n891));
  OAI221_X1 g0691(.A(new_n872), .B1(new_n873), .B2(new_n877), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n871), .B(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n705), .B1(KEYINPUT29), .B2(new_n707), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n493), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n612), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n893), .B(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n307), .B2(new_n632), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT35), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n228), .B1(new_n557), .B2(new_n899), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n900), .B(G116), .C1(new_n899), .C2(new_n557), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT36), .ZN(new_n902));
  OAI21_X1  g0702(.A(G77), .B1(new_n360), .B2(new_n218), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n230), .A2(new_n903), .B1(G50), .B2(new_n218), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n904), .A2(G1), .A3(new_n285), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n898), .A2(new_n902), .A3(new_n905), .ZN(G367));
  NAND2_X1  g0706(.A1(new_n658), .A2(new_n661), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n578), .B(new_n582), .C1(new_n563), .C2(new_n639), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n613), .A2(new_n638), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  OR3_X1    g0711(.A1(new_n907), .A2(KEYINPUT42), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n582), .B1(new_n328), .B2(new_n908), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n639), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT42), .B1(new_n907), .B2(new_n911), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n912), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n544), .A2(new_n638), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n553), .A2(new_n917), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n617), .A2(new_n917), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(KEYINPUT43), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n916), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n920), .A2(KEYINPUT43), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n659), .A2(new_n911), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n922), .A2(new_n923), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n925), .B1(new_n924), .B2(new_n926), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n667), .B(KEYINPUT41), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  XOR2_X1   g0731(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n662), .B2(new_n910), .ZN(new_n933));
  INV_X1    g0733(.A(new_n661), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n656), .B(new_n652), .C1(new_n654), .C2(new_n653), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n934), .B1(new_n935), .B2(new_n651), .ZN(new_n936));
  INV_X1    g0736(.A(new_n932), .ZN(new_n937));
  NOR4_X1   g0737(.A1(new_n936), .A2(new_n660), .A3(new_n911), .A4(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n933), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT44), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n662), .B2(new_n910), .ZN(new_n941));
  OAI211_X1 g0741(.A(KEYINPUT44), .B(new_n911), .C1(new_n936), .C2(new_n660), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AND3_X1   g0743(.A1(new_n939), .A2(new_n659), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n659), .B1(new_n939), .B2(new_n943), .ZN(new_n945));
  OAI21_X1  g0745(.A(KEYINPUT105), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n659), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n947), .A2(KEYINPUT105), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n935), .A2(new_n651), .A3(new_n934), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n936), .A2(KEYINPUT106), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT106), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n907), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n779), .A2(new_n949), .A3(new_n950), .A4(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n952), .A2(new_n949), .A3(new_n950), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n646), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n708), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n946), .A2(new_n948), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n931), .B1(new_n957), .B2(new_n709), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n929), .B1(new_n958), .B2(new_n712), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n738), .A2(new_n218), .ZN(new_n960));
  XNOR2_X1  g0760(.A(KEYINPUT108), .B(G137), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n731), .A2(new_n360), .B1(new_n721), .B2(new_n962), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n960), .B(new_n963), .C1(G143), .C2(new_n737), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n270), .B1(new_n202), .B2(new_n742), .C1(new_n718), .C2(new_n208), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(G150), .B2(new_n729), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n964), .B(new_n966), .C1(new_n755), .C2(new_n744), .ZN(new_n967));
  OAI21_X1  g0767(.A(KEYINPUT46), .B1(new_n732), .B2(new_n244), .ZN(new_n968));
  OR3_X1    g0768(.A1(new_n731), .A2(KEYINPUT46), .A3(new_n244), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n357), .B1(new_n744), .B2(new_n802), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(new_n799), .B2(new_n795), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n718), .A2(new_n210), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(G107), .B2(new_n739), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n722), .A2(G317), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n970), .A2(new_n972), .A3(new_n974), .A4(new_n975), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n736), .A2(new_n741), .B1(new_n728), .B2(new_n505), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT107), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n967), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT47), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n715), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n765), .B1(new_n223), .B2(new_n396), .C1(new_n241), .C2(new_n767), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n918), .A2(new_n764), .A3(new_n919), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n981), .A2(new_n713), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n959), .A2(new_n984), .ZN(G387));
  NAND2_X1  g0785(.A1(new_n953), .A2(new_n955), .ZN(new_n986));
  AOI22_X1  g0786(.A1(G322), .A2(new_n737), .B1(new_n745), .B2(G311), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n987), .B1(new_n505), .B2(new_n742), .C1(new_n747), .C2(new_n728), .ZN(new_n988));
  XOR2_X1   g0788(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n989));
  XNOR2_X1  g0789(.A(new_n988), .B(new_n989), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n802), .B2(new_n731), .C1(new_n738), .C2(new_n796), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT49), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n719), .A2(G116), .B1(G326), .B2(new_n722), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n992), .A2(new_n357), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n270), .B1(new_n721), .B2(new_n417), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n995), .B(new_n973), .C1(G68), .C2(new_n799), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n396), .A2(new_n738), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n731), .A2(new_n208), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n997), .B(new_n998), .C1(new_n375), .C2(new_n745), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n729), .A2(G50), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n737), .A2(G159), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n996), .A2(new_n999), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n716), .B1(new_n994), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n665), .B1(G68), .B2(G77), .ZN(new_n1004));
  INV_X1    g0804(.A(G45), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n374), .A2(G50), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT50), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1004), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n767), .B1(new_n238), .B2(G45), .ZN(new_n1009));
  AND3_X1   g0809(.A1(new_n665), .A2(new_n223), .A3(new_n270), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1008), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n666), .A2(new_n255), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n714), .B(new_n1003), .C1(new_n765), .C2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n935), .A2(new_n651), .A3(new_n764), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n712), .A2(new_n986), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n667), .B1(new_n709), .B2(new_n986), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1016), .B1(new_n1017), .B2(new_n956), .ZN(G393));
  OAI21_X1  g0818(.A(KEYINPUT110), .B1(new_n944), .B2(new_n945), .ZN(new_n1019));
  AND2_X1   g0819(.A1(new_n941), .A2(new_n942), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n660), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n907), .A2(new_n1021), .A3(new_n910), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n937), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n662), .A2(new_n910), .A3(new_n932), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n947), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT110), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n939), .A2(new_n659), .A3(new_n943), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1019), .A2(new_n712), .A3(new_n1029), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n736), .A2(new_n747), .B1(new_n728), .B2(new_n741), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT111), .Z(new_n1032));
  OAI22_X1  g0832(.A1(new_n1032), .A2(KEYINPUT52), .B1(new_n802), .B2(new_n742), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(KEYINPUT52), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n719), .A2(G107), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(G322), .A2(new_n722), .B1(new_n739), .B2(G116), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n270), .B1(new_n751), .B2(new_n795), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n1033), .B(new_n1038), .C1(G303), .C2(new_n745), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G150), .A2(new_n737), .B1(new_n729), .B2(G159), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n270), .B1(new_n202), .B2(new_n744), .C1(new_n1040), .C2(KEYINPUT51), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G68), .A2(new_n751), .B1(new_n719), .B2(G87), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1040), .A2(KEYINPUT51), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n738), .A2(new_n208), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G143), .B2(new_n722), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1042), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1041), .B(new_n1046), .C1(new_n375), .C2(new_n799), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n715), .B1(new_n1039), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n911), .A2(new_n764), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n247), .A2(new_n766), .B1(G97), .B2(new_n666), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n765), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1048), .A2(new_n1049), .A3(new_n713), .A4(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1030), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n956), .B1(new_n1028), .B2(new_n1026), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n709), .A2(new_n986), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1055), .B1(new_n1056), .B2(KEYINPUT105), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1054), .B1(new_n1057), .B2(new_n948), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1053), .B1(new_n1058), .B2(new_n667), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(G390));
  INV_X1    g0860(.A(new_n828), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n891), .B1(new_n875), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1062), .A2(new_n880), .A3(new_n889), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n853), .B1(new_n888), .B2(KEYINPUT38), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n891), .B(KEYINPUT112), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n703), .A2(new_n639), .A3(new_n824), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n874), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1061), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1067), .A2(new_n1070), .A3(KEYINPUT113), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT113), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n857), .A2(new_n859), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n1073), .A2(new_n885), .A3(new_n886), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n851), .B1(new_n1074), .B2(new_n883), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1065), .B1(new_n1075), .B2(new_n853), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n638), .B(new_n785), .C1(new_n702), .C2(new_n624), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n828), .B1(new_n1077), .B2(new_n874), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1072), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1063), .B1(new_n1071), .B2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n829), .A2(new_n631), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n493), .A2(G330), .A3(new_n823), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n895), .A2(new_n612), .A3(new_n1083), .ZN(new_n1084));
  OAI211_X1 g0884(.A(G330), .B(new_n824), .C1(new_n690), .C2(new_n697), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n1061), .ZN(new_n1086));
  AND3_X1   g0886(.A1(new_n823), .A2(new_n824), .A3(new_n828), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(G330), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n876), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1077), .A2(new_n874), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n823), .A2(G330), .A3(new_n824), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n1061), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1091), .B(new_n1093), .C1(new_n1085), .C2(new_n1061), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1084), .B1(new_n1090), .B2(new_n1094), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1085), .A2(new_n1061), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1096), .B(new_n1063), .C1(new_n1071), .C2(new_n1079), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1082), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n667), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT114), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(KEYINPUT113), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1076), .A2(new_n1078), .A3(new_n1072), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1102), .A2(new_n1103), .B1(new_n890), .B2(new_n1062), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1097), .B1(new_n1104), .B2(new_n1088), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1084), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1081), .B1(new_n1061), .B2(new_n1085), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1094), .B1(new_n1107), .B2(new_n875), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g0910(.A(KEYINPUT114), .B(new_n667), .C1(new_n1105), .C2(new_n1109), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1101), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n890), .A2(new_n762), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n790), .A2(new_n375), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n731), .A2(new_n417), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  XOR2_X1   g0917(.A(KEYINPUT54), .B(G143), .Z(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n1119), .A2(new_n742), .B1(new_n808), .B2(new_n728), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(G128), .B2(new_n737), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n357), .B1(new_n722), .B2(G125), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n962), .A2(new_n744), .B1(new_n738), .B2(new_n755), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n719), .B2(G50), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1117), .A2(new_n1121), .A3(new_n1122), .A4(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(G283), .A2(new_n737), .B1(new_n799), .B2(G97), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n255), .B2(new_n744), .ZN(new_n1127));
  OR2_X1    g0927(.A1(new_n1127), .A2(KEYINPUT116), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n733), .A2(G87), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n1127), .A2(KEYINPUT116), .B1(G68), .B2(new_n719), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n270), .B(new_n1044), .C1(G116), .C2(new_n729), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n721), .A2(new_n802), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1125), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  XOR2_X1   g0934(.A(new_n1134), .B(KEYINPUT117), .Z(new_n1135));
  AOI211_X1 g0935(.A(new_n714), .B(new_n1114), .C1(new_n1135), .C2(new_n715), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1113), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n1105), .B2(new_n711), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1112), .A2(new_n1139), .ZN(G378));
  XNOR2_X1  g0940(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n422), .A2(new_n842), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n448), .A2(new_n461), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1143), .B1(new_n448), .B2(new_n461), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1142), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n448), .A2(new_n461), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1143), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n448), .A2(new_n461), .A3(new_n1143), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1149), .A2(new_n1150), .A3(new_n1141), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1146), .A2(new_n1151), .A3(KEYINPUT120), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n867), .A2(G330), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1152), .B1(new_n867), .B2(G330), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n892), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1152), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1087), .A2(new_n1064), .A3(new_n832), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n829), .A2(new_n830), .B1(new_n853), .B2(new_n852), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(KEYINPUT40), .A2(new_n1157), .B1(new_n1158), .B2(new_n833), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1156), .B1(new_n1159), .B2(new_n631), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n890), .A2(new_n891), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n872), .B1(new_n877), .B2(new_n873), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n867), .A2(new_n1152), .A3(G330), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1160), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1155), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1146), .A2(new_n1151), .A3(new_n762), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n713), .B1(new_n790), .B2(G50), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n718), .A2(new_n360), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n736), .A2(new_n244), .B1(new_n728), .B2(new_n255), .ZN(new_n1170));
  OR2_X1    g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(G283), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n721), .A2(new_n1172), .ZN(new_n1173));
  NOR4_X1   g0973(.A1(new_n1171), .A2(new_n960), .A3(new_n998), .A4(new_n1173), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n396), .A2(new_n742), .B1(new_n210), .B2(new_n744), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT118), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1174), .A2(new_n310), .A3(new_n357), .A4(new_n1176), .ZN(new_n1177));
  XOR2_X1   g0977(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n1178));
  XNOR2_X1  g0978(.A(new_n1177), .B(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n202), .B1(new_n263), .B2(G41), .ZN(new_n1180));
  INV_X1    g0980(.A(G124), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n290), .B1(new_n721), .B2(new_n1181), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n751), .A2(new_n1118), .B1(G125), .B2(new_n737), .ZN(new_n1183));
  INV_X1    g0983(.A(G128), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n728), .A2(new_n1184), .B1(new_n742), .B2(new_n810), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G150), .B2(new_n739), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1183), .B(new_n1186), .C1(new_n808), .C2(new_n744), .ZN(new_n1187));
  AOI211_X1 g0987(.A(G41), .B(new_n1182), .C1(new_n1187), .C2(KEYINPUT59), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1188), .B1(KEYINPUT59), .B2(new_n1187), .C1(new_n755), .C2(new_n718), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1179), .A2(new_n1180), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1168), .B1(new_n1190), .B2(new_n715), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n1166), .A2(new_n712), .B1(new_n1167), .B2(new_n1191), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1098), .A2(new_n1106), .B1(new_n1155), .B2(new_n1165), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n667), .B1(new_n1193), .B2(KEYINPUT57), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1106), .B1(new_n1105), .B2(new_n1109), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n1166), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT57), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1192), .B1(new_n1194), .B2(new_n1198), .ZN(G375));
  AOI22_X1  g0999(.A1(new_n719), .A2(G77), .B1(G116), .B2(new_n745), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1200), .B(new_n357), .C1(new_n255), .C2(new_n742), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n728), .A2(new_n1172), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n721), .A2(new_n505), .ZN(new_n1203));
  NOR4_X1   g1003(.A1(new_n1201), .A2(new_n997), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n210), .B2(new_n732), .C1(new_n802), .C2(new_n736), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT121), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G132), .A2(new_n737), .B1(new_n745), .B2(new_n1118), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n728), .B2(new_n962), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT122), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n357), .B1(new_n733), .B2(G159), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n742), .A2(new_n417), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1211), .B(new_n1169), .C1(G50), .C2(new_n739), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1210), .B(new_n1212), .C1(new_n1184), .C2(new_n721), .ZN(new_n1213));
  XOR2_X1   g1013(.A(new_n1213), .B(KEYINPUT123), .Z(new_n1214));
  OAI21_X1  g1014(.A(new_n1206), .B1(new_n1209), .B2(new_n1214), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT124), .Z(new_n1216));
  OAI221_X1 g1016(.A(new_n713), .B1(G68), .B2(new_n790), .C1(new_n1216), .C2(new_n716), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n762), .B2(new_n1061), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n712), .B2(new_n1108), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1090), .A2(new_n1084), .A3(new_n1094), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1109), .A2(new_n1220), .A3(new_n930), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1219), .A2(new_n1221), .ZN(G381));
  NOR2_X1   g1022(.A1(G375), .A2(G378), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n959), .A2(new_n984), .A3(new_n1059), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(G384), .ZN(new_n1227));
  INV_X1    g1027(.A(G381), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(G393), .A2(G396), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .A4(new_n1229), .ZN(G407));
  OAI211_X1 g1030(.A(G407), .B(G213), .C1(G343), .C2(new_n1224), .ZN(G409));
  NAND2_X1  g1031(.A1(new_n637), .A2(G213), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1193), .A2(new_n930), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1112), .A2(new_n1139), .A3(new_n1192), .A4(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1166), .A2(new_n712), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1167), .A2(new_n1191), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n667), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1193), .A2(KEYINPUT57), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1237), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1111), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT114), .B1(new_n1098), .B2(new_n667), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1138), .B1(new_n1244), .B2(new_n1110), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1232), .B(new_n1234), .C1(new_n1241), .C2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT60), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1220), .A2(new_n1247), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1090), .A2(new_n1084), .A3(KEYINPUT60), .A4(new_n1094), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1248), .A2(new_n667), .A3(new_n1109), .A4(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1219), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1227), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1250), .A2(new_n1219), .A3(G384), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT62), .B1(new_n1246), .B2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n637), .A2(G213), .A3(G2897), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1256), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1252), .A2(new_n1253), .A3(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT61), .B1(new_n1246), .B2(new_n1260), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(G375), .A2(G378), .B1(G213), .B2(new_n637), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT62), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1254), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .A4(new_n1234), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1255), .A2(new_n1261), .A3(new_n1265), .ZN(new_n1266));
  XOR2_X1   g1066(.A(G393), .B(G396), .Z(new_n1267));
  NAND2_X1  g1067(.A1(new_n1225), .A2(KEYINPUT127), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1059), .B1(new_n959), .B2(new_n984), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1267), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(G387), .A2(G390), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1267), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1271), .A2(KEYINPUT127), .A3(new_n1225), .A4(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1266), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1246), .A2(KEYINPUT125), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT126), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1252), .A2(new_n1253), .A3(new_n1258), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1258), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1277), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1257), .A2(new_n1259), .A3(KEYINPUT126), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(G375), .A2(G378), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT125), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1283), .A2(new_n1284), .A3(new_n1232), .A4(new_n1234), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1276), .A2(new_n1282), .A3(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT63), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1287), .B1(new_n1246), .B2(new_n1254), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1262), .A2(KEYINPUT63), .A3(new_n1264), .A4(new_n1234), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT61), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1270), .A2(new_n1290), .A3(new_n1273), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1286), .A2(new_n1288), .A3(new_n1289), .A4(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1275), .A2(new_n1292), .ZN(G405));
  NAND2_X1  g1093(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1294), .A2(new_n1240), .A3(new_n667), .ZN(new_n1295));
  AOI22_X1  g1095(.A1(new_n1295), .A2(new_n1192), .B1(new_n1139), .B2(new_n1112), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1223), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1274), .A2(new_n1297), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1270), .B(new_n1273), .C1(new_n1223), .C2(new_n1296), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1298), .A2(new_n1264), .A3(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1264), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(G402));
endmodule


