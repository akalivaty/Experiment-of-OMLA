//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n808, new_n809, new_n810, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(KEYINPUT23), .ZN(new_n203));
  NAND2_X1  g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT65), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT65), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n206), .A2(G169gat), .A3(G176gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n202), .A2(KEYINPUT23), .ZN(new_n209));
  AND3_X1   g008(.A1(new_n203), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n212));
  INV_X1    g011(.A(G183gat), .ZN(new_n213));
  INV_X1    g012(.A(G190gat), .ZN(new_n214));
  AOI22_X1  g013(.A1(new_n211), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT24), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n215), .B(new_n218), .C1(new_n212), .C2(new_n211), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT25), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n210), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n216), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n208), .A2(KEYINPUT69), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT69), .B1(new_n208), .B2(new_n224), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT26), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n202), .A2(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n223), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT27), .B(G183gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(new_n214), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT28), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n232), .A2(KEYINPUT68), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(KEYINPUT68), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n231), .A2(new_n214), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n222), .B1(new_n230), .B2(new_n237), .ZN(new_n238));
  XOR2_X1   g037(.A(G127gat), .B(G134gat), .Z(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(KEYINPUT71), .B(KEYINPUT1), .Z(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT70), .B(G120gat), .ZN(new_n242));
  INV_X1    g041(.A(G113gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n243), .A2(G120gat), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n240), .B(new_n241), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G113gat), .B(G120gat), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n239), .B1(KEYINPUT1), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n251), .A2(new_n213), .A3(new_n214), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n252), .A2(new_n218), .A3(new_n253), .A4(new_n211), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT67), .ZN(new_n255));
  AND2_X1   g054(.A1(new_n253), .A2(new_n211), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n256), .A2(new_n257), .A3(new_n218), .A4(new_n252), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n210), .A2(new_n255), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT25), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n238), .A2(KEYINPUT72), .A3(new_n250), .A4(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n208), .A2(new_n224), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n208), .A2(KEYINPUT69), .A3(new_n224), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(new_n229), .A3(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(new_n216), .A3(new_n237), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n267), .A2(new_n260), .A3(new_n221), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n249), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT72), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n270), .B1(new_n268), .B2(new_n249), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n261), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(G227gat), .A2(G233gat), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT32), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT33), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G15gat), .B(G43gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(G71gat), .ZN(new_n280));
  INV_X1    g079(.A(G99gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n276), .A2(new_n278), .A3(new_n282), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n261), .A2(new_n271), .A3(new_n273), .A4(new_n269), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT34), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT32), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n287), .B1(new_n272), .B2(new_n274), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT33), .B1(new_n272), .B2(new_n274), .ZN(new_n289));
  INV_X1    g088(.A(new_n282), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n283), .A2(new_n286), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT74), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n283), .A2(new_n286), .A3(KEYINPUT74), .A4(new_n291), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AND2_X1   g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G141gat), .B(G148gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT2), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n301), .B1(G155gat), .B2(G162gat), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n299), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G148gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G141gat), .ZN(new_n305));
  INV_X1    g104(.A(G141gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G148gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G155gat), .B(G162gat), .ZN(new_n309));
  INV_X1    g108(.A(G155gat), .ZN(new_n310));
  INV_X1    g109(.A(G162gat), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT2), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n308), .A2(new_n309), .A3(new_n312), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n303), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n314), .A2(new_n246), .A3(new_n248), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT4), .ZN(new_n317));
  NAND2_X1  g116(.A1(G225gat), .A2(G233gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT3), .ZN(new_n320));
  AND3_X1   g119(.A1(new_n303), .A2(new_n313), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n320), .B1(new_n303), .B2(new_n313), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n319), .B1(new_n323), .B2(new_n249), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n317), .B(new_n318), .C1(new_n324), .C2(new_n316), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n303), .A2(new_n313), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n249), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT78), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(new_n328), .A3(new_n315), .ZN(new_n329));
  INV_X1    g128(.A(new_n318), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n249), .A2(KEYINPUT78), .A3(new_n326), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n325), .A2(KEYINPUT5), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n321), .ZN(new_n334));
  INV_X1    g133(.A(new_n322), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n334), .A2(new_n249), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n336), .A2(KEYINPUT4), .A3(new_n315), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n316), .A2(new_n319), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT5), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(new_n340), .A3(new_n318), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n333), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n343));
  XNOR2_X1  g142(.A(G57gat), .B(G85gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G1gat), .B(G29gat), .ZN(new_n346));
  XOR2_X1   g145(.A(new_n345), .B(new_n346), .Z(new_n347));
  NAND2_X1  g146(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT6), .ZN(new_n349));
  INV_X1    g148(.A(new_n347), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n333), .A2(new_n341), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n348), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n342), .A2(KEYINPUT6), .A3(new_n347), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(G211gat), .A2(G218gat), .ZN(new_n355));
  OR2_X1    g154(.A1(G211gat), .A2(G218gat), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT22), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G197gat), .B(G204gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT75), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n356), .A2(new_n355), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n362), .B1(KEYINPUT22), .B2(new_n359), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G226gat), .A2(G233gat), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n268), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT29), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n268), .A2(new_n369), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n365), .B(new_n368), .C1(new_n370), .C2(new_n367), .ZN(new_n371));
  INV_X1    g170(.A(new_n368), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n367), .B1(new_n268), .B2(new_n369), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n364), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G8gat), .B(G36gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(G64gat), .B(G92gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n371), .A2(new_n374), .A3(KEYINPUT30), .A4(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n378), .B1(new_n371), .B2(new_n374), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT76), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n371), .A2(new_n374), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n377), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT76), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n385), .A3(new_n379), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n371), .A2(new_n374), .A3(new_n378), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT30), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AND4_X1   g188(.A1(new_n354), .A2(new_n382), .A3(new_n386), .A4(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT31), .B(G50gat), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n364), .B1(KEYINPUT29), .B2(new_n321), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT3), .B1(new_n365), .B2(new_n369), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n392), .B1(new_n393), .B2(new_n314), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(G78gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n394), .A2(G78gat), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n391), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OR2_X1    g197(.A1(new_n394), .A2(G78gat), .ZN(new_n399));
  INV_X1    g198(.A(new_n391), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(new_n400), .A3(new_n395), .ZN(new_n401));
  NAND2_X1  g200(.A1(G228gat), .A2(G233gat), .ZN(new_n402));
  INV_X1    g201(.A(G22gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(G106gat), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n398), .A2(new_n401), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n405), .B1(new_n398), .B2(new_n401), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR3_X1   g207(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n409));
  AOI221_X4 g208(.A(new_n287), .B1(KEYINPUT33), .B2(new_n282), .C1(new_n272), .C2(new_n274), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT73), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n286), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT73), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n283), .A2(new_n413), .A3(new_n291), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n411), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n296), .A2(new_n390), .A3(new_n408), .A4(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT35), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n283), .A2(new_n291), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n412), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n389), .A2(new_n384), .A3(new_n379), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT35), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n420), .A2(new_n421), .A3(new_n354), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n296), .A2(new_n419), .A3(new_n408), .A4(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT81), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n294), .A2(new_n295), .B1(new_n412), .B2(new_n418), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n426), .A2(KEYINPUT81), .A3(new_n408), .A4(new_n422), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n417), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n296), .A2(new_n415), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT36), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT36), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  OR2_X1    g231(.A1(new_n390), .A2(new_n408), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n337), .A2(new_n330), .A3(new_n338), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n434), .A2(KEYINPUT39), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n435), .A2(new_n347), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n329), .A2(new_n331), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n434), .B(KEYINPUT39), .C1(new_n437), .C2(new_n330), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT40), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT80), .ZN(new_n440));
  OR2_X1    g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n439), .A2(new_n440), .B1(new_n347), .B2(new_n342), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n389), .A2(new_n384), .A3(new_n379), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n436), .A2(KEYINPUT40), .A3(new_n438), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n441), .A2(new_n442), .A3(new_n443), .A4(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n354), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT38), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT37), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n383), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n371), .A2(new_n374), .A3(KEYINPUT37), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n378), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n446), .B1(new_n447), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n447), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n387), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n408), .B(new_n445), .C1(new_n452), .C2(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n430), .A2(new_n432), .A3(new_n433), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n428), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT94), .ZN(new_n458));
  NAND2_X1  g257(.A1(G85gat), .A2(G92gat), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT7), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT90), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT90), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT7), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n460), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT91), .B1(new_n459), .B2(KEYINPUT7), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n460), .A2(new_n462), .A3(new_n464), .A4(KEYINPUT91), .ZN(new_n468));
  NAND2_X1  g267(.A1(G99gat), .A2(G106gat), .ZN(new_n469));
  INV_X1    g268(.A(G85gat), .ZN(new_n470));
  INV_X1    g269(.A(G92gat), .ZN(new_n471));
  AOI22_X1  g270(.A1(KEYINPUT8), .A2(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n467), .A2(new_n468), .A3(new_n472), .ZN(new_n473));
  XOR2_X1   g272(.A(G99gat), .B(G106gat), .Z(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n474), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n467), .A2(new_n476), .A3(new_n468), .A4(new_n472), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(KEYINPUT92), .A3(new_n477), .ZN(new_n478));
  OR3_X1    g277(.A1(new_n473), .A2(KEYINPUT92), .A3(new_n474), .ZN(new_n479));
  NOR2_X1   g278(.A1(G29gat), .A2(G36gat), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT14), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n480), .B(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(G29gat), .A2(G36gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G43gat), .B(G50gat), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(KEYINPUT15), .A3(new_n485), .ZN(new_n486));
  OR2_X1    g285(.A1(new_n485), .A2(KEYINPUT15), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(KEYINPUT15), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n483), .B(KEYINPUT83), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n487), .A2(new_n482), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT17), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n486), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n491), .B1(new_n486), .B2(new_n490), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n478), .B(new_n479), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n486), .A2(new_n490), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n494), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G190gat), .B(G218gat), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n494), .A2(new_n497), .A3(new_n498), .A4(new_n500), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(KEYINPUT93), .A3(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G134gat), .B(G162gat), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n502), .A2(KEYINPUT93), .A3(new_n503), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT93), .B1(new_n502), .B2(new_n503), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n509), .B1(new_n512), .B2(new_n508), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT89), .B(G183gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(G127gat), .B(G155gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G15gat), .B(G22gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT84), .ZN(new_n519));
  INV_X1    g318(.A(G1gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n518), .A2(KEYINPUT84), .A3(G1gat), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT16), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  OR2_X1    g324(.A1(new_n518), .A2(G1gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT85), .ZN(new_n527));
  AOI21_X1  g326(.A(G8gat), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(G8gat), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n518), .A2(G1gat), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n530), .B1(new_n531), .B2(KEYINPUT85), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n532), .A2(new_n521), .A3(new_n522), .A4(new_n524), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT86), .ZN(new_n535));
  XNOR2_X1  g334(.A(G57gat), .B(G64gat), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  XOR2_X1   g337(.A(G71gat), .B(G78gat), .Z(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT21), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n534), .A2(new_n541), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n538), .A2(new_n539), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n538), .A2(new_n539), .ZN(new_n544));
  XOR2_X1   g343(.A(KEYINPUT87), .B(KEYINPUT21), .Z(new_n545));
  OR3_X1    g344(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G231gat), .A2(G233gat), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n549), .B(KEYINPUT88), .Z(new_n550));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n546), .A3(new_n541), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n550), .B1(new_n548), .B2(new_n551), .ZN(new_n554));
  XNOR2_X1  g353(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n555));
  INV_X1    g354(.A(G211gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NOR3_X1   g356(.A1(new_n553), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n557), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n548), .A2(new_n551), .ZN(new_n560));
  INV_X1    g359(.A(new_n550), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n559), .B1(new_n562), .B2(new_n552), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n517), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n557), .B1(new_n553), .B2(new_n554), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n562), .A2(new_n552), .A3(new_n559), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(new_n516), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n458), .B1(new_n513), .B2(new_n568), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n564), .A2(new_n567), .ZN(new_n570));
  INV_X1    g369(.A(new_n511), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n571), .A2(new_n504), .A3(new_n508), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n510), .A2(new_n507), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n570), .A2(new_n574), .A3(KEYINPUT94), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n569), .A2(new_n575), .ZN(new_n576));
  AND2_X1   g375(.A1(new_n457), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n540), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n478), .A2(new_n479), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT10), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n540), .A2(new_n475), .A3(new_n477), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n495), .A2(KEYINPUT10), .A3(new_n540), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G230gat), .A2(G233gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n585), .B1(new_n579), .B2(new_n581), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G120gat), .B(G148gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(G176gat), .B(G204gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n586), .A2(new_n588), .A3(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n585), .B(KEYINPUT95), .Z(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n595), .B1(new_n582), .B2(new_n583), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n591), .B1(new_n596), .B2(new_n587), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n593), .A2(KEYINPUT96), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT96), .ZN(new_n599));
  OAI211_X1 g398(.A(new_n599), .B(new_n591), .C1(new_n596), .C2(new_n587), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n534), .B1(new_n492), .B2(new_n493), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n496), .A2(new_n529), .A3(new_n533), .ZN(new_n604));
  NAND2_X1  g403(.A1(G229gat), .A2(G233gat), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT18), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n605), .B(KEYINPUT13), .Z(new_n609));
  INV_X1    g408(.A(new_n604), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n496), .B1(new_n529), .B2(new_n533), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n603), .A2(KEYINPUT18), .A3(new_n604), .A4(new_n605), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n608), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G169gat), .B(G197gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G113gat), .B(G141gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n614), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n608), .A2(new_n620), .A3(new_n612), .A4(new_n613), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n602), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n577), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n446), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g428(.A1(new_n627), .A2(new_n443), .ZN(new_n630));
  NAND2_X1  g429(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n523), .A2(new_n530), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT42), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n635), .B(new_n636), .C1(new_n530), .C2(new_n630), .ZN(G1325gat));
  AOI21_X1  g436(.A(G15gat), .B1(new_n627), .B2(new_n426), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n430), .A2(new_n432), .ZN(new_n639));
  AND2_X1   g438(.A1(new_n639), .A2(G15gat), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n638), .B1(new_n627), .B2(new_n640), .ZN(G1326gat));
  INV_X1    g440(.A(new_n408), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(new_n403), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT97), .B(KEYINPUT43), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(G1327gat));
  AOI21_X1  g445(.A(new_n574), .B1(new_n428), .B2(new_n456), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n647), .A2(KEYINPUT99), .A3(KEYINPUT44), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT44), .B1(new_n647), .B2(KEYINPUT99), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n648), .A2(new_n649), .A3(new_n570), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n601), .B(KEYINPUT98), .Z(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n650), .A2(new_n624), .A3(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(G29gat), .B1(new_n653), .B2(new_n354), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n647), .A2(new_n626), .A3(new_n568), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n655), .A2(G29gat), .A3(new_n354), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n656), .B(KEYINPUT45), .Z(new_n657));
  NAND2_X1  g456(.A1(new_n654), .A2(new_n657), .ZN(G1328gat));
  OR3_X1    g457(.A1(new_n653), .A2(KEYINPUT100), .A3(new_n420), .ZN(new_n659));
  OAI21_X1  g458(.A(KEYINPUT100), .B1(new_n653), .B2(new_n420), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n659), .A2(G36gat), .A3(new_n660), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n655), .A2(G36gat), .A3(new_n420), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT46), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(G1329gat));
  INV_X1    g463(.A(new_n426), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n655), .A2(G43gat), .A3(new_n665), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n650), .A2(new_n624), .A3(new_n639), .A4(new_n652), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n666), .B1(new_n667), .B2(G43gat), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT47), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n668), .A2(KEYINPUT101), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n666), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n457), .A2(KEYINPUT99), .A3(new_n513), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n647), .A2(KEYINPUT99), .A3(KEYINPUT44), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n674), .A2(new_n624), .A3(new_n568), .A4(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n639), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n676), .A2(new_n677), .A3(new_n651), .ZN(new_n678));
  INV_X1    g477(.A(G43gat), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n671), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT101), .ZN(new_n681));
  AOI21_X1  g480(.A(KEYINPUT47), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n670), .A2(new_n682), .ZN(G1330gat));
  NOR3_X1   g482(.A1(new_n676), .A2(new_n408), .A3(new_n651), .ZN(new_n684));
  INV_X1    g483(.A(G50gat), .ZN(new_n685));
  OAI21_X1  g484(.A(KEYINPUT103), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n655), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n655), .A2(new_n687), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n688), .A2(new_n685), .A3(new_n642), .A4(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(new_n684), .B2(new_n685), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n686), .A2(new_n691), .A3(KEYINPUT48), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT48), .ZN(new_n693));
  OAI221_X1 g492(.A(new_n690), .B1(KEYINPUT103), .B2(new_n693), .C1(new_n684), .C2(new_n685), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n692), .A2(new_n694), .ZN(G1331gat));
  AOI21_X1  g494(.A(new_n652), .B1(new_n428), .B2(new_n456), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n576), .A2(new_n625), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n354), .B(KEYINPUT104), .Z(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(G57gat), .ZN(G1332gat));
  INV_X1    g501(.A(KEYINPUT49), .ZN(new_n703));
  INV_X1    g502(.A(G64gat), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n443), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT105), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n699), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n703), .A2(new_n704), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1333gat));
  OAI21_X1  g508(.A(G71gat), .B1(new_n698), .B2(new_n677), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n665), .A2(G71gat), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n710), .B1(new_n698), .B2(new_n711), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n712), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g512(.A1(new_n699), .A2(new_n642), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g514(.A1(new_n570), .A2(new_n624), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n674), .A2(new_n602), .A3(new_n675), .A4(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(G85gat), .B1(new_n717), .B2(new_n354), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n647), .A2(new_n716), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n719), .A2(KEYINPUT51), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(KEYINPUT51), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(new_n602), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n446), .A2(new_n470), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n718), .B1(new_n722), .B2(new_n723), .ZN(G1336gat));
  OAI21_X1  g523(.A(G92gat), .B1(new_n717), .B2(new_n420), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(KEYINPUT51), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n719), .B(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n651), .A2(new_n471), .A3(new_n443), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n730), .B(KEYINPUT106), .Z(new_n731));
  OAI21_X1  g530(.A(new_n725), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(KEYINPUT52), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT108), .ZN(new_n734));
  INV_X1    g533(.A(new_n730), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n720), .A2(new_n721), .A3(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT109), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT52), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n738), .B(new_n725), .C1(new_n736), .C2(new_n737), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT108), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n732), .A2(new_n740), .A3(KEYINPUT52), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n734), .A2(new_n739), .A3(new_n741), .ZN(G1337gat));
  OAI21_X1  g541(.A(G99gat), .B1(new_n717), .B2(new_n677), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n426), .A2(new_n281), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n722), .B2(new_n744), .ZN(G1338gat));
  OAI21_X1  g544(.A(G106gat), .B1(new_n717), .B2(new_n408), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n652), .A2(G106gat), .A3(new_n408), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n746), .B1(new_n729), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT53), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT53), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n746), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n720), .A2(new_n721), .A3(new_n747), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT110), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AND4_X1   g553(.A1(KEYINPUT110), .A2(new_n746), .A3(new_n751), .A4(new_n753), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n750), .B1(new_n754), .B2(new_n755), .ZN(G1339gat));
  AND4_X1   g555(.A1(new_n625), .A2(new_n569), .A3(new_n575), .A4(new_n601), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n605), .B1(new_n603), .B2(new_n604), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n610), .A2(new_n611), .A3(new_n609), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n619), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n623), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n761), .A2(new_n598), .A3(new_n600), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(KEYINPUT113), .ZN(new_n763));
  XNOR2_X1  g562(.A(KEYINPUT111), .B(KEYINPUT54), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n596), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n582), .A2(new_n595), .A3(new_n583), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(KEYINPUT54), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n582), .A2(new_n583), .B1(G230gat), .B2(G233gat), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n765), .B(new_n591), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n586), .A2(KEYINPUT54), .A3(new_n766), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n772), .A2(KEYINPUT55), .A3(new_n591), .A4(new_n765), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n771), .A2(new_n624), .A3(new_n593), .A4(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n761), .A2(new_n598), .A3(new_n775), .A4(new_n600), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n763), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n574), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n572), .A2(new_n773), .A3(new_n593), .A4(new_n573), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n623), .A2(new_n760), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n780), .B1(new_n769), .B2(new_n770), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT112), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n773), .A2(new_n593), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT112), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n785), .A2(new_n513), .A3(new_n786), .A4(new_n781), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n778), .A2(new_n783), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n757), .B1(new_n788), .B2(new_n568), .ZN(new_n789));
  OAI21_X1  g588(.A(KEYINPUT114), .B1(new_n789), .B2(new_n642), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n354), .A2(new_n443), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n783), .A2(new_n787), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n570), .B1(new_n793), .B2(new_n778), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n792), .B(new_n408), .C1(new_n794), .C2(new_n757), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n790), .A2(new_n426), .A3(new_n791), .A4(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(G113gat), .B1(new_n796), .B2(new_n625), .ZN(new_n797));
  INV_X1    g596(.A(new_n789), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n798), .A2(new_n420), .A3(new_n700), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n429), .A2(new_n642), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n624), .A2(new_n243), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n797), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  XOR2_X1   g602(.A(new_n803), .B(KEYINPUT115), .Z(G1340gat));
  OAI21_X1  g603(.A(G120gat), .B1(new_n796), .B2(new_n652), .ZN(new_n805));
  OR2_X1    g604(.A1(new_n601), .A2(new_n242), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n801), .B2(new_n806), .ZN(G1341gat));
  INV_X1    g606(.A(G127gat), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n796), .A2(new_n808), .A3(new_n568), .ZN(new_n809));
  INV_X1    g608(.A(new_n801), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n570), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n809), .B1(new_n808), .B2(new_n811), .ZN(G1342gat));
  NOR3_X1   g611(.A1(new_n801), .A2(G134gat), .A3(new_n574), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT56), .ZN(new_n814));
  OR2_X1    g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n814), .ZN(new_n816));
  OAI21_X1  g615(.A(G134gat), .B1(new_n796), .B2(new_n574), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(G1343gat));
  OR2_X1    g617(.A1(new_n769), .A2(KEYINPUT116), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT55), .B1(new_n769), .B2(KEYINPUT116), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n784), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT117), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n624), .B1(new_n821), .B2(KEYINPUT117), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n762), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n574), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n793), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n757), .B1(new_n827), .B2(new_n568), .ZN(new_n828));
  OAI21_X1  g627(.A(KEYINPUT57), .B1(new_n828), .B2(new_n408), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n798), .A2(new_n830), .A3(new_n642), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n639), .A2(new_n354), .A3(new_n443), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n829), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(G141gat), .B1(new_n833), .B2(new_n625), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n639), .A2(new_n408), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n799), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n837), .A2(new_n306), .A3(new_n624), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n819), .A2(new_n820), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n842), .B1(new_n843), .B2(new_n784), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n844), .A2(new_n624), .A3(new_n822), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n513), .B1(new_n845), .B2(new_n762), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n779), .A2(new_n782), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n568), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n757), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n408), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n841), .B1(new_n850), .B2(KEYINPUT57), .ZN(new_n851));
  INV_X1    g650(.A(new_n847), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n570), .B1(new_n826), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n642), .B1(new_n853), .B2(new_n757), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(KEYINPUT118), .A3(new_n830), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n789), .A2(new_n830), .A3(new_n408), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n859), .A2(KEYINPUT59), .A3(new_n602), .A4(new_n832), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n833), .A2(new_n601), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n860), .B1(KEYINPUT59), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(G148gat), .B1(new_n837), .B2(new_n602), .ZN(new_n863));
  AOI22_X1  g662(.A1(new_n862), .A2(G148gat), .B1(new_n863), .B2(KEYINPUT59), .ZN(G1345gat));
  NOR3_X1   g663(.A1(new_n833), .A2(new_n310), .A3(new_n568), .ZN(new_n865));
  AOI21_X1  g664(.A(G155gat), .B1(new_n837), .B2(new_n570), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(G1346gat));
  NOR3_X1   g666(.A1(new_n833), .A2(new_n311), .A3(new_n574), .ZN(new_n868));
  AOI21_X1  g667(.A(G162gat), .B1(new_n837), .B2(new_n513), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n868), .A2(new_n869), .ZN(G1347gat));
  NOR2_X1   g669(.A1(new_n700), .A2(new_n420), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n790), .A2(new_n795), .A3(new_n426), .A4(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(G169gat), .B1(new_n872), .B2(new_n625), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n789), .A2(new_n446), .A3(new_n420), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n625), .A2(G169gat), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n800), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n873), .A2(new_n876), .ZN(G1348gat));
  AND3_X1   g676(.A1(new_n874), .A2(new_n602), .A3(new_n800), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n651), .A2(G176gat), .ZN(new_n879));
  OAI22_X1  g678(.A1(new_n878), .A2(G176gat), .B1(new_n872), .B2(new_n879), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT119), .ZN(G1349gat));
  NOR2_X1   g680(.A1(KEYINPUT120), .A2(KEYINPUT60), .ZN(new_n882));
  OAI21_X1  g681(.A(G183gat), .B1(new_n872), .B2(new_n568), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n874), .A2(new_n570), .A3(new_n231), .A4(new_n800), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(KEYINPUT120), .A2(KEYINPUT60), .ZN(new_n886));
  XOR2_X1   g685(.A(new_n885), .B(new_n886), .Z(G1350gat));
  OAI21_X1  g686(.A(G190gat), .B1(new_n872), .B2(new_n574), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g689(.A(KEYINPUT121), .B(G190gat), .C1(new_n872), .C2(new_n574), .ZN(new_n891));
  NAND2_X1  g690(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NOR2_X1   g692(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n874), .A2(new_n214), .A3(new_n513), .A4(new_n800), .ZN(new_n896));
  INV_X1    g695(.A(new_n894), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n890), .A2(new_n891), .A3(new_n892), .A4(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n895), .A2(KEYINPUT123), .A3(new_n896), .A4(new_n898), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1351gat));
  NAND2_X1  g702(.A1(new_n677), .A2(new_n871), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT126), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n859), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(G197gat), .B1(new_n906), .B2(new_n625), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n835), .A2(new_n443), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n908), .A2(KEYINPUT124), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n789), .A2(new_n446), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(KEYINPUT124), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n912), .A2(G197gat), .A3(new_n625), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT125), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n907), .A2(new_n914), .ZN(G1352gat));
  OAI21_X1  g714(.A(G204gat), .B1(new_n906), .B2(new_n652), .ZN(new_n916));
  OR3_X1    g715(.A1(new_n912), .A2(G204gat), .A3(new_n601), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(KEYINPUT62), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n917), .A2(KEYINPUT62), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n916), .A2(new_n918), .A3(new_n919), .ZN(G1353gat));
  OR3_X1    g719(.A1(new_n912), .A2(G211gat), .A3(new_n568), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n859), .A2(new_n570), .A3(new_n677), .A4(new_n871), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n922), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT63), .B1(new_n922), .B2(G211gat), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(G1354gat));
  NAND3_X1  g724(.A1(new_n859), .A2(new_n905), .A3(KEYINPUT127), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n857), .B1(new_n851), .B2(new_n855), .ZN(new_n928));
  INV_X1    g727(.A(new_n905), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n926), .A2(new_n513), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(G218gat), .ZN(new_n932));
  OR3_X1    g731(.A1(new_n912), .A2(G218gat), .A3(new_n574), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1355gat));
endmodule


