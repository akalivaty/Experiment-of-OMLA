

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761;

  NOR2_X1 U376 ( .A1(n598), .A2(n597), .ZN(n683) );
  NOR2_X1 U377 ( .A1(G953), .A2(G237), .ZN(n492) );
  NOR2_X1 U378 ( .A1(n596), .A2(n578), .ZN(n672) );
  AND2_X4 U379 ( .A1(n374), .A2(n634), .ZN(n725) );
  NOR2_X2 U380 ( .A1(n601), .A2(KEYINPUT44), .ZN(n602) );
  XNOR2_X1 U381 ( .A(n390), .B(KEYINPUT35), .ZN(n586) );
  NOR2_X1 U382 ( .A1(n588), .A2(n580), .ZN(n581) );
  NAND2_X1 U383 ( .A1(n382), .A2(n380), .ZN(n410) );
  AND2_X1 U384 ( .A1(n386), .A2(n383), .ZN(n382) );
  NOR2_X1 U385 ( .A1(n611), .A2(KEYINPUT83), .ZN(n606) );
  XNOR2_X1 U386 ( .A(n375), .B(n589), .ZN(n698) );
  NOR2_X2 U387 ( .A1(n530), .A2(n529), .ZN(n693) );
  OR2_X1 U388 ( .A1(n583), .A2(n656), .ZN(n375) );
  XOR2_X1 U389 ( .A(n709), .B(n708), .Z(n710) );
  NAND2_X1 U390 ( .A1(n394), .A2(n391), .ZN(n535) );
  AND2_X1 U391 ( .A1(n396), .A2(n395), .ZN(n394) );
  XOR2_X1 U392 ( .A(n717), .B(n716), .Z(n718) );
  INV_X1 U393 ( .A(n625), .ZN(n353) );
  NAND2_X1 U394 ( .A1(n376), .A2(n362), .ZN(n747) );
  XNOR2_X1 U395 ( .A(n354), .B(KEYINPUT84), .ZN(n388) );
  NAND2_X1 U396 ( .A1(n635), .A2(n634), .ZN(n354) );
  INV_X1 U397 ( .A(G128), .ZN(n420) );
  NAND2_X1 U398 ( .A1(n401), .A2(n693), .ZN(n542) );
  XNOR2_X1 U399 ( .A(n402), .B(KEYINPUT77), .ZN(n401) );
  NAND2_X1 U400 ( .A1(n593), .A2(n363), .ZN(n402) );
  AND2_X1 U401 ( .A1(n600), .A2(n413), .ZN(n412) );
  XNOR2_X1 U402 ( .A(G902), .B(KEYINPUT15), .ZN(n610) );
  XNOR2_X1 U403 ( .A(n400), .B(G140), .ZN(n476) );
  XNOR2_X1 U404 ( .A(G125), .B(KEYINPUT10), .ZN(n400) );
  XNOR2_X1 U405 ( .A(n423), .B(G953), .ZN(n447) );
  INV_X1 U406 ( .A(KEYINPUT64), .ZN(n423) );
  XOR2_X1 U407 ( .A(G137), .B(KEYINPUT71), .Z(n505) );
  XNOR2_X1 U408 ( .A(KEYINPUT74), .B(G110), .ZN(n421) );
  NAND2_X1 U409 ( .A1(n435), .A2(G214), .ZN(n637) );
  NAND2_X1 U410 ( .A1(n393), .A2(n392), .ZN(n391) );
  NOR2_X1 U411 ( .A1(n355), .A2(G902), .ZN(n392) );
  XNOR2_X1 U412 ( .A(n509), .B(G469), .ZN(n549) );
  XNOR2_X1 U413 ( .A(n481), .B(n480), .ZN(n648) );
  NOR2_X1 U414 ( .A1(n726), .A2(G902), .ZN(n481) );
  XNOR2_X1 U415 ( .A(G128), .B(G146), .ZN(n470) );
  XOR2_X1 U416 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n472) );
  XOR2_X1 U417 ( .A(G113), .B(G104), .Z(n441) );
  XNOR2_X1 U418 ( .A(n476), .B(n398), .ZN(n438) );
  XNOR2_X1 U419 ( .A(n436), .B(n399), .ZN(n398) );
  XNOR2_X1 U420 ( .A(KEYINPUT100), .B(KEYINPUT101), .ZN(n436) );
  XNOR2_X1 U421 ( .A(KEYINPUT99), .B(KEYINPUT11), .ZN(n399) );
  XNOR2_X1 U422 ( .A(G131), .B(G143), .ZN(n439) );
  XNOR2_X1 U423 ( .A(n487), .B(n486), .ZN(n745) );
  INV_X1 U424 ( .A(n418), .ZN(n385) );
  BUF_X1 U425 ( .A(n550), .Z(n407) );
  AND2_X1 U426 ( .A1(n407), .A2(n482), .ZN(n573) );
  BUF_X1 U427 ( .A(n648), .Z(n408) );
  INV_X1 U428 ( .A(n407), .ZN(n409) );
  NOR2_X1 U429 ( .A1(n407), .A2(n360), .ZN(n646) );
  XNOR2_X1 U430 ( .A(n525), .B(n403), .ZN(n593) );
  INV_X1 U431 ( .A(KEYINPUT103), .ZN(n403) );
  OR2_X1 U432 ( .A1(n699), .A2(n696), .ZN(n525) );
  NAND2_X1 U433 ( .A1(n355), .A2(G902), .ZN(n395) );
  XNOR2_X1 U434 ( .A(G113), .B(G137), .ZN(n489) );
  XOR2_X1 U435 ( .A(KEYINPUT5), .B(KEYINPUT97), .Z(n495) );
  NOR2_X1 U436 ( .A1(n552), .A2(n702), .ZN(n553) );
  XNOR2_X1 U437 ( .A(KEYINPUT3), .B(G119), .ZN(n427) );
  XOR2_X1 U438 ( .A(G107), .B(G122), .Z(n450) );
  XNOR2_X1 U439 ( .A(n747), .B(KEYINPUT80), .ZN(n611) );
  XNOR2_X1 U440 ( .A(KEYINPUT18), .B(KEYINPUT81), .ZN(n378) );
  AND2_X1 U441 ( .A1(n748), .A2(G224), .ZN(n426) );
  XNOR2_X1 U442 ( .A(G125), .B(KEYINPUT17), .ZN(n424) );
  XNOR2_X1 U443 ( .A(n549), .B(n364), .ZN(n550) );
  XNOR2_X1 U444 ( .A(n431), .B(KEYINPUT94), .ZN(n432) );
  OR2_X1 U445 ( .A1(n652), .A2(n514), .ZN(n516) );
  AND2_X1 U446 ( .A1(n648), .A2(n649), .ZN(n360) );
  NOR2_X1 U447 ( .A1(n747), .A2(n627), .ZN(n616) );
  OR2_X1 U448 ( .A1(n532), .A2(n519), .ZN(n520) );
  NOR2_X1 U449 ( .A1(n547), .A2(n652), .ZN(n500) );
  XNOR2_X1 U450 ( .A(n535), .B(KEYINPUT102), .ZN(n524) );
  NAND2_X1 U451 ( .A1(n360), .A2(n549), .ZN(n590) );
  XNOR2_X1 U452 ( .A(n475), .B(n474), .ZN(n477) );
  XNOR2_X1 U453 ( .A(n444), .B(n443), .ZN(n717) );
  XNOR2_X1 U454 ( .A(n358), .B(n442), .ZN(n443) );
  XNOR2_X1 U455 ( .A(n508), .B(n507), .ZN(n620) );
  AND2_X1 U456 ( .A1(n384), .A2(n731), .ZN(n383) );
  NAND2_X1 U457 ( .A1(n385), .A2(KEYINPUT116), .ZN(n384) );
  NAND2_X1 U458 ( .A1(n381), .A2(KEYINPUT116), .ZN(n380) );
  INV_X1 U459 ( .A(n585), .ZN(n406) );
  AND2_X1 U460 ( .A1(n580), .A2(n573), .ZN(n419) );
  NAND2_X1 U461 ( .A1(n577), .A2(n409), .ZN(n578) );
  AND2_X1 U462 ( .A1(n524), .A2(n533), .ZN(n696) );
  NAND2_X1 U463 ( .A1(n409), .A2(n408), .ZN(n597) );
  XOR2_X1 U464 ( .A(n446), .B(n445), .Z(n355) );
  AND2_X1 U465 ( .A1(n725), .A2(G478), .ZN(n356) );
  NOR2_X1 U466 ( .A1(n583), .A2(n592), .ZN(n357) );
  XOR2_X1 U467 ( .A(n440), .B(n439), .Z(n358) );
  OR2_X1 U468 ( .A1(G237), .A2(G902), .ZN(n359) );
  XNOR2_X1 U469 ( .A(n581), .B(n416), .ZN(n636) );
  AND2_X1 U470 ( .A1(n568), .A2(n567), .ZN(n361) );
  AND2_X1 U471 ( .A1(n759), .A2(n670), .ZN(n362) );
  XOR2_X1 U472 ( .A(KEYINPUT70), .B(KEYINPUT47), .Z(n363) );
  XOR2_X1 U473 ( .A(KEYINPUT1), .B(KEYINPUT67), .Z(n364) );
  XNOR2_X1 U474 ( .A(KEYINPUT76), .B(KEYINPUT34), .ZN(n365) );
  XOR2_X1 U475 ( .A(n555), .B(KEYINPUT72), .Z(n366) );
  INV_X1 U476 ( .A(G953), .ZN(n731) );
  XOR2_X1 U477 ( .A(n669), .B(KEYINPUT53), .Z(n367) );
  INV_X1 U478 ( .A(KEYINPUT116), .ZN(n411) );
  NOR2_X1 U479 ( .A1(n582), .A2(n572), .ZN(n368) );
  XNOR2_X1 U480 ( .A(n368), .B(KEYINPUT22), .ZN(n574) );
  XNOR2_X1 U481 ( .A(n404), .B(n575), .ZN(n674) );
  XNOR2_X1 U482 ( .A(n369), .B(n370), .ZN(n680) );
  NAND2_X1 U483 ( .A1(n725), .A2(G472), .ZN(n369) );
  XOR2_X1 U484 ( .A(n678), .B(n677), .Z(n370) );
  NAND2_X1 U485 ( .A1(n707), .A2(n610), .ZN(n433) );
  XNOR2_X1 U486 ( .A(n371), .B(n737), .ZN(n707) );
  XNOR2_X1 U487 ( .A(n372), .B(n373), .ZN(n371) );
  XNOR2_X1 U488 ( .A(n422), .B(n426), .ZN(n372) );
  XNOR2_X1 U489 ( .A(n504), .B(n425), .ZN(n373) );
  NAND2_X1 U490 ( .A1(n614), .A2(n615), .ZN(n374) );
  XNOR2_X1 U491 ( .A(n556), .B(n366), .ZN(n376) );
  XNOR2_X2 U492 ( .A(n433), .B(n432), .ZN(n526) );
  BUF_X1 U493 ( .A(n447), .Z(n748) );
  NOR2_X2 U494 ( .A1(n712), .A2(n730), .ZN(n713) );
  NOR2_X2 U495 ( .A1(n720), .A2(n730), .ZN(n721) );
  NOR2_X2 U496 ( .A1(n623), .A2(n730), .ZN(n624) );
  XNOR2_X1 U497 ( .A(n405), .B(n377), .ZN(n422) );
  XNOR2_X1 U498 ( .A(n485), .B(n378), .ZN(n377) );
  XNOR2_X2 U499 ( .A(KEYINPUT4), .B(G146), .ZN(n485) );
  XNOR2_X2 U500 ( .A(n379), .B(n420), .ZN(n405) );
  XNOR2_X2 U501 ( .A(KEYINPUT65), .B(G143), .ZN(n379) );
  INV_X1 U502 ( .A(n388), .ZN(n381) );
  NAND2_X1 U503 ( .A1(n388), .A2(n387), .ZN(n386) );
  AND2_X1 U504 ( .A1(n418), .A2(n411), .ZN(n387) );
  NAND2_X1 U505 ( .A1(n389), .A2(n406), .ZN(n390) );
  XNOR2_X1 U506 ( .A(n584), .B(n365), .ZN(n389) );
  INV_X1 U507 ( .A(n586), .ZN(n760) );
  INV_X1 U508 ( .A(n717), .ZN(n393) );
  NAND2_X1 U509 ( .A1(n717), .A2(n355), .ZN(n396) );
  INV_X1 U510 ( .A(G902), .ZN(n397) );
  NAND2_X1 U511 ( .A1(n574), .A2(n419), .ZN(n404) );
  XNOR2_X1 U512 ( .A(n405), .B(G134), .ZN(n487) );
  XNOR2_X1 U513 ( .A(n570), .B(KEYINPUT0), .ZN(n582) );
  XNOR2_X1 U514 ( .A(n415), .B(KEYINPUT88), .ZN(n603) );
  NOR2_X2 U515 ( .A1(n674), .A2(n672), .ZN(n579) );
  NAND2_X1 U516 ( .A1(n587), .A2(KEYINPUT44), .ZN(n414) );
  XNOR2_X1 U517 ( .A(n473), .B(n472), .ZN(n474) );
  NAND2_X1 U518 ( .A1(n550), .A2(n360), .ZN(n588) );
  NAND2_X1 U519 ( .A1(n557), .A2(n409), .ZN(n558) );
  INV_X1 U520 ( .A(n574), .ZN(n596) );
  XNOR2_X1 U521 ( .A(n410), .B(n367), .ZN(G75) );
  NAND2_X1 U522 ( .A1(n414), .A2(n412), .ZN(n415) );
  NAND2_X1 U523 ( .A1(n586), .A2(KEYINPUT44), .ZN(n413) );
  OR2_X1 U524 ( .A1(n587), .A2(n586), .ZN(n601) );
  BUF_X2 U525 ( .A(n626), .Z(n732) );
  XOR2_X1 U526 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n416) );
  XOR2_X1 U527 ( .A(n503), .B(n502), .Z(n417) );
  AND2_X1 U528 ( .A1(n668), .A2(n667), .ZN(n418) );
  XNOR2_X1 U529 ( .A(n501), .B(G104), .ZN(n503) );
  NOR2_X1 U530 ( .A1(n636), .A2(n583), .ZN(n584) );
  OR2_X1 U531 ( .A1(n748), .A2(G952), .ZN(n679) );
  BUF_X1 U532 ( .A(n674), .Z(n675) );
  XNOR2_X1 U533 ( .A(KEYINPUT69), .B(G101), .ZN(n488) );
  XNOR2_X1 U534 ( .A(n488), .B(n421), .ZN(n504) );
  XNOR2_X1 U535 ( .A(n424), .B(KEYINPUT93), .ZN(n425) );
  XNOR2_X1 U536 ( .A(n441), .B(n450), .ZN(n430) );
  XNOR2_X1 U537 ( .A(n427), .B(G116), .ZN(n490) );
  INV_X1 U538 ( .A(KEYINPUT16), .ZN(n428) );
  XNOR2_X1 U539 ( .A(n490), .B(n428), .ZN(n429) );
  XNOR2_X1 U540 ( .A(n430), .B(n429), .ZN(n737) );
  XNOR2_X1 U541 ( .A(KEYINPUT78), .B(n359), .ZN(n435) );
  AND2_X1 U542 ( .A1(n435), .A2(G210), .ZN(n431) );
  BUF_X1 U543 ( .A(n526), .Z(n434) );
  XNOR2_X1 U544 ( .A(n434), .B(KEYINPUT38), .ZN(n519) );
  INV_X1 U545 ( .A(n519), .ZN(n638) );
  NAND2_X1 U546 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U547 ( .A1(G214), .A2(n492), .ZN(n437) );
  XNOR2_X1 U548 ( .A(n438), .B(n437), .ZN(n444) );
  XOR2_X1 U549 ( .A(KEYINPUT12), .B(G122), .Z(n440) );
  XNOR2_X1 U550 ( .A(G146), .B(n441), .ZN(n442) );
  INV_X1 U551 ( .A(G475), .ZN(n446) );
  INV_X1 U552 ( .A(KEYINPUT13), .ZN(n445) );
  INV_X1 U553 ( .A(n535), .ZN(n458) );
  INV_X1 U554 ( .A(KEYINPUT8), .ZN(n449) );
  NAND2_X1 U555 ( .A1(G234), .A2(n447), .ZN(n448) );
  XNOR2_X1 U556 ( .A(n449), .B(n448), .ZN(n469) );
  NAND2_X1 U557 ( .A1(n469), .A2(G217), .ZN(n454) );
  XOR2_X1 U558 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n452) );
  XNOR2_X1 U559 ( .A(G116), .B(n450), .ZN(n451) );
  XNOR2_X1 U560 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U561 ( .A(n454), .B(n453), .ZN(n456) );
  INV_X1 U562 ( .A(n487), .ZN(n455) );
  XNOR2_X1 U563 ( .A(n456), .B(n455), .ZN(n723) );
  NAND2_X1 U564 ( .A1(n723), .A2(n397), .ZN(n457) );
  INV_X1 U565 ( .A(G478), .ZN(n722) );
  XNOR2_X1 U566 ( .A(n457), .B(n722), .ZN(n533) );
  NAND2_X1 U567 ( .A1(n458), .A2(n533), .ZN(n639) );
  NOR2_X1 U568 ( .A1(n641), .A2(n639), .ZN(n459) );
  XNOR2_X1 U569 ( .A(KEYINPUT41), .B(n459), .ZN(n660) );
  NAND2_X1 U570 ( .A1(n610), .A2(G234), .ZN(n460) );
  XNOR2_X1 U571 ( .A(n460), .B(KEYINPUT96), .ZN(n461) );
  XNOR2_X1 U572 ( .A(KEYINPUT20), .B(n461), .ZN(n478) );
  AND2_X1 U573 ( .A1(n478), .A2(G221), .ZN(n462) );
  XNOR2_X1 U574 ( .A(n462), .B(KEYINPUT21), .ZN(n649) );
  INV_X1 U575 ( .A(n649), .ZN(n468) );
  NOR2_X1 U576 ( .A1(G900), .A2(n748), .ZN(n463) );
  NAND2_X1 U577 ( .A1(G902), .A2(n463), .ZN(n464) );
  NAND2_X1 U578 ( .A1(n731), .A2(G952), .ZN(n565) );
  NAND2_X1 U579 ( .A1(n464), .A2(n565), .ZN(n467) );
  NAND2_X1 U580 ( .A1(G237), .A2(G234), .ZN(n466) );
  INV_X1 U581 ( .A(KEYINPUT14), .ZN(n465) );
  XNOR2_X1 U582 ( .A(n466), .B(n465), .ZN(n665) );
  INV_X1 U583 ( .A(n665), .ZN(n567) );
  NAND2_X1 U584 ( .A1(n467), .A2(n567), .ZN(n513) );
  NOR2_X1 U585 ( .A1(n468), .A2(n513), .ZN(n483) );
  NAND2_X1 U586 ( .A1(G221), .A2(n469), .ZN(n475) );
  XOR2_X1 U587 ( .A(G110), .B(G119), .Z(n471) );
  XNOR2_X1 U588 ( .A(n471), .B(n470), .ZN(n473) );
  XNOR2_X1 U589 ( .A(n476), .B(n505), .ZN(n746) );
  XNOR2_X1 U590 ( .A(n477), .B(n746), .ZN(n726) );
  NAND2_X1 U591 ( .A1(n478), .A2(G217), .ZN(n479) );
  XNOR2_X1 U592 ( .A(KEYINPUT25), .B(n479), .ZN(n480) );
  INV_X1 U593 ( .A(n648), .ZN(n482) );
  NAND2_X1 U594 ( .A1(n483), .A2(n482), .ZN(n484) );
  XOR2_X1 U595 ( .A(KEYINPUT73), .B(n484), .Z(n547) );
  XNOR2_X1 U596 ( .A(n485), .B(G131), .ZN(n486) );
  XNOR2_X1 U597 ( .A(n489), .B(n488), .ZN(n491) );
  XNOR2_X1 U598 ( .A(n491), .B(n490), .ZN(n497) );
  NAND2_X1 U599 ( .A1(n492), .A2(G210), .ZN(n493) );
  XNOR2_X1 U600 ( .A(n493), .B(KEYINPUT79), .ZN(n494) );
  XNOR2_X1 U601 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U602 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U603 ( .A(n745), .B(n498), .ZN(n678) );
  OR2_X1 U604 ( .A1(n678), .A2(G902), .ZN(n499) );
  INV_X1 U605 ( .A(G472), .ZN(n676) );
  XNOR2_X2 U606 ( .A(n499), .B(n676), .ZN(n652) );
  XNOR2_X1 U607 ( .A(n500), .B(KEYINPUT28), .ZN(n510) );
  INV_X1 U608 ( .A(n745), .ZN(n508) );
  XOR2_X1 U609 ( .A(G107), .B(G140), .Z(n501) );
  NAND2_X1 U610 ( .A1(G227), .A2(n447), .ZN(n502) );
  XNOR2_X1 U611 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U612 ( .A(n417), .B(n506), .ZN(n507) );
  NAND2_X1 U613 ( .A1(n620), .A2(n397), .ZN(n509) );
  NAND2_X1 U614 ( .A1(n510), .A2(n549), .ZN(n530) );
  NOR2_X1 U615 ( .A1(n660), .A2(n530), .ZN(n512) );
  INV_X1 U616 ( .A(KEYINPUT42), .ZN(n511) );
  XNOR2_X1 U617 ( .A(n512), .B(n511), .ZN(n761) );
  NOR2_X1 U618 ( .A1(n590), .A2(n513), .ZN(n518) );
  INV_X1 U619 ( .A(n637), .ZN(n514) );
  INV_X1 U620 ( .A(KEYINPUT30), .ZN(n515) );
  XNOR2_X1 U621 ( .A(n516), .B(n515), .ZN(n517) );
  NAND2_X1 U622 ( .A1(n518), .A2(n517), .ZN(n532) );
  XNOR2_X2 U623 ( .A(n520), .B(KEYINPUT39), .ZN(n562) );
  NAND2_X1 U624 ( .A1(n562), .A2(n696), .ZN(n521) );
  XNOR2_X1 U625 ( .A(n521), .B(KEYINPUT40), .ZN(n671) );
  NAND2_X1 U626 ( .A1(n761), .A2(n671), .ZN(n523) );
  XNOR2_X1 U627 ( .A(KEYINPUT87), .B(KEYINPUT46), .ZN(n522) );
  XNOR2_X1 U628 ( .A(n523), .B(n522), .ZN(n554) );
  NOR2_X1 U629 ( .A1(n524), .A2(n533), .ZN(n699) );
  NAND2_X1 U630 ( .A1(n526), .A2(n637), .ZN(n528) );
  INV_X1 U631 ( .A(KEYINPUT19), .ZN(n527) );
  XNOR2_X1 U632 ( .A(n528), .B(n527), .ZN(n563) );
  BUF_X1 U633 ( .A(n563), .Z(n529) );
  NAND2_X1 U634 ( .A1(n693), .A2(n593), .ZN(n531) );
  NAND2_X1 U635 ( .A1(n531), .A2(KEYINPUT47), .ZN(n540) );
  INV_X1 U636 ( .A(n532), .ZN(n538) );
  INV_X1 U637 ( .A(n533), .ZN(n534) );
  NAND2_X1 U638 ( .A1(n535), .A2(n534), .ZN(n585) );
  INV_X1 U639 ( .A(n434), .ZN(n536) );
  NOR2_X1 U640 ( .A1(n585), .A2(n536), .ZN(n537) );
  AND2_X1 U641 ( .A1(n538), .A2(n537), .ZN(n692) );
  INV_X1 U642 ( .A(n692), .ZN(n539) );
  AND2_X1 U643 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U644 ( .A1(n542), .A2(n541), .ZN(n552) );
  INV_X1 U645 ( .A(n696), .ZN(n544) );
  INV_X1 U646 ( .A(KEYINPUT6), .ZN(n543) );
  XNOR2_X1 U647 ( .A(n652), .B(n543), .ZN(n580) );
  NOR2_X1 U648 ( .A1(n544), .A2(n580), .ZN(n545) );
  NAND2_X1 U649 ( .A1(n545), .A2(n637), .ZN(n546) );
  NOR2_X1 U650 ( .A1(n547), .A2(n546), .ZN(n557) );
  AND2_X1 U651 ( .A1(n434), .A2(n557), .ZN(n548) );
  XNOR2_X1 U652 ( .A(n548), .B(KEYINPUT36), .ZN(n551) );
  AND2_X1 U653 ( .A1(n551), .A2(n407), .ZN(n702) );
  NAND2_X1 U654 ( .A1(n554), .A2(n553), .ZN(n556) );
  XNOR2_X1 U655 ( .A(KEYINPUT86), .B(KEYINPUT48), .ZN(n555) );
  XNOR2_X1 U656 ( .A(KEYINPUT104), .B(KEYINPUT43), .ZN(n559) );
  XOR2_X1 U657 ( .A(n559), .B(n558), .Z(n560) );
  NOR2_X1 U658 ( .A1(n560), .A2(n434), .ZN(n561) );
  XNOR2_X1 U659 ( .A(n561), .B(KEYINPUT105), .ZN(n759) );
  NAND2_X1 U660 ( .A1(n562), .A2(n699), .ZN(n670) );
  INV_X1 U661 ( .A(n563), .ZN(n569) );
  NOR2_X1 U662 ( .A1(G898), .A2(n731), .ZN(n564) );
  XOR2_X1 U663 ( .A(KEYINPUT95), .B(n564), .Z(n741) );
  NAND2_X1 U664 ( .A1(n741), .A2(G902), .ZN(n566) );
  NAND2_X1 U665 ( .A1(n566), .A2(n565), .ZN(n568) );
  NAND2_X1 U666 ( .A1(n569), .A2(n361), .ZN(n570) );
  INV_X1 U667 ( .A(n639), .ZN(n571) );
  NAND2_X1 U668 ( .A1(n571), .A2(n649), .ZN(n572) );
  INV_X1 U669 ( .A(n580), .ZN(n595) );
  XOR2_X1 U670 ( .A(KEYINPUT66), .B(KEYINPUT32), .Z(n575) );
  INV_X1 U671 ( .A(n652), .ZN(n576) );
  NOR2_X1 U672 ( .A1(n408), .A2(n576), .ZN(n577) );
  XNOR2_X1 U673 ( .A(n579), .B(KEYINPUT89), .ZN(n587) );
  BUF_X1 U674 ( .A(n582), .Z(n583) );
  XNOR2_X1 U675 ( .A(KEYINPUT31), .B(KEYINPUT98), .ZN(n589) );
  OR2_X1 U676 ( .A1(n588), .A2(n652), .ZN(n656) );
  INV_X1 U677 ( .A(n590), .ZN(n591) );
  NAND2_X1 U678 ( .A1(n591), .A2(n652), .ZN(n592) );
  NOR2_X1 U679 ( .A1(n698), .A2(n357), .ZN(n594) );
  INV_X1 U680 ( .A(n593), .ZN(n642) );
  NOR2_X1 U681 ( .A1(n594), .A2(n642), .ZN(n599) );
  OR2_X1 U682 ( .A1(n596), .A2(n595), .ZN(n598) );
  NOR2_X1 U683 ( .A1(n599), .A2(n683), .ZN(n600) );
  NOR2_X2 U684 ( .A1(n603), .A2(n602), .ZN(n605) );
  INV_X1 U685 ( .A(KEYINPUT45), .ZN(n604) );
  XNOR2_X2 U686 ( .A(n605), .B(n604), .ZN(n626) );
  NAND2_X1 U687 ( .A1(n606), .A2(n626), .ZN(n607) );
  INV_X1 U688 ( .A(KEYINPUT2), .ZN(n627) );
  NAND2_X1 U689 ( .A1(n607), .A2(n627), .ZN(n609) );
  INV_X1 U690 ( .A(n610), .ZN(n608) );
  NAND2_X1 U691 ( .A1(n609), .A2(n608), .ZN(n615) );
  NOR2_X1 U692 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U693 ( .A1(n732), .A2(n612), .ZN(n613) );
  NAND2_X1 U694 ( .A1(n613), .A2(KEYINPUT83), .ZN(n614) );
  XOR2_X1 U695 ( .A(KEYINPUT85), .B(n616), .Z(n617) );
  NAND2_X1 U696 ( .A1(n617), .A2(n732), .ZN(n634) );
  NAND2_X1 U697 ( .A1(n725), .A2(G469), .ZN(n622) );
  XNOR2_X1 U698 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n618) );
  XOR2_X1 U699 ( .A(n618), .B(KEYINPUT57), .Z(n619) );
  XNOR2_X1 U700 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U701 ( .A(n622), .B(n621), .ZN(n623) );
  INV_X1 U702 ( .A(n679), .ZN(n730) );
  XNOR2_X1 U703 ( .A(n624), .B(KEYINPUT120), .ZN(G54) );
  INV_X1 U704 ( .A(n747), .ZN(n625) );
  NAND2_X1 U705 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n629), .A2(KEYINPUT82), .ZN(n633) );
  NOR2_X1 U708 ( .A1(KEYINPUT2), .A2(KEYINPUT82), .ZN(n630) );
  AND2_X1 U709 ( .A1(n747), .A2(n630), .ZN(n631) );
  NAND2_X1 U710 ( .A1(n732), .A2(n631), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n633), .A2(n632), .ZN(n635) );
  OR2_X1 U712 ( .A1(n660), .A2(n636), .ZN(n668) );
  NOR2_X1 U713 ( .A1(n638), .A2(n637), .ZN(n640) );
  NOR2_X1 U714 ( .A1(n640), .A2(n639), .ZN(n644) );
  NOR2_X1 U715 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U716 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U717 ( .A1(n636), .A2(n645), .ZN(n662) );
  XNOR2_X1 U718 ( .A(n646), .B(KEYINPUT50), .ZN(n655) );
  XOR2_X1 U719 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n647) );
  XNOR2_X1 U720 ( .A(KEYINPUT114), .B(n647), .ZN(n651) );
  NOR2_X1 U721 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U722 ( .A(n651), .B(n650), .ZN(n653) );
  NAND2_X1 U723 ( .A1(n653), .A2(n652), .ZN(n654) );
  OR2_X1 U724 ( .A1(n655), .A2(n654), .ZN(n657) );
  NAND2_X1 U725 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U726 ( .A(KEYINPUT51), .B(n658), .ZN(n659) );
  NOR2_X1 U727 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U728 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U729 ( .A(n663), .B(KEYINPUT52), .ZN(n664) );
  NOR2_X1 U730 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U731 ( .A1(n666), .A2(G952), .ZN(n667) );
  INV_X1 U732 ( .A(KEYINPUT117), .ZN(n669) );
  XNOR2_X1 U733 ( .A(n670), .B(G134), .ZN(G36) );
  XNOR2_X1 U734 ( .A(n671), .B(G131), .ZN(G33) );
  XOR2_X1 U735 ( .A(G110), .B(KEYINPUT107), .Z(n673) );
  XOR2_X1 U736 ( .A(n673), .B(n672), .Z(G12) );
  XOR2_X1 U737 ( .A(n675), .B(G119), .Z(G21) );
  XOR2_X1 U738 ( .A(KEYINPUT91), .B(KEYINPUT62), .Z(n677) );
  NAND2_X1 U739 ( .A1(n680), .A2(n679), .ZN(n682) );
  XNOR2_X1 U740 ( .A(KEYINPUT106), .B(KEYINPUT63), .ZN(n681) );
  XNOR2_X1 U741 ( .A(n682), .B(n681), .ZN(G57) );
  XOR2_X1 U742 ( .A(G101), .B(n683), .Z(G3) );
  NAND2_X1 U743 ( .A1(n357), .A2(n696), .ZN(n684) );
  XNOR2_X1 U744 ( .A(n684), .B(G104), .ZN(G6) );
  XOR2_X1 U745 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n686) );
  NAND2_X1 U746 ( .A1(n357), .A2(n699), .ZN(n685) );
  XNOR2_X1 U747 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U748 ( .A(G107), .B(n687), .ZN(G9) );
  XOR2_X1 U749 ( .A(KEYINPUT29), .B(KEYINPUT109), .Z(n689) );
  NAND2_X1 U750 ( .A1(n693), .A2(n699), .ZN(n688) );
  XNOR2_X1 U751 ( .A(n689), .B(n688), .ZN(n691) );
  XOR2_X1 U752 ( .A(G128), .B(KEYINPUT108), .Z(n690) );
  XNOR2_X1 U753 ( .A(n691), .B(n690), .ZN(G30) );
  XOR2_X1 U754 ( .A(G143), .B(n692), .Z(G45) );
  NAND2_X1 U755 ( .A1(n693), .A2(n696), .ZN(n694) );
  XNOR2_X1 U756 ( .A(n694), .B(KEYINPUT110), .ZN(n695) );
  XNOR2_X1 U757 ( .A(G146), .B(n695), .ZN(G48) );
  NAND2_X1 U758 ( .A1(n698), .A2(n696), .ZN(n697) );
  XNOR2_X1 U759 ( .A(n697), .B(G113), .ZN(G15) );
  XOR2_X1 U760 ( .A(G116), .B(KEYINPUT111), .Z(n701) );
  NAND2_X1 U761 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U762 ( .A(n701), .B(n700), .ZN(G18) );
  XNOR2_X1 U763 ( .A(n702), .B(KEYINPUT37), .ZN(n703) );
  XNOR2_X1 U764 ( .A(n703), .B(KEYINPUT112), .ZN(n704) );
  XNOR2_X1 U765 ( .A(G125), .B(n704), .ZN(G27) );
  NAND2_X1 U766 ( .A1(n725), .A2(G210), .ZN(n711) );
  XOR2_X1 U767 ( .A(KEYINPUT90), .B(KEYINPUT55), .Z(n706) );
  XNOR2_X1 U768 ( .A(KEYINPUT118), .B(KEYINPUT54), .ZN(n705) );
  XNOR2_X1 U769 ( .A(n706), .B(n705), .ZN(n709) );
  BUF_X1 U770 ( .A(n707), .Z(n708) );
  XNOR2_X1 U771 ( .A(n711), .B(n710), .ZN(n712) );
  XNOR2_X1 U772 ( .A(n713), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U773 ( .A1(n725), .A2(G475), .ZN(n719) );
  XOR2_X1 U774 ( .A(KEYINPUT92), .B(KEYINPUT68), .Z(n715) );
  XNOR2_X1 U775 ( .A(KEYINPUT121), .B(KEYINPUT59), .ZN(n714) );
  XNOR2_X1 U776 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X1 U777 ( .A(n719), .B(n718), .ZN(n720) );
  XNOR2_X1 U778 ( .A(n721), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U779 ( .A(n356), .B(n723), .ZN(n724) );
  NOR2_X1 U780 ( .A1(n730), .A2(n724), .ZN(G63) );
  NAND2_X1 U781 ( .A1(n725), .A2(G217), .ZN(n728) );
  XNOR2_X1 U782 ( .A(n726), .B(KEYINPUT122), .ZN(n727) );
  XNOR2_X1 U783 ( .A(n728), .B(n727), .ZN(n729) );
  NOR2_X1 U784 ( .A1(n730), .A2(n729), .ZN(G66) );
  NAND2_X1 U785 ( .A1(n732), .A2(n731), .ZN(n736) );
  NAND2_X1 U786 ( .A1(G953), .A2(G224), .ZN(n733) );
  XNOR2_X1 U787 ( .A(KEYINPUT61), .B(n733), .ZN(n734) );
  NAND2_X1 U788 ( .A1(n734), .A2(G898), .ZN(n735) );
  NAND2_X1 U789 ( .A1(n736), .A2(n735), .ZN(n743) );
  XNOR2_X1 U790 ( .A(G110), .B(n737), .ZN(n738) );
  XNOR2_X1 U791 ( .A(n738), .B(KEYINPUT123), .ZN(n739) );
  XNOR2_X1 U792 ( .A(n739), .B(G101), .ZN(n740) );
  NOR2_X1 U793 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U794 ( .A(n743), .B(n742), .ZN(n744) );
  XNOR2_X1 U795 ( .A(KEYINPUT124), .B(n744), .ZN(G69) );
  XOR2_X1 U796 ( .A(n746), .B(n745), .Z(n751) );
  XNOR2_X1 U797 ( .A(n353), .B(n751), .ZN(n749) );
  NAND2_X1 U798 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U799 ( .A(KEYINPUT125), .B(n750), .Z(n757) );
  XNOR2_X1 U800 ( .A(n751), .B(G227), .ZN(n752) );
  XNOR2_X1 U801 ( .A(n752), .B(KEYINPUT126), .ZN(n753) );
  NAND2_X1 U802 ( .A1(n753), .A2(G900), .ZN(n754) );
  XOR2_X1 U803 ( .A(KEYINPUT127), .B(n754), .Z(n755) );
  NAND2_X1 U804 ( .A1(G953), .A2(n755), .ZN(n756) );
  NAND2_X1 U805 ( .A1(n757), .A2(n756), .ZN(G72) );
  XOR2_X1 U806 ( .A(G140), .B(KEYINPUT113), .Z(n758) );
  XNOR2_X1 U807 ( .A(n759), .B(n758), .ZN(G42) );
  XNOR2_X1 U808 ( .A(n760), .B(G122), .ZN(G24) );
  XNOR2_X1 U809 ( .A(G137), .B(n761), .ZN(G39) );
endmodule

