//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n568, new_n570, new_n571, new_n572, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1180;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G120), .Z(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT65), .Z(G319));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  AND3_X1   g035(.A1(new_n460), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(KEYINPUT67), .B1(new_n460), .B2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND4_X1  g040(.A1(new_n464), .A2(KEYINPUT68), .A3(G137), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n463), .A2(new_n462), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n460), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n467), .A2(G137), .A3(new_n465), .A4(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n465), .A2(G101), .A3(G2104), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n475));
  INV_X1    g050(.A(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT3), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n462), .A2(new_n477), .A3(G125), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n475), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  AOI211_X1 g056(.A(KEYINPUT66), .B(new_n465), .C1(new_n478), .C2(new_n479), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n474), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT69), .ZN(G160));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n487));
  INV_X1    g062(.A(G124), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n467), .A2(G2105), .A3(new_n468), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n464), .A2(new_n465), .ZN(new_n490));
  INV_X1    g065(.A(G136), .ZN(new_n491));
  OAI221_X1 g066(.A(new_n487), .B1(new_n488), .B2(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n492), .B(new_n493), .ZN(G162));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  AND4_X1   g072(.A1(new_n495), .A2(new_n497), .A3(new_n462), .A4(new_n477), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n467), .A2(G138), .A3(new_n465), .A4(new_n468), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(KEYINPUT4), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n467), .A2(G126), .A3(G2105), .A4(new_n468), .ZN(new_n501));
  OR2_X1    g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n502), .B(G2104), .C1(G114), .C2(new_n465), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n500), .A2(new_n504), .ZN(G164));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT6), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  XOR2_X1   g088(.A(new_n513), .B(KEYINPUT71), .Z(new_n514));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n515));
  OAI21_X1  g090(.A(G543), .B1(new_n515), .B2(KEYINPUT5), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n517), .A2(new_n515), .A3(KEYINPUT5), .A4(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n507), .A2(new_n509), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  OAI221_X1 g100(.A(new_n514), .B1(new_n523), .B2(new_n524), .C1(new_n525), .C2(new_n506), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  INV_X1    g102(.A(KEYINPUT76), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(KEYINPUT75), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(KEYINPUT75), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT7), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n530), .A2(KEYINPUT7), .A3(new_n531), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G89), .ZN(new_n537));
  AOI211_X1 g112(.A(new_n537), .B(new_n510), .C1(new_n519), .C2(new_n520), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n528), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n521), .A2(G89), .A3(new_n522), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n540), .A2(KEYINPUT76), .A3(new_n534), .A4(new_n535), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n522), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G51), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(G63), .ZN(new_n546));
  AOI211_X1 g121(.A(new_n546), .B(new_n506), .C1(new_n519), .C2(new_n520), .ZN(new_n547));
  OAI21_X1  g122(.A(KEYINPUT74), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT74), .ZN(new_n550));
  OAI211_X1 g125(.A(new_n549), .B(new_n550), .C1(new_n544), .C2(new_n543), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n542), .A2(new_n552), .ZN(G286));
  INV_X1    g128(.A(G286), .ZN(G168));
  AOI22_X1  g129(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(new_n506), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n512), .A2(G52), .ZN(new_n557));
  INV_X1    g132(.A(G90), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n523), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n556), .A2(new_n559), .ZN(G171));
  AOI22_X1  g135(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n561), .A2(new_n506), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n512), .A2(G43), .ZN(new_n563));
  INV_X1    g138(.A(G81), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n523), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  AND3_X1   g142(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G36), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT77), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(G188));
  XOR2_X1   g148(.A(KEYINPUT78), .B(KEYINPUT9), .Z(new_n574));
  NAND3_X1  g149(.A1(new_n512), .A2(G53), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(KEYINPUT79), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT79), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n512), .A2(new_n577), .A3(G53), .A4(new_n574), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT9), .ZN(new_n579));
  AND2_X1   g154(.A1(new_n512), .A2(G53), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n576), .B(new_n578), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n523), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G91), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n521), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(new_n506), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n581), .A2(new_n583), .A3(new_n585), .ZN(G299));
  INV_X1    g161(.A(G171), .ZN(G301));
  OR2_X1    g162(.A1(new_n521), .A2(G74), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n588), .A2(G651), .B1(G49), .B2(new_n512), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n582), .A2(G87), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(G288));
  AOI22_X1  g166(.A1(new_n521), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n506), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n512), .A2(G48), .ZN(new_n594));
  INV_X1    g169(.A(G86), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n523), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(new_n506), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n512), .A2(G47), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n523), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n521), .A2(G66), .ZN(new_n607));
  INV_X1    g182(.A(G79), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(new_n511), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(G651), .B1(G54), .B2(new_n512), .ZN(new_n610));
  INV_X1    g185(.A(G92), .ZN(new_n611));
  OAI21_X1  g186(.A(KEYINPUT10), .B1(new_n523), .B2(new_n611), .ZN(new_n612));
  OR3_X1    g187(.A1(new_n523), .A2(KEYINPUT10), .A3(new_n611), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n606), .B1(new_n615), .B2(G868), .ZN(G284));
  OAI21_X1  g191(.A(new_n606), .B1(new_n615), .B2(G868), .ZN(G321));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(G299), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G168), .B2(new_n618), .ZN(G297));
  OAI21_X1  g195(.A(new_n619), .B1(G168), .B2(new_n618), .ZN(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n615), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND2_X1  g198(.A1(new_n615), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n566), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g202(.A(new_n489), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G123), .ZN(new_n629));
  INV_X1    g204(.A(G135), .ZN(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n465), .A2(G111), .ZN(new_n632));
  OAI221_X1 g207(.A(new_n629), .B1(new_n630), .B2(new_n490), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2096), .Z(new_n634));
  NAND3_X1  g209(.A1(new_n465), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT81), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(KEYINPUT80), .B(G2100), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n634), .B(new_n641), .C1(new_n638), .C2(new_n637), .ZN(G156));
  XOR2_X1   g217(.A(G2427), .B(G2430), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT83), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT82), .B(G2438), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(KEYINPUT14), .ZN(new_n649));
  XOR2_X1   g224(.A(G2443), .B(G2446), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G1341), .B(G1348), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n651), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n654), .B(new_n655), .Z(new_n656));
  AND2_X1   g231(.A1(new_n656), .A2(G14), .ZN(G401));
  XOR2_X1   g232(.A(G2067), .B(G2678), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n661), .A2(KEYINPUT17), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n659), .A2(new_n660), .ZN(new_n663));
  AOI21_X1  g238(.A(KEYINPUT18), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2096), .ZN(new_n665));
  XOR2_X1   g240(.A(G2072), .B(G2078), .Z(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n661), .B2(KEYINPUT18), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n665), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT84), .B(G2100), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G227));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT85), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT20), .Z(new_n678));
  NOR2_X1   g253(.A1(new_n673), .A2(new_n674), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n680), .A2(new_n672), .A3(new_n675), .ZN(new_n681));
  OAI211_X1 g256(.A(new_n678), .B(new_n681), .C1(new_n672), .C2(new_n680), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT86), .B(G1981), .Z(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n685), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G229));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G25), .ZN(new_n692));
  INV_X1    g267(.A(new_n490), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G131), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n628), .A2(G119), .ZN(new_n695));
  OR2_X1    g270(.A1(G95), .A2(G2105), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n696), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n694), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n692), .B1(new_n699), .B2(new_n691), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT35), .B(G1991), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT87), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n700), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n604), .A2(G16), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G16), .B2(G24), .ZN(new_n705));
  INV_X1    g280(.A(G1986), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n703), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n589), .B2(new_n590), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT33), .B(G1976), .Z(new_n712));
  AND2_X1   g287(.A1(new_n710), .A2(G23), .ZN(new_n713));
  OR3_X1    g288(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n712), .B1(new_n711), .B2(new_n713), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT89), .B(KEYINPUT90), .Z(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n717), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n714), .A2(new_n719), .A3(new_n715), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  OR2_X1    g297(.A1(G16), .A2(G22), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G303), .B2(new_n710), .ZN(new_n724));
  INV_X1    g299(.A(G1971), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n597), .A2(new_n710), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n710), .A2(G6), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT88), .B(G1981), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT32), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  OR3_X1    g306(.A1(new_n727), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n727), .B2(new_n728), .ZN(new_n733));
  OAI211_X1 g308(.A(G1971), .B(new_n723), .C1(G303), .C2(new_n710), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n726), .A2(new_n732), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(KEYINPUT91), .B1(new_n722), .B2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n735), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT91), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n737), .A2(new_n738), .A3(new_n721), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(KEYINPUT34), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT34), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n736), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n709), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n744), .A2(KEYINPUT92), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n744), .A2(KEYINPUT92), .A3(KEYINPUT93), .A4(KEYINPUT36), .ZN(new_n746));
  INV_X1    g321(.A(new_n709), .ZN(new_n747));
  INV_X1    g322(.A(new_n743), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n742), .B1(new_n736), .B2(new_n739), .ZN(new_n749));
  OAI211_X1 g324(.A(KEYINPUT93), .B(new_n747), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT36), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n746), .A2(new_n752), .ZN(new_n753));
  OR2_X1    g328(.A1(G16), .A2(G21), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G286), .B2(new_n710), .ZN(new_n755));
  INV_X1    g330(.A(G1966), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT100), .B(KEYINPUT30), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G28), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n755), .A2(new_n756), .B1(new_n691), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT31), .B(G11), .ZN(new_n761));
  AND3_X1   g336(.A1(new_n757), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G1961), .ZN(new_n763));
  NAND2_X1  g338(.A1(G171), .A2(G16), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G5), .B2(G16), .ZN(new_n765));
  OAI221_X1 g340(.A(new_n762), .B1(new_n691), .B2(new_n633), .C1(new_n763), .C2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT101), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n765), .A2(new_n763), .ZN(new_n769));
  NOR2_X1   g344(.A1(G29), .A2(G35), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G162), .B2(G29), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT29), .Z(new_n772));
  INV_X1    g347(.A(G2090), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(G299), .A2(G16), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n710), .A2(KEYINPUT23), .A3(G20), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT23), .ZN(new_n777));
  INV_X1    g352(.A(G20), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n778), .B2(G16), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n775), .A2(new_n776), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1956), .ZN(new_n781));
  NOR2_X1   g356(.A1(G164), .A2(new_n691), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G27), .B2(new_n691), .ZN(new_n783));
  INV_X1    g358(.A(G2078), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  NOR3_X1   g361(.A1(new_n781), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT25), .Z(new_n789));
  INV_X1    g364(.A(G139), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n490), .B2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT98), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n462), .A2(new_n477), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n795), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n796));
  OAI22_X1  g371(.A1(new_n793), .A2(new_n794), .B1(new_n465), .B2(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G33), .B(new_n797), .S(G29), .Z(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(G2072), .ZN(new_n799));
  NOR2_X1   g374(.A1(G4), .A2(G16), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n615), .B2(G16), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT94), .B(G1348), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n774), .A2(new_n787), .A3(new_n799), .A4(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n798), .A2(G2072), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n772), .B2(new_n773), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n691), .A2(G26), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT97), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT28), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n628), .A2(G128), .ZN(new_n810));
  INV_X1    g385(.A(G140), .ZN(new_n811));
  OAI21_X1  g386(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n465), .A2(G116), .ZN(new_n813));
  OAI221_X1 g388(.A(new_n810), .B1(new_n811), .B2(new_n490), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G29), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n815), .A2(KEYINPUT96), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(KEYINPUT96), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n809), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(G2067), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  OR2_X1    g395(.A1(KEYINPUT24), .A2(G34), .ZN(new_n821));
  NAND2_X1  g396(.A1(KEYINPUT24), .A2(G34), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n821), .A2(new_n691), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G160), .B2(new_n691), .ZN(new_n824));
  INV_X1    g399(.A(G2084), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n806), .A2(new_n820), .A3(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n804), .A2(new_n827), .ZN(new_n828));
  AND3_X1   g403(.A1(new_n768), .A2(new_n769), .A3(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT102), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n693), .A2(G141), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n628), .A2(G129), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n465), .A2(G105), .A3(G2104), .ZN(new_n833));
  NAND3_X1  g408(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT26), .Z(new_n835));
  NAND4_X1  g410(.A1(new_n831), .A2(new_n832), .A3(new_n833), .A4(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT99), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(G29), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(G29), .B2(G32), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT27), .B(G1996), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(G16), .A2(G19), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(new_n566), .B2(G16), .ZN(new_n845));
  XOR2_X1   g420(.A(KEYINPUT95), .B(G1341), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n829), .A2(new_n830), .A3(new_n843), .A4(new_n847), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n768), .A2(new_n828), .A3(new_n847), .A4(new_n769), .ZN(new_n849));
  OAI21_X1  g424(.A(KEYINPUT102), .B1(new_n849), .B2(new_n842), .ZN(new_n850));
  AOI211_X1 g425(.A(new_n745), .B(new_n753), .C1(new_n848), .C2(new_n850), .ZN(G311));
  NAND2_X1  g426(.A1(new_n848), .A2(new_n850), .ZN(new_n852));
  INV_X1    g427(.A(new_n753), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n852), .B(new_n853), .C1(KEYINPUT92), .C2(new_n744), .ZN(G150));
  AOI22_X1  g429(.A1(new_n582), .A2(G93), .B1(G55), .B2(new_n512), .ZN(new_n855));
  AOI22_X1  g430(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n855), .B1(new_n506), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(G860), .ZN(new_n858));
  XOR2_X1   g433(.A(KEYINPUT103), .B(KEYINPUT37), .Z(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n857), .B(new_n566), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT39), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n615), .A2(G559), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT38), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n862), .B(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n860), .B1(new_n865), .B2(G860), .ZN(G145));
  INV_X1    g441(.A(new_n504), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT104), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n869));
  INV_X1    g444(.A(new_n498), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI211_X1 g446(.A(KEYINPUT104), .B(new_n498), .C1(new_n499), .C2(KEYINPUT4), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n867), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n814), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n837), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT105), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n875), .B1(new_n876), .B2(new_n797), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n877), .B(new_n636), .Z(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(G160), .B(new_n633), .ZN(new_n880));
  INV_X1    g455(.A(G162), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n797), .A2(new_n876), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n698), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n880), .B(G162), .ZN(new_n886));
  INV_X1    g461(.A(new_n884), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n693), .A2(G142), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n628), .A2(G130), .ZN(new_n890));
  OAI21_X1  g465(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT106), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n892), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n893), .B(new_n894), .C1(G118), .C2(new_n465), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n889), .A2(new_n890), .A3(new_n895), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n885), .A2(new_n888), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n896), .B1(new_n885), .B2(new_n888), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n879), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n896), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n886), .A2(new_n887), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n882), .A2(new_n884), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n885), .A2(new_n888), .A3(new_n896), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(new_n878), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n899), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g483(.A1(new_n857), .A2(new_n618), .ZN(new_n909));
  XNOR2_X1  g484(.A(G288), .B(new_n597), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n910), .A2(G290), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(G290), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n912), .A2(G166), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(G166), .B1(new_n912), .B2(new_n913), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT42), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n861), .B(new_n624), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n614), .B(G299), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  XOR2_X1   g496(.A(new_n919), .B(KEYINPUT41), .Z(new_n922));
  AOI21_X1  g497(.A(new_n921), .B1(new_n922), .B2(new_n918), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n917), .B(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n909), .B1(new_n924), .B2(new_n618), .ZN(G295));
  OAI21_X1  g500(.A(new_n909), .B1(new_n924), .B2(new_n618), .ZN(G331));
  XNOR2_X1  g501(.A(G286), .B(G301), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(new_n861), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n920), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n922), .A2(new_n928), .ZN(new_n931));
  OAI22_X1  g506(.A1(new_n930), .A2(new_n931), .B1(new_n914), .B2(new_n915), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT107), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n906), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n916), .B(new_n929), .C1(new_n922), .C2(new_n928), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n935), .B1(new_n932), .B2(KEYINPUT107), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT43), .ZN(new_n937));
  NOR3_X1   g512(.A1(new_n934), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n932), .A2(new_n935), .A3(new_n906), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n939), .A2(new_n937), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT44), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n934), .A2(new_n936), .A3(KEYINPUT43), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n941), .B1(new_n945), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g521(.A(G1384), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n873), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT45), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n483), .A2(new_n472), .A3(G40), .A4(new_n473), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OR2_X1    g527(.A1(new_n837), .A2(G1996), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n814), .B(new_n819), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n837), .A2(G1996), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n699), .A2(new_n702), .ZN(new_n958));
  OR2_X1    g533(.A1(new_n699), .A2(new_n702), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(G290), .A2(G1986), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n961), .A2(KEYINPUT108), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n604), .A2(new_n706), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n962), .B(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n952), .B1(new_n960), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G288), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(G1976), .ZN(new_n967));
  AND4_X1   g542(.A1(G40), .A2(new_n483), .A3(new_n472), .A4(new_n473), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n968), .A2(new_n947), .A3(new_n873), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n970));
  XNOR2_X1  g545(.A(KEYINPUT111), .B(G8), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n970), .B1(new_n969), .B2(new_n971), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n967), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT113), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI211_X1 g551(.A(KEYINPUT113), .B(new_n967), .C1(new_n972), .C2(new_n973), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(new_n977), .A3(KEYINPUT52), .ZN(new_n978));
  OR2_X1    g553(.A1(new_n972), .A2(new_n973), .ZN(new_n979));
  NAND2_X1  g554(.A1(G305), .A2(G1981), .ZN(new_n980));
  OR3_X1    g555(.A1(new_n593), .A2(new_n596), .A3(G1981), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT115), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT49), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n982), .B(new_n985), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n979), .B(new_n986), .C1(new_n983), .C2(new_n984), .ZN(new_n987));
  INV_X1    g562(.A(G1976), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT52), .B1(G288), .B2(new_n988), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n967), .B(new_n989), .C1(new_n972), .C2(new_n973), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT114), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT114), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n979), .A2(new_n992), .A3(new_n967), .A4(new_n989), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n978), .A2(new_n987), .A3(new_n991), .A4(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n947), .B1(new_n500), .B2(new_n504), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n949), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT109), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT109), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n996), .A2(new_n999), .A3(new_n949), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n998), .A2(new_n968), .A3(new_n1000), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n873), .A2(KEYINPUT45), .A3(new_n947), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n995), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n951), .B1(new_n997), .B2(KEYINPUT109), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n873), .A2(KEYINPUT45), .A3(new_n947), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1004), .A2(new_n1005), .A3(KEYINPUT110), .A4(new_n1000), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n725), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n951), .B1(KEYINPUT50), .B2(new_n996), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n873), .A2(new_n1010), .A3(new_n947), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1012), .A2(G2090), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1008), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(G303), .A2(G8), .ZN(new_n1016));
  XOR2_X1   g591(.A(new_n1016), .B(KEYINPUT55), .Z(new_n1017));
  NAND3_X1  g592(.A1(new_n1015), .A2(G8), .A3(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n994), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n972), .A2(new_n973), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n987), .A2(new_n988), .A3(new_n966), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1020), .B1(new_n1021), .B2(new_n981), .ZN(new_n1022));
  OR2_X1    g597(.A1(new_n500), .A2(new_n504), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1023), .A2(KEYINPUT45), .A3(new_n947), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n950), .A2(new_n968), .A3(new_n1024), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1025), .A2(new_n756), .B1(new_n1026), .B2(new_n825), .ZN(new_n1027));
  INV_X1    g602(.A(new_n971), .ZN(new_n1028));
  OR3_X1    g603(.A1(new_n1027), .A2(G286), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(KEYINPUT117), .B(KEYINPUT63), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n1019), .A2(new_n1022), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1010), .B1(new_n873), .B2(new_n947), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1023), .A2(new_n1010), .A3(new_n947), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n1035), .A2(new_n1037), .A3(new_n951), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n773), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1028), .B1(new_n1008), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1018), .B1(new_n1040), .B2(new_n1017), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n994), .A2(KEYINPUT116), .ZN(new_n1042));
  XNOR2_X1  g617(.A(new_n990), .B(new_n992), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1043), .A2(new_n1044), .A3(new_n987), .A4(new_n978), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1041), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT62), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT123), .B1(G168), .B2(new_n1028), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT123), .ZN(new_n1049));
  NAND3_X1  g624(.A1(G286), .A2(new_n1049), .A3(new_n971), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1027), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G8), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1053), .B(KEYINPUT51), .C1(new_n1027), .C2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT51), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1058), .B(new_n1052), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1047), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1056), .A2(new_n1059), .A3(KEYINPUT62), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1003), .A2(new_n784), .A3(new_n1006), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT125), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1026), .A2(G1961), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT125), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1063), .A2(new_n1069), .A3(new_n1064), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n950), .A2(new_n968), .A3(new_n1024), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1064), .A2(G2078), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1066), .A2(new_n1068), .A3(new_n1070), .A4(new_n1073), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1062), .A2(G171), .A3(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1046), .A2(new_n1061), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G1348), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1012), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n969), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n819), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1078), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(G1348), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n969), .A2(G2067), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT120), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1082), .A2(new_n1085), .A3(new_n615), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT121), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n581), .A2(new_n583), .A3(new_n585), .A4(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1091), .B(new_n1092), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1093), .A2(KEYINPUT122), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1093), .A2(KEYINPUT122), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1035), .A2(new_n951), .ZN(new_n1096));
  AOI21_X1  g671(.A(G1956), .B1(new_n1096), .B2(new_n1036), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT56), .B(G2072), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1004), .A2(new_n1005), .A3(new_n1000), .A4(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  OAI22_X1  g675(.A1(new_n1094), .A2(new_n1095), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1082), .A2(new_n1085), .A3(new_n1102), .A4(new_n615), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1087), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1092), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1091), .B(new_n1105), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1099), .B(new_n1106), .C1(new_n1038), .C2(G1956), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT119), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n948), .A2(KEYINPUT50), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1109), .A2(new_n1036), .A3(new_n968), .ZN(new_n1110));
  INV_X1    g685(.A(G1956), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1112), .A2(new_n1113), .A3(new_n1099), .A4(new_n1106), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1104), .A2(new_n1108), .A3(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1093), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1108), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT61), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1101), .A2(KEYINPUT61), .A3(new_n1107), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1004), .A2(new_n1005), .A3(new_n1000), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT58), .B(G1341), .ZN(new_n1122));
  OAI22_X1  g697(.A1(new_n1121), .A2(G1996), .B1(new_n1079), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n566), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1124), .B(KEYINPUT59), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1119), .A2(new_n1120), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1081), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1083), .A2(new_n1084), .A3(KEYINPUT120), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1127), .A2(new_n1128), .A3(KEYINPUT60), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT60), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n615), .ZN(new_n1131));
  OAI211_X1 g706(.A(KEYINPUT60), .B(new_n614), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1129), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1115), .B1(new_n1126), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1046), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1063), .A2(new_n1069), .A3(new_n1064), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1069), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1139), .A2(G301), .A3(new_n1068), .A4(new_n1073), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n950), .A2(G40), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1141), .B1(G2105), .B2(new_n480), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1142), .A2(new_n474), .A3(new_n1005), .A4(new_n1072), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1066), .A2(new_n1068), .A3(new_n1070), .A4(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(G171), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1140), .A2(new_n1145), .A3(KEYINPUT54), .ZN(new_n1146));
  NOR4_X1   g721(.A1(new_n1137), .A2(new_n1138), .A3(G171), .A4(new_n1067), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1147), .A2(new_n1143), .B1(G171), .B2(new_n1074), .ZN(new_n1148));
  XNOR2_X1  g723(.A(KEYINPUT124), .B(KEYINPUT54), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1146), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1034), .B(new_n1076), .C1(new_n1136), .C2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1054), .B1(new_n1008), .B2(new_n1014), .ZN(new_n1152));
  OAI21_X1  g727(.A(KEYINPUT63), .B1(new_n1152), .B2(new_n1017), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n994), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1046), .A2(new_n1030), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1154), .B1(new_n1155), .B2(new_n1032), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n965), .B1(new_n1151), .B2(new_n1156), .ZN(new_n1157));
  OAI22_X1  g732(.A1(new_n956), .A2(new_n958), .B1(G2067), .B2(new_n814), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1158), .A2(new_n952), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n950), .A2(G1996), .A3(new_n951), .ZN(new_n1160));
  OR2_X1    g735(.A1(new_n1160), .A2(KEYINPUT46), .ZN(new_n1161));
  INV_X1    g736(.A(new_n954), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n952), .B1(new_n1162), .B2(new_n837), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1160), .A2(KEYINPUT46), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1161), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1165), .B(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n960), .A2(new_n952), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n952), .A2(new_n961), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1169), .B(KEYINPUT127), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1170), .B(KEYINPUT48), .ZN(new_n1171));
  AOI211_X1 g746(.A(new_n1159), .B(new_n1167), .C1(new_n1168), .C2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1157), .A2(new_n1172), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g748(.A(G319), .ZN(new_n1175));
  AOI211_X1 g749(.A(new_n1175), .B(G227), .C1(new_n656), .C2(G14), .ZN(new_n1176));
  NAND2_X1  g750(.A1(new_n907), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g751(.A(new_n689), .B1(new_n942), .B2(new_n944), .ZN(new_n1178));
  NOR2_X1   g752(.A1(new_n1177), .A2(new_n1178), .ZN(G308));
  INV_X1    g753(.A(new_n945), .ZN(new_n1180));
  NAND4_X1  g754(.A1(new_n1180), .A2(new_n689), .A3(new_n907), .A4(new_n1176), .ZN(G225));
endmodule


