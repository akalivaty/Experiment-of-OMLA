

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582;

  XNOR2_X1 U326 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U327 ( .A(KEYINPUT28), .B(n470), .Z(n528) );
  XOR2_X1 U328 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n294) );
  XOR2_X1 U329 ( .A(G43GAT), .B(G134GAT), .Z(n295) );
  XOR2_X1 U330 ( .A(n372), .B(n371), .Z(n296) );
  XNOR2_X1 U331 ( .A(KEYINPUT121), .B(KEYINPUT54), .ZN(n467) );
  XNOR2_X1 U332 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U333 ( .A(n367), .B(KEYINPUT100), .ZN(n368) );
  XNOR2_X1 U334 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U335 ( .A(n379), .B(n295), .ZN(n380) );
  XNOR2_X1 U336 ( .A(n536), .B(n368), .ZN(n580) );
  NOR2_X1 U337 ( .A1(n474), .A2(n473), .ZN(n562) );
  NOR2_X1 U338 ( .A1(n504), .A2(n490), .ZN(n521) );
  XNOR2_X1 U339 ( .A(n381), .B(n380), .ZN(n525) );
  XNOR2_X1 U340 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n475) );
  XNOR2_X1 U341 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U342 ( .A(n476), .B(n475), .ZN(G1351GAT) );
  XNOR2_X1 U343 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n314) );
  XOR2_X1 U344 ( .A(KEYINPUT76), .B(KEYINPUT75), .Z(n298) );
  XNOR2_X1 U345 ( .A(KEYINPUT74), .B(KEYINPUT73), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n298), .B(n297), .ZN(n313) );
  XOR2_X1 U347 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n300) );
  NAND2_X1 U348 ( .A1(G230GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U349 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U350 ( .A(n301), .B(KEYINPUT31), .Z(n305) );
  XNOR2_X1 U351 ( .A(G99GAT), .B(G106GAT), .ZN(n302) );
  XNOR2_X1 U352 ( .A(n302), .B(G85GAT), .ZN(n361) );
  XNOR2_X1 U353 ( .A(G71GAT), .B(G57GAT), .ZN(n303) );
  XNOR2_X1 U354 ( .A(n303), .B(KEYINPUT13), .ZN(n343) );
  XNOR2_X1 U355 ( .A(n361), .B(n343), .ZN(n304) );
  XNOR2_X1 U356 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U357 ( .A(G176GAT), .B(G64GAT), .Z(n403) );
  XOR2_X1 U358 ( .A(KEYINPUT72), .B(n403), .Z(n307) );
  XOR2_X1 U359 ( .A(G148GAT), .B(G78GAT), .Z(n385) );
  XNOR2_X1 U360 ( .A(G204GAT), .B(n385), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U362 ( .A(n309), .B(n308), .Z(n311) );
  XNOR2_X1 U363 ( .A(G120GAT), .B(G92GAT), .ZN(n310) );
  XNOR2_X1 U364 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n313), .B(n312), .ZN(n571) );
  XNOR2_X1 U366 ( .A(n314), .B(n571), .ZN(n555) );
  XOR2_X1 U367 ( .A(G197GAT), .B(G22GAT), .Z(n316) );
  XNOR2_X1 U368 ( .A(G50GAT), .B(G36GAT), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U370 ( .A(n317), .B(G15GAT), .Z(n319) );
  XOR2_X1 U371 ( .A(G113GAT), .B(G1GAT), .Z(n433) );
  XNOR2_X1 U372 ( .A(G169GAT), .B(n433), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n319), .B(n318), .ZN(n325) );
  XOR2_X1 U374 ( .A(G29GAT), .B(G43GAT), .Z(n321) );
  XNOR2_X1 U375 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n320) );
  XNOR2_X1 U376 ( .A(n321), .B(n320), .ZN(n358) );
  XOR2_X1 U377 ( .A(n358), .B(KEYINPUT67), .Z(n323) );
  NAND2_X1 U378 ( .A1(G229GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U379 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U380 ( .A(n325), .B(n324), .Z(n333) );
  XOR2_X1 U381 ( .A(KEYINPUT30), .B(KEYINPUT70), .Z(n327) );
  XNOR2_X1 U382 ( .A(G141GAT), .B(KEYINPUT71), .ZN(n326) );
  XNOR2_X1 U383 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U384 ( .A(G8GAT), .B(KEYINPUT69), .Z(n329) );
  XNOR2_X1 U385 ( .A(KEYINPUT29), .B(KEYINPUT68), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U387 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U388 ( .A(n333), .B(n332), .Z(n567) );
  NAND2_X1 U389 ( .A1(n555), .A2(n567), .ZN(n334) );
  XNOR2_X1 U390 ( .A(n334), .B(KEYINPUT106), .ZN(n504) );
  XOR2_X1 U391 ( .A(KEYINPUT14), .B(G64GAT), .Z(n336) );
  XNOR2_X1 U392 ( .A(G1GAT), .B(G78GAT), .ZN(n335) );
  XNOR2_X1 U393 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U394 ( .A(KEYINPUT84), .B(KEYINPUT12), .Z(n338) );
  XNOR2_X1 U395 ( .A(KEYINPUT83), .B(KEYINPUT82), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U397 ( .A(n340), .B(n339), .ZN(n350) );
  XOR2_X1 U398 ( .A(KEYINPUT81), .B(G211GAT), .Z(n342) );
  XNOR2_X1 U399 ( .A(G8GAT), .B(G183GAT), .ZN(n341) );
  XNOR2_X1 U400 ( .A(n342), .B(n341), .ZN(n406) );
  XOR2_X1 U401 ( .A(KEYINPUT15), .B(n343), .Z(n345) );
  NAND2_X1 U402 ( .A1(G231GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U404 ( .A(n406), .B(n346), .Z(n348) );
  XOR2_X1 U405 ( .A(G15GAT), .B(G127GAT), .Z(n370) );
  XOR2_X1 U406 ( .A(G22GAT), .B(G155GAT), .Z(n386) );
  XNOR2_X1 U407 ( .A(n370), .B(n386), .ZN(n347) );
  XNOR2_X1 U408 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U409 ( .A(n350), .B(n349), .Z(n575) );
  XOR2_X1 U410 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n352) );
  XNOR2_X1 U411 ( .A(KEYINPUT66), .B(KEYINPUT11), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n352), .B(n351), .ZN(n366) );
  XOR2_X1 U413 ( .A(KEYINPUT10), .B(KEYINPUT77), .Z(n354) );
  NAND2_X1 U414 ( .A1(G232GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U415 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U416 ( .A(n355), .B(KEYINPUT79), .ZN(n360) );
  XOR2_X1 U417 ( .A(G92GAT), .B(G218GAT), .Z(n357) );
  XNOR2_X1 U418 ( .A(G36GAT), .B(G190GAT), .ZN(n356) );
  XNOR2_X1 U419 ( .A(n357), .B(n356), .ZN(n408) );
  XNOR2_X1 U420 ( .A(n358), .B(n408), .ZN(n359) );
  XNOR2_X1 U421 ( .A(n360), .B(n359), .ZN(n364) );
  XOR2_X1 U422 ( .A(G50GAT), .B(G162GAT), .Z(n389) );
  XOR2_X1 U423 ( .A(G134GAT), .B(KEYINPUT78), .Z(n429) );
  XNOR2_X1 U424 ( .A(n389), .B(n429), .ZN(n362) );
  XNOR2_X1 U425 ( .A(n366), .B(n365), .ZN(n551) );
  XOR2_X1 U426 ( .A(KEYINPUT80), .B(n551), .Z(n536) );
  INV_X1 U427 ( .A(KEYINPUT36), .ZN(n367) );
  INV_X1 U428 ( .A(KEYINPUT97), .ZN(n448) );
  XNOR2_X1 U429 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n369) );
  XNOR2_X1 U430 ( .A(n294), .B(n369), .ZN(n409) );
  XOR2_X1 U431 ( .A(n409), .B(n370), .Z(n372) );
  NAND2_X1 U432 ( .A1(G227GAT), .A2(G233GAT), .ZN(n371) );
  XOR2_X1 U433 ( .A(KEYINPUT0), .B(G120GAT), .Z(n428) );
  XNOR2_X1 U434 ( .A(n296), .B(n428), .ZN(n381) );
  XOR2_X1 U435 ( .A(KEYINPUT20), .B(G99GAT), .Z(n374) );
  XNOR2_X1 U436 ( .A(G113GAT), .B(G190GAT), .ZN(n373) );
  XNOR2_X1 U437 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U438 ( .A(G71GAT), .B(G176GAT), .Z(n376) );
  XNOR2_X1 U439 ( .A(KEYINPUT86), .B(G183GAT), .ZN(n375) );
  XNOR2_X1 U440 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U441 ( .A(n378), .B(n377), .Z(n379) );
  XOR2_X1 U442 ( .A(G204GAT), .B(KEYINPUT21), .Z(n383) );
  XNOR2_X1 U443 ( .A(G197GAT), .B(KEYINPUT89), .ZN(n382) );
  XNOR2_X1 U444 ( .A(n383), .B(n382), .ZN(n413) );
  XNOR2_X1 U445 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n384) );
  XOR2_X1 U446 ( .A(n384), .B(KEYINPUT2), .Z(n437) );
  XNOR2_X1 U447 ( .A(n413), .B(n437), .ZN(n400) );
  XOR2_X1 U448 ( .A(n386), .B(n385), .Z(n388) );
  NAND2_X1 U449 ( .A1(G228GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U450 ( .A(n388), .B(n387), .ZN(n390) );
  XOR2_X1 U451 ( .A(n390), .B(n389), .Z(n398) );
  XOR2_X1 U452 ( .A(KEYINPUT22), .B(G211GAT), .Z(n392) );
  XNOR2_X1 U453 ( .A(G218GAT), .B(G106GAT), .ZN(n391) );
  XNOR2_X1 U454 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U455 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n394) );
  XNOR2_X1 U456 ( .A(KEYINPUT87), .B(KEYINPUT88), .ZN(n393) );
  XNOR2_X1 U457 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U458 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U459 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U460 ( .A(n400), .B(n399), .ZN(n470) );
  NOR2_X1 U461 ( .A1(n525), .A2(n470), .ZN(n401) );
  XOR2_X1 U462 ( .A(KEYINPUT26), .B(n401), .Z(n402) );
  XOR2_X1 U463 ( .A(KEYINPUT94), .B(n402), .Z(n565) );
  XOR2_X1 U464 ( .A(KEYINPUT93), .B(n403), .Z(n405) );
  NAND2_X1 U465 ( .A1(G226GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U466 ( .A(n405), .B(n404), .ZN(n407) );
  XOR2_X1 U467 ( .A(n407), .B(n406), .Z(n411) );
  XNOR2_X1 U468 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U469 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U470 ( .A(n413), .B(n412), .ZN(n519) );
  XNOR2_X1 U471 ( .A(n519), .B(KEYINPUT27), .ZN(n443) );
  NAND2_X1 U472 ( .A1(n565), .A2(n443), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n414), .B(KEYINPUT95), .ZN(n419) );
  NAND2_X1 U474 ( .A1(n519), .A2(n525), .ZN(n415) );
  NAND2_X1 U475 ( .A1(n415), .A2(n470), .ZN(n416) );
  XNOR2_X1 U476 ( .A(n416), .B(KEYINPUT96), .ZN(n417) );
  XNOR2_X1 U477 ( .A(KEYINPUT25), .B(n417), .ZN(n418) );
  NOR2_X1 U478 ( .A1(n419), .A2(n418), .ZN(n442) );
  XOR2_X1 U479 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n421) );
  XNOR2_X1 U480 ( .A(KEYINPUT90), .B(KEYINPUT92), .ZN(n420) );
  XNOR2_X1 U481 ( .A(n421), .B(n420), .ZN(n441) );
  XOR2_X1 U482 ( .A(G85GAT), .B(G162GAT), .Z(n423) );
  XNOR2_X1 U483 ( .A(G29GAT), .B(G127GAT), .ZN(n422) );
  XNOR2_X1 U484 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U485 ( .A(KEYINPUT1), .B(G57GAT), .Z(n425) );
  XNOR2_X1 U486 ( .A(G155GAT), .B(G148GAT), .ZN(n424) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U488 ( .A(n427), .B(n426), .Z(n435) );
  XOR2_X1 U489 ( .A(n429), .B(n428), .Z(n431) );
  NAND2_X1 U490 ( .A1(G225GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U491 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U492 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U494 ( .A(n436), .B(KEYINPUT91), .Z(n439) );
  XOR2_X1 U495 ( .A(n437), .B(KEYINPUT6), .Z(n438) );
  XNOR2_X1 U496 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U497 ( .A(n441), .B(n440), .ZN(n517) );
  NOR2_X1 U498 ( .A1(n442), .A2(n517), .ZN(n446) );
  NAND2_X1 U499 ( .A1(n443), .A2(n517), .ZN(n523) );
  OR2_X1 U500 ( .A1(n528), .A2(n525), .ZN(n444) );
  NOR2_X1 U501 ( .A1(n523), .A2(n444), .ZN(n445) );
  NOR2_X1 U502 ( .A1(n446), .A2(n445), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n448), .B(n447), .ZN(n480) );
  NOR2_X1 U504 ( .A1(n580), .A2(n480), .ZN(n449) );
  NAND2_X1 U505 ( .A1(n575), .A2(n449), .ZN(n450) );
  XOR2_X1 U506 ( .A(KEYINPUT37), .B(n450), .Z(n490) );
  NAND2_X1 U507 ( .A1(n521), .A2(n528), .ZN(n454) );
  XOR2_X1 U508 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n452) );
  XNOR2_X1 U509 ( .A(G106GAT), .B(KEYINPUT110), .ZN(n451) );
  XNOR2_X1 U510 ( .A(n454), .B(n453), .ZN(G1339GAT) );
  INV_X1 U511 ( .A(KEYINPUT55), .ZN(n472) );
  XOR2_X1 U512 ( .A(KEYINPUT47), .B(KEYINPUT113), .Z(n459) );
  XOR2_X1 U513 ( .A(KEYINPUT112), .B(n575), .Z(n563) );
  INV_X1 U514 ( .A(n567), .ZN(n553) );
  NAND2_X1 U515 ( .A1(n553), .A2(n555), .ZN(n455) );
  XOR2_X1 U516 ( .A(KEYINPUT46), .B(n455), .Z(n456) );
  NOR2_X1 U517 ( .A1(n563), .A2(n456), .ZN(n457) );
  NAND2_X1 U518 ( .A1(n457), .A2(n551), .ZN(n458) );
  XNOR2_X1 U519 ( .A(n459), .B(n458), .ZN(n464) );
  NOR2_X1 U520 ( .A1(n580), .A2(n575), .ZN(n460) );
  XNOR2_X1 U521 ( .A(n460), .B(KEYINPUT45), .ZN(n461) );
  NAND2_X1 U522 ( .A1(n461), .A2(n571), .ZN(n462) );
  NOR2_X1 U523 ( .A1(n553), .A2(n462), .ZN(n463) );
  NOR2_X1 U524 ( .A1(n464), .A2(n463), .ZN(n465) );
  XNOR2_X1 U525 ( .A(KEYINPUT48), .B(n465), .ZN(n524) );
  XOR2_X1 U526 ( .A(n519), .B(KEYINPUT120), .Z(n466) );
  NOR2_X1 U527 ( .A1(n524), .A2(n466), .ZN(n468) );
  NOR2_X1 U528 ( .A1(n469), .A2(n517), .ZN(n566) );
  NAND2_X1 U529 ( .A1(n566), .A2(n470), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n472), .B(n471), .ZN(n474) );
  INV_X1 U531 ( .A(n525), .ZN(n473) );
  NAND2_X1 U532 ( .A1(n536), .A2(n562), .ZN(n476) );
  XOR2_X1 U533 ( .A(KEYINPUT85), .B(KEYINPUT16), .Z(n478) );
  OR2_X1 U534 ( .A1(n536), .A2(n575), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n478), .B(n477), .ZN(n479) );
  NOR2_X1 U536 ( .A1(n480), .A2(n479), .ZN(n481) );
  XOR2_X1 U537 ( .A(KEYINPUT98), .B(n481), .Z(n505) );
  NAND2_X1 U538 ( .A1(n553), .A2(n571), .ZN(n491) );
  NOR2_X1 U539 ( .A1(n505), .A2(n491), .ZN(n488) );
  NAND2_X1 U540 ( .A1(n517), .A2(n488), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(KEYINPUT34), .ZN(n483) );
  XNOR2_X1 U542 ( .A(G1GAT), .B(n483), .ZN(G1324GAT) );
  NAND2_X1 U543 ( .A1(n519), .A2(n488), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n484), .B(G8GAT), .ZN(G1325GAT) );
  XNOR2_X1 U545 ( .A(KEYINPUT99), .B(KEYINPUT35), .ZN(n486) );
  AND2_X1 U546 ( .A1(n488), .A2(n525), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U548 ( .A(G15GAT), .B(n487), .Z(G1326GAT) );
  NAND2_X1 U549 ( .A1(n528), .A2(n488), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n489), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U551 ( .A1(n491), .A2(n490), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n492), .B(KEYINPUT38), .ZN(n501) );
  NAND2_X1 U553 ( .A1(n517), .A2(n501), .ZN(n494) );
  XOR2_X1 U554 ( .A(G29GAT), .B(KEYINPUT39), .Z(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  NAND2_X1 U556 ( .A1(n501), .A2(n519), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n495), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n497) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(KEYINPUT102), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U561 ( .A(KEYINPUT101), .B(n498), .Z(n500) );
  NAND2_X1 U562 ( .A1(n525), .A2(n501), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(G1330GAT) );
  XNOR2_X1 U564 ( .A(G50GAT), .B(KEYINPUT104), .ZN(n503) );
  NAND2_X1 U565 ( .A1(n528), .A2(n501), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n503), .B(n502), .ZN(G1331GAT) );
  XOR2_X1 U567 ( .A(G57GAT), .B(KEYINPUT105), .Z(n507) );
  NOR2_X1 U568 ( .A1(n505), .A2(n504), .ZN(n513) );
  NAND2_X1 U569 ( .A1(n513), .A2(n517), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n507), .B(n506), .ZN(n509) );
  XOR2_X1 U571 ( .A(KEYINPUT42), .B(KEYINPUT107), .Z(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(G1332GAT) );
  NAND2_X1 U573 ( .A1(n519), .A2(n513), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n510), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U575 ( .A1(n513), .A2(n525), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n511), .B(KEYINPUT108), .ZN(n512) );
  XNOR2_X1 U577 ( .A(G71GAT), .B(n512), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n515) );
  NAND2_X1 U579 ( .A1(n513), .A2(n528), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(n516) );
  XOR2_X1 U581 ( .A(G78GAT), .B(n516), .Z(G1335GAT) );
  NAND2_X1 U582 ( .A1(n521), .A2(n517), .ZN(n518) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n518), .ZN(G1336GAT) );
  NAND2_X1 U584 ( .A1(n519), .A2(n521), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n520), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U586 ( .A1(n521), .A2(n525), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n522), .B(G99GAT), .ZN(G1338GAT) );
  NOR2_X1 U588 ( .A1(n524), .A2(n523), .ZN(n540) );
  NAND2_X1 U589 ( .A1(n525), .A2(n540), .ZN(n526) );
  XNOR2_X1 U590 ( .A(KEYINPUT114), .B(n526), .ZN(n527) );
  NOR2_X1 U591 ( .A1(n528), .A2(n527), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n553), .A2(n537), .ZN(n529) );
  XNOR2_X1 U593 ( .A(G113GAT), .B(n529), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n531) );
  NAND2_X1 U595 ( .A1(n537), .A2(n555), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(n533) );
  XOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT115), .Z(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  NAND2_X1 U599 ( .A1(n563), .A2(n537), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n534), .B(KEYINPUT50), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(G134GAT), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U603 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  NAND2_X1 U605 ( .A1(n565), .A2(n540), .ZN(n550) );
  NOR2_X1 U606 ( .A1(n567), .A2(n550), .ZN(n542) );
  XNOR2_X1 U607 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(G1344GAT) );
  INV_X1 U609 ( .A(n555), .ZN(n543) );
  NOR2_X1 U610 ( .A1(n543), .A2(n550), .ZN(n548) );
  XOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n545) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U614 ( .A(KEYINPUT118), .B(n546), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NOR2_X1 U616 ( .A1(n575), .A2(n550), .ZN(n549) );
  XOR2_X1 U617 ( .A(G155GAT), .B(n549), .Z(G1346GAT) );
  NOR2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U619 ( .A(G162GAT), .B(n552), .Z(G1347GAT) );
  NAND2_X1 U620 ( .A1(n553), .A2(n562), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G169GAT), .B(n554), .ZN(G1348GAT) );
  NAND2_X1 U622 ( .A1(n555), .A2(n562), .ZN(n561) );
  XOR2_X1 U623 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n557) );
  XNOR2_X1 U624 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(n559) );
  XOR2_X1 U626 ( .A(G176GAT), .B(KEYINPUT122), .Z(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(G1349GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n569) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n579) );
  OR2_X1 U633 ( .A1(n579), .A2(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n573) );
  OR2_X1 U637 ( .A1(n579), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U639 ( .A(G204GAT), .B(n574), .Z(G1353GAT) );
  OR2_X1 U640 ( .A1(n579), .A2(n575), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n578) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n582) );
  NOR2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(n582), .B(n581), .Z(G1355GAT) );
endmodule

