//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1247, new_n1248,
    new_n1249, new_n1251, new_n1252, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1325, new_n1326;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n207), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  OR2_X1    g0016(.A1(new_n216), .A2(KEYINPUT0), .ZN(new_n217));
  INV_X1    g0017(.A(G50), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n206), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(new_n211), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n216), .A2(KEYINPUT0), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n217), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT65), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(KEYINPUT66), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n228), .A2(KEYINPUT66), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n213), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n234), .A2(KEYINPUT1), .ZN(new_n235));
  AND2_X1   g0035(.A1(new_n234), .A2(KEYINPUT1), .ZN(new_n236));
  NOR3_X1   g0036(.A1(new_n225), .A2(new_n235), .A3(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G358));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT67), .ZN(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G68), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n220), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT8), .A2(G58), .ZN(new_n256));
  OR2_X1    g0056(.A1(KEYINPUT68), .A2(G58), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT68), .A2(G58), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n256), .B1(new_n259), .B2(KEYINPUT8), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G150), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT69), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(new_n211), .A3(new_n262), .ZN(new_n267));
  OAI21_X1  g0067(.A(KEYINPUT69), .B1(G20), .B2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  OAI22_X1  g0070(.A1(new_n261), .A2(new_n264), .B1(new_n265), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n211), .B1(new_n206), .B2(new_n218), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n255), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n218), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n255), .ZN(new_n277));
  OR2_X1    g0077(.A1(new_n277), .A2(KEYINPUT70), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(KEYINPUT70), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n210), .A2(G20), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n273), .B(new_n276), .C1(new_n218), .C2(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT3), .B(G33), .ZN(new_n283));
  INV_X1    g0083(.A(G1698), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(G222), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G77), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n283), .A2(G1698), .ZN(new_n287));
  INV_X1    g0087(.A(G223), .ZN(new_n288));
  OAI221_X1 g0088(.A(new_n285), .B1(new_n286), .B2(new_n283), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(G1), .A3(G13), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G41), .ZN(new_n294));
  INV_X1    g0094(.A(G45), .ZN(new_n295));
  AOI21_X1  g0095(.A(G1), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n296), .A2(new_n291), .A3(G274), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n292), .A2(new_n296), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n297), .B1(G226), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n293), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G179), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n293), .A2(new_n303), .A3(new_n299), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n282), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n282), .B(KEYINPUT9), .ZN(new_n306));
  INV_X1    g0106(.A(G190), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n300), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(G200), .B2(new_n300), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT10), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n306), .A2(new_n312), .A3(new_n309), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n305), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n283), .A2(G232), .A3(G1698), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n283), .A2(G226), .A3(new_n284), .ZN(new_n316));
  INV_X1    g0116(.A(G97), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n315), .B(new_n316), .C1(new_n262), .C2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n292), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n297), .B1(G238), .B2(new_n298), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT13), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT13), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n319), .A2(new_n323), .A3(new_n320), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G200), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n270), .A2(new_n218), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n264), .A2(new_n286), .B1(new_n211), .B2(G68), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n255), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT11), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI211_X1 g0131(.A(KEYINPUT11), .B(new_n255), .C1(new_n327), .C2(new_n328), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT74), .B1(new_n274), .B2(G68), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT12), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n333), .B(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n277), .A2(G68), .A3(new_n280), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n331), .B(new_n332), .C1(KEYINPUT75), .C2(new_n337), .ZN(new_n338));
  AND2_X1   g0138(.A1(new_n337), .A2(KEYINPUT75), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n322), .A2(G190), .A3(new_n324), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n326), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n325), .A2(G169), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT14), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n322), .A2(G179), .A3(new_n324), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT14), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n325), .A2(new_n347), .A3(G169), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n345), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n340), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n343), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G87), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT15), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT15), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G87), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n356), .A2(new_n263), .B1(G20), .B2(G77), .ZN(new_n357));
  AND2_X1   g0157(.A1(KEYINPUT8), .A2(G58), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(new_n256), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n269), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n255), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n280), .A2(G77), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n277), .A2(new_n364), .B1(new_n286), .B2(new_n275), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n362), .A2(KEYINPUT71), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT71), .ZN(new_n367));
  INV_X1    g0167(.A(new_n255), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n357), .B2(new_n360), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n274), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n370), .A2(new_n363), .B1(G77), .B2(new_n274), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n367), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n366), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n283), .A2(G232), .A3(new_n284), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n283), .A2(G238), .A3(G1698), .ZN(new_n375));
  INV_X1    g0175(.A(G107), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n374), .B(new_n375), .C1(new_n376), .C2(new_n283), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n292), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n297), .B1(G244), .B2(new_n298), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n301), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n378), .A2(new_n303), .A3(new_n379), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n373), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT72), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n366), .A2(new_n372), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n380), .A2(G200), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n384), .B1(new_n366), .B2(new_n372), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT73), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n373), .A2(KEYINPUT72), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT73), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n390), .A2(new_n391), .A3(new_n385), .A4(new_n386), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n378), .A2(G190), .A3(new_n379), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n389), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AND4_X1   g0194(.A1(new_n314), .A2(new_n351), .A3(new_n383), .A4(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT17), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT3), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(G33), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n397), .A2(new_n399), .A3(G226), .A4(G1698), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n397), .A2(new_n399), .A3(G223), .A4(new_n284), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n400), .B(new_n401), .C1(new_n262), .C2(new_n352), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n292), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n291), .A2(G274), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n298), .A2(G232), .B1(new_n404), .B2(new_n296), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n406), .A2(G190), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT76), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n403), .A2(new_n405), .A3(KEYINPUT76), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G200), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n407), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT16), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n202), .B1(new_n257), .B2(new_n258), .ZN(new_n415));
  OAI21_X1  g0215(.A(G20), .B1(new_n415), .B2(new_n206), .ZN(new_n416));
  INV_X1    g0216(.A(G159), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n416), .B1(new_n417), .B2(new_n270), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT7), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n283), .B2(G20), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n397), .A2(new_n399), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n421), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n202), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n414), .B1(new_n418), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n420), .A2(new_n422), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(G68), .ZN(new_n426));
  AND2_X1   g0226(.A1(KEYINPUT68), .A2(G58), .ZN(new_n427));
  NOR2_X1   g0227(.A1(KEYINPUT68), .A2(G58), .ZN(new_n428));
  OAI21_X1  g0228(.A(G68), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n429), .A2(new_n205), .A3(new_n203), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n430), .A2(G20), .B1(G159), .B2(new_n269), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n426), .A2(new_n431), .A3(KEYINPUT16), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n424), .A2(new_n255), .A3(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n278), .A2(new_n279), .A3(new_n280), .A4(new_n260), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n261), .A2(new_n275), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n396), .B1(new_n413), .B2(new_n438), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n403), .A2(new_n405), .A3(KEYINPUT76), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT76), .B1(new_n403), .B2(new_n405), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n301), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n406), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n303), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n426), .A2(new_n431), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n368), .B1(new_n446), .B2(new_n414), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n436), .B1(new_n447), .B2(new_n432), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT18), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT18), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n438), .A2(new_n450), .A3(new_n444), .A4(new_n442), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n412), .B1(new_n440), .B2(new_n441), .ZN(new_n452));
  INV_X1    g0252(.A(new_n407), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n454), .A2(new_n448), .A3(KEYINPUT17), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n439), .A2(new_n449), .A3(new_n451), .A4(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT77), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OR2_X1    g0258(.A1(new_n456), .A2(new_n457), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n395), .A2(KEYINPUT78), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT78), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n314), .A2(new_n351), .A3(new_n383), .A4(new_n394), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n459), .A2(new_n458), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT87), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n397), .A2(new_n399), .A3(new_n211), .A4(G87), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT22), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT22), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n283), .A2(new_n469), .A3(new_n211), .A4(G87), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT24), .ZN(new_n472));
  NAND2_X1  g0272(.A1(G33), .A2(G116), .ZN(new_n473));
  OR3_X1    g0273(.A1(new_n473), .A2(KEYINPUT84), .A3(G20), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT23), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(new_n211), .B2(G107), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n376), .A2(KEYINPUT23), .A3(G20), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT84), .B1(new_n473), .B2(G20), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n474), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n471), .A2(new_n472), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n472), .B1(new_n471), .B2(new_n480), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n255), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n210), .A2(G33), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n274), .A2(new_n484), .A3(new_n220), .A4(new_n254), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n275), .A2(KEYINPUT25), .A3(new_n376), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT25), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n274), .B2(G107), .ZN(new_n489));
  AOI22_X1  g0289(.A1(G107), .A2(new_n486), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT5), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(G41), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n210), .B(G45), .C1(new_n294), .C2(KEYINPUT5), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT79), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n491), .A2(G41), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n496), .A2(KEYINPUT79), .A3(new_n210), .A4(G45), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n404), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n493), .A2(new_n494), .ZN(new_n499));
  INV_X1    g0299(.A(new_n492), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n499), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n501), .A2(G264), .A3(new_n291), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n397), .A2(new_n399), .A3(G257), .A4(G1698), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n397), .A2(new_n399), .A3(G250), .A4(new_n284), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G294), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n292), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n502), .A2(KEYINPUT86), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT86), .B1(new_n502), .B2(new_n507), .ZN(new_n509));
  OAI211_X1 g0309(.A(G179), .B(new_n498), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT85), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n502), .B(new_n498), .C1(new_n507), .C2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT85), .B1(new_n506), .B2(new_n292), .ZN(new_n513));
  OAI21_X1  g0313(.A(G169), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI221_X4 g0314(.A(new_n466), .B1(new_n483), .B2(new_n490), .C1(new_n510), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n510), .A2(new_n514), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n483), .A2(new_n490), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT87), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n517), .ZN(new_n520));
  INV_X1    g0320(.A(new_n498), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n502), .A2(new_n507), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT86), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n502), .A2(new_n507), .A3(KEYINPUT86), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n521), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n526), .A2(G200), .ZN(new_n527));
  NOR3_X1   g0327(.A1(new_n512), .A2(new_n513), .A3(G190), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n520), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AND2_X1   g0329(.A1(new_n519), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G283), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n397), .A2(new_n399), .A3(G250), .A4(G1698), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n397), .A2(new_n399), .A3(G244), .A4(new_n284), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT4), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n531), .B(new_n532), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n292), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n501), .A2(G257), .A3(new_n291), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n498), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT6), .ZN(new_n540));
  NOR3_X1   g0340(.A1(new_n540), .A2(new_n317), .A3(G107), .ZN(new_n541));
  XNOR2_X1  g0341(.A(G97), .B(G107), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n541), .B1(new_n542), .B2(new_n540), .ZN(new_n543));
  OAI22_X1  g0343(.A1(new_n543), .A2(new_n211), .B1(new_n286), .B2(new_n270), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n376), .B1(new_n420), .B2(new_n422), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n255), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n274), .A2(G97), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n547), .B1(new_n486), .B2(G97), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n539), .A2(new_n301), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT80), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n538), .A2(new_n550), .A3(new_n498), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n550), .B1(new_n538), .B2(new_n498), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n303), .B(new_n537), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n537), .ZN(new_n555));
  INV_X1    g0355(.A(G257), .ZN(new_n556));
  AOI211_X1 g0356(.A(new_n556), .B(new_n292), .C1(new_n495), .C2(new_n497), .ZN(new_n557));
  OAI21_X1  g0357(.A(KEYINPUT80), .B1(new_n557), .B2(new_n521), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n538), .A2(new_n550), .A3(new_n498), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n555), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n560), .A2(new_n412), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n546), .B(new_n548), .C1(new_n539), .C2(new_n307), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n554), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n486), .A2(G116), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n531), .B(new_n211), .C1(G33), .C2(new_n317), .ZN(new_n565));
  INV_X1    g0365(.A(G116), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G20), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n565), .A2(new_n255), .A3(new_n567), .ZN(new_n568));
  XOR2_X1   g0368(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n275), .A2(new_n566), .ZN(new_n571));
  NOR2_X1   g0371(.A1(KEYINPUT83), .A2(KEYINPUT20), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n565), .A2(new_n255), .A3(new_n567), .A4(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n564), .A2(new_n570), .A3(new_n571), .A4(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n501), .A2(G270), .A3(new_n291), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n398), .A2(G33), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n577));
  OAI21_X1  g0377(.A(G303), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n397), .A2(new_n399), .A3(G264), .A4(G1698), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n397), .A2(new_n399), .A3(G257), .A4(new_n284), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n292), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n575), .A2(new_n582), .A3(new_n498), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n574), .B1(new_n583), .B2(G200), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n307), .B2(new_n583), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n583), .A2(G169), .A3(new_n574), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT21), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n303), .B1(new_n581), .B2(new_n292), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n574), .A2(new_n589), .A3(new_n498), .A4(new_n575), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n583), .A2(KEYINPUT21), .A3(G169), .A4(new_n574), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n585), .A2(new_n588), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n356), .A2(new_n274), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n485), .A2(new_n352), .ZN(new_n594));
  XNOR2_X1  g0394(.A(KEYINPUT82), .B(G87), .ZN(new_n595));
  NOR2_X1   g0395(.A1(G97), .A2(G107), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n211), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n283), .A2(new_n211), .A3(G68), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT19), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n264), .B2(new_n317), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  AOI211_X1 g0404(.A(new_n593), .B(new_n594), .C1(new_n604), .C2(new_n255), .ZN(new_n605));
  INV_X1    g0405(.A(G250), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n295), .B2(G1), .ZN(new_n607));
  INV_X1    g0407(.A(G274), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n210), .A2(new_n608), .A3(G45), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n291), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n397), .A2(new_n399), .A3(G238), .A4(new_n284), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n397), .A2(new_n399), .A3(G244), .A4(G1698), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(new_n613), .A3(new_n473), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n611), .B1(new_n614), .B2(new_n292), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G190), .ZN(new_n616));
  INV_X1    g0416(.A(new_n615), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G200), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n605), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n615), .A2(new_n303), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT81), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n604), .A2(new_n255), .ZN(new_n623));
  INV_X1    g0423(.A(new_n593), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n486), .A2(new_n356), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n617), .A2(new_n301), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n622), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n620), .A2(new_n621), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n619), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n563), .A2(new_n592), .A3(new_n630), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n465), .A2(new_n530), .A3(new_n631), .ZN(G372));
  NAND3_X1  g0432(.A1(new_n626), .A2(new_n620), .A3(new_n627), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n619), .A2(new_n633), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n554), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT26), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(KEYINPUT26), .B1(new_n630), .B2(new_n554), .ZN(new_n639));
  INV_X1    g0439(.A(new_n562), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n537), .B1(new_n551), .B2(new_n552), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(G200), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n640), .A2(new_n642), .B1(new_n553), .B2(new_n549), .ZN(new_n643));
  INV_X1    g0443(.A(new_n635), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n529), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n516), .A2(new_n517), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n638), .B(new_n639), .C1(new_n645), .C2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n465), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n449), .A2(new_n451), .ZN(new_n651));
  INV_X1    g0451(.A(new_n383), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n349), .A2(new_n350), .B1(new_n342), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n439), .A2(new_n455), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n651), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n311), .A2(new_n313), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n305), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n650), .A2(new_n657), .ZN(G369));
  NAND3_X1  g0458(.A1(new_n210), .A2(new_n211), .A3(G13), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(G213), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G343), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n530), .B1(new_n520), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n516), .A2(new_n517), .A3(new_n664), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n647), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n574), .A2(new_n664), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n592), .B2(new_n670), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(G330), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n668), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n664), .B(KEYINPUT88), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n516), .A2(new_n517), .A3(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n647), .A2(new_n664), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n519), .A2(new_n529), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n675), .A2(new_n677), .A3(new_n679), .ZN(G399));
  INV_X1    g0480(.A(new_n214), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(G41), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n597), .A2(G116), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G1), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n219), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n685), .B1(new_n686), .B2(new_n683), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT28), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n649), .A2(new_n676), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n689), .A2(KEYINPUT29), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n646), .A2(new_n466), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT87), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(new_n692), .A3(new_n647), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n693), .A2(new_n529), .A3(new_n643), .A4(new_n644), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n636), .A2(new_n637), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n630), .A2(new_n554), .A3(KEYINPUT26), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n633), .B(KEYINPUT92), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n664), .B1(new_n694), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT29), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n690), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT31), .ZN(new_n702));
  XNOR2_X1  g0502(.A(KEYINPUT89), .B(KEYINPUT30), .ZN(new_n703));
  AND4_X1   g0503(.A1(new_n498), .A2(new_n589), .A3(new_n615), .A4(new_n575), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n537), .A2(new_n498), .A3(new_n538), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n508), .A2(new_n509), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n703), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n589), .A2(new_n615), .A3(new_n498), .A4(new_n575), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(new_n539), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT30), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n524), .A2(new_n525), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n526), .A2(new_n560), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n614), .A2(new_n292), .ZN(new_n715));
  AOI21_X1  g0515(.A(G179), .B1(new_n715), .B2(new_n610), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n583), .A2(new_n716), .A3(KEYINPUT90), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT90), .B1(new_n583), .B2(new_n716), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI22_X1  g0519(.A1(new_n708), .A2(new_n713), .B1(new_n714), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n664), .B1(new_n720), .B2(KEYINPUT91), .ZN(new_n721));
  INV_X1    g0521(.A(new_n718), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n498), .B1(new_n508), .B2(new_n509), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n583), .A2(new_n716), .A3(KEYINPUT90), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n722), .A2(new_n723), .A3(new_n641), .A4(new_n724), .ZN(new_n725));
  NOR4_X1   g0525(.A1(new_n707), .A2(KEYINPUT30), .A3(new_n539), .A4(new_n709), .ZN(new_n726));
  INV_X1    g0526(.A(new_n703), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n727), .B1(new_n710), .B2(new_n712), .ZN(new_n728));
  OAI211_X1 g0528(.A(KEYINPUT91), .B(new_n725), .C1(new_n726), .C2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n702), .B1(new_n721), .B2(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n631), .A2(new_n519), .A3(new_n529), .A4(new_n676), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n725), .B1(new_n726), .B2(new_n728), .ZN(new_n733));
  INV_X1    g0533(.A(new_n676), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(KEYINPUT31), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n731), .A2(new_n732), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G330), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n701), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n688), .B1(new_n739), .B2(G1), .ZN(G364));
  INV_X1    g0540(.A(G13), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G20), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n210), .B1(new_n742), .B2(G45), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n682), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n214), .A2(new_n283), .ZN(new_n746));
  INV_X1    g0546(.A(G355), .ZN(new_n747));
  OAI22_X1  g0547(.A1(new_n746), .A2(new_n747), .B1(G116), .B2(new_n214), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n681), .A2(new_n283), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n750), .B1(new_n219), .B2(new_n295), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n252), .A2(G45), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n748), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n220), .B1(G20), .B2(new_n301), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n745), .B1(new_n753), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n211), .A2(new_n303), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n761), .A2(new_n307), .A3(new_n412), .ZN(new_n762));
  NOR4_X1   g0562(.A1(new_n211), .A2(new_n303), .A3(new_n412), .A4(G190), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n283), .B1(new_n286), .B2(new_n762), .C1(new_n764), .C2(new_n202), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n761), .A2(G190), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n412), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G179), .A2(G200), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n211), .B1(new_n769), .B2(G190), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n768), .A2(new_n218), .B1(new_n770), .B2(new_n317), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n765), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n766), .A2(G200), .ZN(new_n773));
  NOR4_X1   g0573(.A1(new_n211), .A2(new_n412), .A3(G179), .A4(G190), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n773), .A2(new_n259), .B1(G107), .B2(new_n774), .ZN(new_n775));
  NOR4_X1   g0575(.A1(new_n211), .A2(new_n307), .A3(new_n412), .A4(G179), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n772), .B(new_n775), .C1(new_n595), .C2(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n769), .A2(G20), .A3(new_n307), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT93), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n779), .A2(new_n780), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G159), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT32), .ZN(new_n786));
  INV_X1    g0586(.A(G311), .ZN(new_n787));
  XOR2_X1   g0587(.A(KEYINPUT33), .B(G317), .Z(new_n788));
  OAI221_X1 g0588(.A(new_n421), .B1(new_n787), .B2(new_n762), .C1(new_n764), .C2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n774), .ZN(new_n790));
  INV_X1    g0590(.A(G283), .ZN(new_n791));
  INV_X1    g0591(.A(G294), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n790), .A2(new_n791), .B1(new_n792), .B2(new_n770), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n767), .A2(G326), .B1(G303), .B2(new_n776), .ZN(new_n795));
  INV_X1    g0595(.A(G322), .ZN(new_n796));
  INV_X1    g0596(.A(new_n773), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n794), .B(new_n795), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n783), .B(KEYINPUT94), .ZN(new_n799));
  INV_X1    g0599(.A(G329), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n778), .A2(new_n786), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n760), .B1(new_n802), .B2(new_n757), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n756), .B(KEYINPUT95), .Z(new_n804));
  OAI21_X1  g0604(.A(new_n803), .B1(new_n672), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n745), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n673), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n672), .A2(G330), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(G396));
  INV_X1    g0609(.A(G303), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n768), .A2(new_n810), .B1(new_n376), .B2(new_n777), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n797), .A2(new_n792), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n421), .B1(new_n770), .B2(new_n317), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n790), .A2(new_n352), .ZN(new_n814));
  NOR4_X1   g0614(.A1(new_n811), .A2(new_n812), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n762), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n816), .A2(G116), .B1(new_n763), .B2(G283), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT96), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n815), .B(new_n818), .C1(new_n787), .C2(new_n799), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n816), .A2(G159), .B1(new_n763), .B2(G150), .ZN(new_n820));
  INV_X1    g0620(.A(G143), .ZN(new_n821));
  INV_X1    g0621(.A(G137), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n820), .B1(new_n797), .B2(new_n821), .C1(new_n822), .C2(new_n768), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n823), .B(KEYINPUT34), .Z(new_n824));
  AOI21_X1  g0624(.A(new_n421), .B1(new_n776), .B2(G50), .ZN(new_n825));
  INV_X1    g0625(.A(new_n770), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n826), .A2(new_n259), .B1(new_n774), .B2(G68), .ZN(new_n827));
  INV_X1    g0627(.A(G132), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n825), .B(new_n827), .C1(new_n799), .C2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n819), .B1(new_n824), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n757), .A2(new_n754), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n830), .A2(new_n757), .B1(new_n286), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n383), .A2(new_n664), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n373), .A2(new_n664), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n394), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n833), .B1(new_n835), .B2(new_n383), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n832), .B1(new_n836), .B2(new_n755), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n745), .ZN(new_n838));
  INV_X1    g0638(.A(new_n836), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n689), .B(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n737), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n806), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n840), .A2(new_n737), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n838), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT97), .Z(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(G384));
  NOR2_X1   g0646(.A1(new_n742), .A2(new_n210), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT100), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT91), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n733), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n850), .A2(KEYINPUT31), .A3(new_n664), .A4(new_n729), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n732), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT99), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n731), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n850), .A2(new_n664), .A3(new_n729), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n855), .A2(KEYINPUT99), .A3(new_n702), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n852), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n350), .B(new_n664), .C1(new_n349), .C2(new_n343), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n348), .A2(new_n346), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n347), .B1(new_n325), .B2(G169), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n350), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n350), .A2(new_n664), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n861), .A2(new_n342), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n836), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n848), .B1(new_n857), .B2(new_n865), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n732), .A2(new_n851), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n665), .B1(new_n733), .B2(new_n849), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n853), .B(KEYINPUT31), .C1(new_n868), .C2(new_n729), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT99), .B1(new_n855), .B2(new_n702), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n867), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n865), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n871), .A2(KEYINPUT100), .A3(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT40), .ZN(new_n874));
  INV_X1    g0674(.A(new_n662), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n438), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n456), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n448), .B1(new_n445), .B2(new_n662), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n413), .A2(new_n438), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT37), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n454), .A2(new_n448), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n438), .A2(new_n444), .A3(new_n442), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT37), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n882), .A2(new_n883), .A3(new_n884), .A4(new_n876), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n878), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT38), .ZN(new_n888));
  INV_X1    g0688(.A(new_n885), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n411), .A2(new_n301), .B1(new_n303), .B2(new_n443), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n438), .B1(new_n890), .B2(new_n875), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n884), .B1(new_n891), .B2(new_n882), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT98), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n887), .A2(new_n888), .A3(new_n893), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n878), .B(new_n886), .C1(KEYINPUT98), .C2(KEYINPUT38), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n874), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n866), .A2(new_n873), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n878), .A2(new_n886), .A3(new_n888), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n888), .B1(new_n878), .B2(new_n886), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n871), .A2(new_n901), .A3(new_n872), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n897), .B1(KEYINPUT40), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n465), .A2(new_n871), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  INV_X1    g0707(.A(G330), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n701), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n465), .A2(new_n911), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n912), .A2(new_n657), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT39), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n887), .A2(new_n888), .A3(new_n893), .ZN(new_n915));
  INV_X1    g0715(.A(new_n895), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n887), .A2(KEYINPUT38), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n914), .B1(new_n918), .B2(new_n898), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n349), .A2(new_n350), .A3(new_n665), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n858), .A2(new_n863), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n649), .A2(new_n836), .A3(new_n676), .ZN(new_n925));
  INV_X1    g0725(.A(new_n833), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n901), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n651), .B2(new_n875), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n923), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n913), .B(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n847), .B1(new_n910), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n931), .B2(new_n910), .ZN(new_n933));
  INV_X1    g0733(.A(new_n543), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n934), .A2(KEYINPUT35), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(KEYINPUT35), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n935), .A2(G116), .A3(new_n221), .A4(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT36), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n219), .A2(G77), .A3(new_n429), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(G50), .B2(new_n202), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n940), .A2(G1), .A3(new_n741), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n933), .A2(new_n938), .A3(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT101), .Z(G367));
  OAI21_X1  g0743(.A(new_n679), .B1(new_n668), .B2(new_n678), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(new_n673), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n945), .A2(new_n738), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT44), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n679), .A2(new_n677), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n546), .A2(new_n548), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n643), .B1(new_n949), .B2(new_n676), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n734), .A2(new_n549), .A3(new_n553), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n948), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT104), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n954), .A2(KEYINPUT104), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n947), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n954), .A2(KEYINPUT104), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n959), .A2(KEYINPUT44), .A3(new_n955), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n948), .A2(new_n953), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT45), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n958), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT105), .ZN(new_n964));
  INV_X1    g0764(.A(new_n675), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n958), .A2(new_n960), .A3(new_n675), .A4(new_n962), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n946), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n964), .B1(new_n963), .B2(new_n965), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n739), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n682), .B(KEYINPUT41), .Z(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n744), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n530), .A2(new_n678), .A3(new_n952), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(KEYINPUT42), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT103), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n561), .A2(new_n562), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n554), .B1(new_n519), .B2(new_n977), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n974), .A2(KEYINPUT42), .B1(new_n676), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n605), .A2(new_n665), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n634), .A2(new_n981), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n982), .A2(KEYINPUT102), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n982), .B(KEYINPUT102), .C1(new_n635), .C2(new_n981), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n980), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT43), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n976), .A2(new_n991), .A3(new_n985), .A4(new_n979), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n675), .A2(new_n953), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n994), .B1(new_n990), .B2(new_n992), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(KEYINPUT106), .B1(new_n973), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT106), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n969), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n1002), .A2(new_n966), .A3(new_n946), .A4(new_n967), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n971), .B1(new_n1003), .B2(new_n739), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n998), .B(new_n1001), .C1(new_n1004), .C2(new_n744), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1000), .A2(new_n1005), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n773), .A2(G150), .B1(G68), .B2(new_n826), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT107), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n259), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n768), .A2(new_n821), .B1(new_n1009), .B2(new_n777), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n790), .A2(new_n286), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n1010), .A2(new_n421), .A3(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n816), .A2(G50), .B1(new_n763), .B2(G159), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT108), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n784), .A2(G137), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1008), .A2(new_n1012), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT109), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n790), .A2(new_n317), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n768), .A2(new_n787), .B1(new_n770), .B2(new_n376), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n1018), .B(new_n1019), .C1(G303), .C2(new_n773), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n784), .A2(G317), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n421), .B1(new_n762), .B2(new_n791), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G294), .B2(new_n763), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n776), .A2(G116), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT46), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1020), .A2(new_n1021), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1017), .A2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT47), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n757), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n749), .A2(new_n244), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n759), .B1(new_n681), .B2(new_n356), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n806), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1029), .B(new_n1032), .C1(new_n804), .C2(new_n986), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1006), .A2(new_n1033), .ZN(G387));
  INV_X1    g0834(.A(new_n945), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n668), .A2(new_n804), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n749), .B1(new_n241), .B2(new_n295), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n684), .B2(new_n746), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n359), .A2(new_n218), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT50), .Z(new_n1040));
  AOI21_X1  g0840(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1040), .A2(new_n684), .A3(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n1038), .A2(new_n1042), .B1(new_n376), .B2(new_n681), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n745), .B1(new_n1043), .B2(new_n759), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT110), .Z(new_n1045));
  OAI22_X1  g0845(.A1(new_n261), .A2(new_n764), .B1(new_n202), .B2(new_n762), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT111), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n797), .A2(new_n218), .B1(new_n768), .B2(new_n417), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n356), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1049), .A2(new_n770), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n777), .A2(new_n286), .ZN(new_n1051));
  NOR3_X1   g0851(.A1(new_n1048), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n421), .B(new_n1018), .C1(new_n784), .C2(G150), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1047), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n816), .A2(G303), .B1(new_n763), .B2(G311), .ZN(new_n1055));
  INV_X1    g0855(.A(G317), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1055), .B1(new_n797), .B2(new_n1056), .C1(new_n796), .C2(new_n768), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT112), .Z(new_n1058));
  INV_X1    g0858(.A(KEYINPUT48), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n777), .A2(new_n792), .B1(new_n791), .B2(new_n770), .ZN(new_n1062));
  NOR3_X1   g0862(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(KEYINPUT49), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n784), .A2(G326), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n283), .B1(new_n774), .B2(G116), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1063), .A2(KEYINPUT49), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1054), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1069), .A2(KEYINPUT113), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n757), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n1069), .B2(KEYINPUT113), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1045), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1035), .A2(new_n744), .B1(new_n1036), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n946), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n682), .B(KEYINPUT114), .Z(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1035), .A2(new_n739), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1074), .B1(new_n1077), .B2(new_n1078), .ZN(G393));
  NOR2_X1   g0879(.A1(new_n249), .A2(new_n750), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n758), .B1(new_n317), .B2(new_n214), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n745), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(G311), .A2(new_n773), .B1(new_n767), .B2(G317), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT52), .Z(new_n1084));
  NAND2_X1  g0884(.A1(new_n826), .A2(G116), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n816), .A2(G294), .B1(new_n763), .B2(G303), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n283), .B1(new_n774), .B2(G107), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1088), .B1(new_n791), .B2(new_n777), .C1(new_n783), .C2(new_n796), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT115), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G150), .A2(new_n767), .B1(new_n773), .B2(G159), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT51), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n764), .A2(new_n218), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n421), .B(new_n1093), .C1(new_n359), .C2(new_n816), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n770), .A2(new_n286), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1095), .B(new_n814), .C1(G68), .C2(new_n776), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1094), .B(new_n1096), .C1(new_n821), .C2(new_n783), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n1087), .A2(new_n1090), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1082), .B1(new_n1098), .B2(new_n757), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n756), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1099), .B1(new_n952), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n963), .A2(new_n965), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n967), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1101), .B1(new_n1103), .B2(new_n743), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1076), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n1075), .B2(new_n1103), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1104), .B1(new_n1003), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(G390));
  OAI22_X1  g0908(.A1(new_n768), .A2(new_n791), .B1(new_n202), .B2(new_n790), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n421), .B1(new_n317), .B2(new_n762), .C1(new_n764), .C2(new_n376), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1109), .B(new_n1110), .C1(G87), .C2(new_n776), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1095), .B1(new_n773), .B2(G116), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT117), .Z(new_n1113));
  OAI211_X1 g0913(.A(new_n1111), .B(new_n1113), .C1(new_n792), .C2(new_n799), .ZN(new_n1114));
  INV_X1    g0914(.A(G128), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n797), .A2(new_n828), .B1(new_n768), .B2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT54), .B(G143), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n283), .B1(new_n762), .B2(new_n1117), .C1(new_n764), .C2(new_n822), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n790), .A2(new_n218), .B1(new_n417), .B2(new_n770), .ZN(new_n1119));
  NOR3_X1   g0919(.A1(new_n1116), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n776), .A2(G150), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT53), .Z(new_n1122));
  INV_X1    g0922(.A(G125), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1120), .B(new_n1122), .C1(new_n1123), .C2(new_n799), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1071), .B1(new_n1114), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n831), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n745), .B1(new_n260), .B2(new_n1126), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1125), .B(new_n1127), .C1(new_n921), .C2(new_n754), .ZN(new_n1128));
  AOI21_X1  g0928(.A(KEYINPUT39), .B1(new_n894), .B2(new_n895), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n922), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n1129), .A2(new_n919), .B1(new_n927), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1130), .B1(new_n894), .B2(new_n895), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n835), .A2(new_n383), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n833), .B1(new_n699), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1132), .B1(new_n1134), .B2(new_n924), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n736), .A2(G330), .A3(new_n836), .A4(new_n864), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1131), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n871), .A2(G330), .A3(new_n872), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1128), .B1(new_n1140), .B2(new_n744), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n857), .A2(new_n908), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n465), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n912), .A2(new_n1143), .A3(new_n657), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n924), .B1(new_n737), .B2(new_n839), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n1138), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n925), .A2(new_n926), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n871), .A2(G330), .A3(new_n836), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1150), .A2(KEYINPUT116), .A3(new_n924), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1136), .A2(new_n1134), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(KEYINPUT116), .B1(new_n1150), .B2(new_n924), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1149), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1145), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1140), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1076), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1140), .B1(new_n1145), .B2(new_n1155), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1141), .B1(new_n1158), .B2(new_n1159), .ZN(G378));
  AOI21_X1  g0960(.A(new_n908), .B1(new_n902), .B2(new_n874), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n282), .A2(new_n875), .ZN(new_n1162));
  OR2_X1    g0962(.A1(new_n314), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n314), .A2(new_n1162), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1165), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n897), .A2(new_n1161), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1168), .B1(new_n897), .B2(new_n1161), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n930), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n897), .A2(new_n1161), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1168), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n928), .B1(new_n651), .B2(new_n875), .C1(new_n921), .C2(new_n922), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n897), .A2(new_n1161), .A3(new_n1168), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1171), .A2(new_n1177), .A3(KEYINPUT120), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT120), .B1(new_n1171), .B2(new_n1177), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n744), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1168), .A2(new_n754), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n745), .B1(G50), .B2(new_n1126), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT119), .ZN(new_n1183));
  NOR3_X1   g0983(.A1(new_n1051), .A2(G41), .A3(new_n283), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n1009), .B2(new_n790), .C1(new_n799), .C2(new_n791), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT118), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n764), .A2(new_n317), .B1(new_n1049), .B2(new_n762), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(G68), .B2(new_n826), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(G107), .A2(new_n773), .B1(new_n767), .B2(G116), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1186), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT58), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(G33), .A2(G41), .ZN(new_n1194));
  AOI211_X1 g0994(.A(G50), .B(new_n1194), .C1(new_n421), .C2(new_n294), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n764), .A2(new_n828), .B1(new_n762), .B2(new_n822), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1117), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1196), .B1(new_n776), .B2(new_n1197), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n767), .A2(G125), .B1(G150), .B2(new_n826), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1198), .B(new_n1199), .C1(new_n1115), .C2(new_n797), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1201));
  INV_X1    g1001(.A(G124), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1194), .B1(new_n417), .B2(new_n790), .C1(new_n783), .C2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n1200), .B2(KEYINPUT59), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1195), .B1(new_n1201), .B2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1192), .A2(new_n1193), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1183), .B1(new_n1206), .B2(new_n757), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1181), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1180), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1144), .B1(new_n1155), .B2(new_n1140), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT57), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1210), .A2(new_n1213), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1175), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(KEYINPUT121), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT121), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1171), .A2(new_n1177), .A3(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1215), .A2(new_n1217), .A3(new_n1219), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n1220), .A2(new_n1076), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1209), .B1(new_n1214), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(G375));
  INV_X1    g1023(.A(new_n1155), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n1144), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1225), .A2(new_n972), .A3(new_n1156), .ZN(new_n1226));
  XOR2_X1   g1026(.A(new_n743), .B(KEYINPUT122), .Z(new_n1227));
  NAND2_X1  g1027(.A1(new_n924), .A2(new_n754), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n745), .B1(G68), .B2(new_n1126), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1229), .B(KEYINPUT123), .Z(new_n1230));
  AOI22_X1  g1030(.A1(new_n767), .A2(G294), .B1(G97), .B2(new_n776), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n791), .B2(new_n797), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n421), .B1(new_n376), .B2(new_n762), .C1(new_n764), .C2(new_n566), .ZN(new_n1233));
  NOR4_X1   g1033(.A1(new_n1232), .A2(new_n1233), .A3(new_n1011), .A4(new_n1050), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n810), .B2(new_n799), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n283), .B1(new_n762), .B2(new_n265), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n259), .B2(new_n774), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n776), .A2(G159), .B1(new_n826), .B2(G50), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1237), .B(new_n1238), .C1(new_n799), .C2(new_n1115), .ZN(new_n1239));
  XOR2_X1   g1039(.A(new_n1239), .B(KEYINPUT124), .Z(new_n1240));
  AOI22_X1  g1040(.A1(new_n767), .A2(G132), .B1(new_n763), .B2(new_n1197), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n822), .B2(new_n797), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1235), .B1(new_n1240), .B2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1230), .B1(new_n1243), .B2(new_n757), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1155), .A2(new_n1227), .B1(new_n1228), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1226), .A2(new_n1245), .ZN(G381));
  NOR3_X1   g1046(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1107), .ZN(new_n1248));
  NOR4_X1   g1048(.A1(G387), .A2(G378), .A3(new_n1248), .A4(G381), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1222), .ZN(G407));
  INV_X1    g1050(.A(G378), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1222), .A2(new_n663), .A3(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(G407), .A2(G213), .A3(new_n1252), .ZN(G409));
  INV_X1    g1053(.A(KEYINPUT126), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1219), .A2(new_n1217), .A3(new_n1227), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1255), .A2(new_n1208), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT120), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n1169), .A2(new_n1170), .A3(new_n930), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1257), .B1(new_n1258), .B2(new_n1216), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1171), .A2(new_n1177), .A3(KEYINPUT120), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1261), .A2(new_n972), .A3(new_n1211), .ZN(new_n1262));
  AOI21_X1  g1062(.A(G378), .B1(new_n1256), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT125), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n1222), .B2(G378), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1208), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(new_n1261), .B2(new_n744), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT57), .B1(new_n1261), .B2(new_n1211), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1220), .A2(new_n1076), .ZN(new_n1270));
  OAI211_X1 g1070(.A(G378), .B(new_n1268), .C1(new_n1269), .C2(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1271), .A2(KEYINPUT125), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1264), .B1(new_n1266), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(G213), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1274), .A2(G343), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT63), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT60), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1225), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1224), .A2(KEYINPUT60), .A3(new_n1144), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1279), .A2(new_n1076), .A3(new_n1156), .A4(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1245), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(G384), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1281), .A2(new_n845), .A3(new_n1245), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1277), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1273), .A2(new_n1276), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1275), .A2(G2897), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1287), .B(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1271), .A2(KEYINPUT125), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1221), .A2(new_n1214), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1292), .A2(new_n1265), .A3(G378), .A4(new_n1268), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1263), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1290), .B1(new_n1294), .B2(new_n1275), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT61), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(G387), .A2(new_n1107), .ZN(new_n1297));
  XNOR2_X1  g1097(.A(G393), .B(G396), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1006), .A2(new_n1033), .A3(G390), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1297), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(G390), .B1(new_n1006), .B2(new_n1033), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1033), .ZN(new_n1303));
  AOI211_X1 g1103(.A(new_n1303), .B(new_n1107), .C1(new_n1000), .C2(new_n1005), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1298), .B1(new_n1302), .B2(new_n1304), .ZN(new_n1305));
  AND2_X1   g1105(.A1(new_n1301), .A2(new_n1305), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1286), .A2(new_n1295), .A3(new_n1296), .A4(new_n1306), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1294), .A2(new_n1275), .ZN(new_n1308));
  AOI21_X1  g1108(.A(KEYINPUT63), .B1(new_n1308), .B2(new_n1287), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1254), .B1(new_n1307), .B2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1273), .A2(new_n1276), .ZN(new_n1311));
  AOI21_X1  g1111(.A(KEYINPUT61), .B1(new_n1311), .B2(new_n1290), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1273), .A2(new_n1276), .A3(new_n1287), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1277), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1301), .A2(new_n1305), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1315), .B1(new_n1308), .B2(new_n1285), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1312), .A2(new_n1314), .A3(new_n1316), .A4(KEYINPUT126), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1310), .A2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1313), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1312), .ZN(new_n1320));
  XNOR2_X1  g1120(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1313), .A2(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1315), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1318), .A2(new_n1323), .ZN(G405));
  OAI22_X1  g1124(.A1(new_n1266), .A2(new_n1272), .B1(G378), .B2(new_n1222), .ZN(new_n1325));
  XNOR2_X1  g1125(.A(new_n1325), .B(new_n1287), .ZN(new_n1326));
  XNOR2_X1  g1126(.A(new_n1326), .B(new_n1315), .ZN(G402));
endmodule


