//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n756, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n849,
    new_n850, new_n851, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  XOR2_X1   g001(.A(KEYINPUT69), .B(G71gat), .Z(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G99gat), .ZN(new_n204));
  XOR2_X1   g003(.A(G15gat), .B(G43gat), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(KEYINPUT24), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G183gat), .B(G190gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT24), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT23), .ZN(new_n214));
  INV_X1    g013(.A(G169gat), .ZN(new_n215));
  INV_X1    g014(.A(G176gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT25), .B1(new_n219), .B2(KEYINPUT23), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n212), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n223));
  INV_X1    g022(.A(G190gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT27), .B(G183gat), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G183gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT27), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT27), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G183gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n228), .A2(new_n230), .A3(new_n224), .A4(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(new_n207), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n226), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT64), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(G169gat), .B2(G176gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT26), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n213), .A2(new_n238), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n217), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n222), .B1(new_n234), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n235), .A2(new_n237), .A3(KEYINPUT23), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n244), .A2(new_n218), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n227), .A2(G190gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n224), .A2(G183gat), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n211), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT65), .B1(new_n248), .B2(new_n208), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n209), .B(new_n250), .C1(new_n210), .C2(new_n211), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n245), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT25), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n243), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G113gat), .B(G120gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G127gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n258), .A2(G134gat), .ZN(new_n259));
  INV_X1    g058(.A(G134gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n260), .A2(G127gat), .ZN(new_n261));
  OAI22_X1  g060(.A1(new_n255), .A2(new_n257), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G120gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(G113gat), .ZN(new_n264));
  INV_X1    g063(.A(G113gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G120gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G127gat), .B(G134gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n267), .A2(new_n268), .A3(new_n256), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n262), .A2(new_n269), .A3(KEYINPUT68), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT68), .B1(new_n262), .B2(new_n269), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n254), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G227gat), .ZN(new_n275));
  INV_X1    g074(.A(G233gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n272), .A2(new_n243), .A3(new_n253), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n274), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT33), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n206), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n277), .B1(new_n274), .B2(new_n278), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT34), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI211_X1 g083(.A(KEYINPUT34), .B(new_n277), .C1(new_n274), .C2(new_n278), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n281), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NOR3_X1   g086(.A1(new_n281), .A2(new_n284), .A3(new_n285), .ZN(new_n288));
  AND2_X1   g087(.A1(new_n279), .A2(KEYINPUT32), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NOR3_X1   g089(.A1(new_n287), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n284), .A2(new_n285), .ZN(new_n292));
  INV_X1    g091(.A(new_n281), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n289), .B1(new_n294), .B2(new_n286), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n202), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  NOR3_X1   g096(.A1(new_n291), .A2(new_n295), .A3(new_n202), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XOR2_X1   g098(.A(G1gat), .B(G29gat), .Z(new_n300));
  XNOR2_X1  g099(.A(G57gat), .B(G85gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  XOR2_X1   g103(.A(new_n304), .B(KEYINPUT85), .Z(new_n305));
  INV_X1    g104(.A(G155gat), .ZN(new_n306));
  INV_X1    g105(.A(G162gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G141gat), .B(G148gat), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n310), .B(KEYINPUT72), .C1(KEYINPUT2), .C2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT72), .ZN(new_n313));
  INV_X1    g112(.A(G148gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G141gat), .ZN(new_n315));
  INV_X1    g114(.A(G141gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(G148gat), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT2), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n308), .A2(new_n309), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n313), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n312), .A2(new_n320), .ZN(new_n321));
  XOR2_X1   g120(.A(KEYINPUT76), .B(KEYINPUT3), .Z(new_n322));
  OAI21_X1  g121(.A(new_n309), .B1(new_n308), .B2(KEYINPUT2), .ZN(new_n323));
  AND2_X1   g122(.A1(KEYINPUT73), .A2(G141gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(KEYINPUT73), .A2(G141gat), .ZN(new_n325));
  NOR3_X1   g124(.A1(new_n324), .A2(new_n325), .A3(new_n314), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT74), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n327), .B1(new_n316), .B2(G148gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n314), .A2(KEYINPUT74), .A3(G141gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OAI211_X1 g129(.A(KEYINPUT75), .B(new_n323), .C1(new_n326), .C2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT73), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n316), .ZN(new_n334));
  NAND2_X1  g133(.A1(KEYINPUT73), .A2(G141gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n334), .A2(G148gat), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n336), .A2(new_n328), .A3(new_n329), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT75), .B1(new_n337), .B2(new_n323), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n321), .B(new_n322), .C1(new_n332), .C2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n262), .A2(new_n269), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n323), .B1(new_n326), .B2(new_n330), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT75), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI22_X1  g142(.A1(new_n343), .A2(new_n331), .B1(new_n320), .B2(new_n312), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT3), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n339), .B(new_n340), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT4), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n321), .B1(new_n332), .B2(new_n338), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n347), .B1(new_n348), .B2(new_n272), .ZN(new_n349));
  INV_X1    g148(.A(new_n340), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n344), .A2(KEYINPUT4), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n346), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(G225gat), .A2(G233gat), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n305), .B1(new_n355), .B2(KEYINPUT39), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n348), .A2(new_n340), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n344), .A2(new_n350), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(KEYINPUT39), .B1(new_n359), .B2(new_n354), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n360), .B1(new_n352), .B2(new_n354), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n356), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT40), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n347), .B1(new_n273), .B2(new_n344), .ZN(new_n364));
  NOR3_X1   g163(.A1(new_n348), .A2(KEYINPUT4), .A3(new_n340), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n353), .B(new_n346), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT77), .B(KEYINPUT5), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n367), .B1(new_n359), .B2(new_n354), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  AND3_X1   g168(.A1(new_n349), .A2(new_n367), .A3(new_n351), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n350), .B1(new_n348), .B2(KEYINPUT3), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n354), .B1(new_n371), .B2(new_n339), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n305), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n363), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n362), .A2(KEYINPUT40), .ZN(new_n378));
  OR2_X1    g177(.A1(KEYINPUT70), .A2(KEYINPUT22), .ZN(new_n379));
  NAND2_X1  g178(.A1(G211gat), .A2(G218gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(KEYINPUT70), .A2(KEYINPUT22), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G211gat), .B(G218gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(G197gat), .B(G204gat), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n383), .B1(new_n382), .B2(new_n384), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(G226gat), .A2(G233gat), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT29), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n390), .B1(new_n254), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n389), .B1(new_n243), .B2(new_n253), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n388), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n254), .A2(new_n390), .ZN(new_n395));
  INV_X1    g194(.A(new_n388), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT29), .B1(new_n243), .B2(new_n253), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n395), .B(new_n396), .C1(new_n390), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  XOR2_X1   g198(.A(G8gat), .B(G36gat), .Z(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(KEYINPUT71), .ZN(new_n401));
  XNOR2_X1  g200(.A(G64gat), .B(G92gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n399), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n394), .A2(new_n403), .A3(new_n398), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(KEYINPUT30), .A3(new_n406), .ZN(new_n407));
  OR3_X1    g206(.A1(new_n399), .A2(KEYINPUT30), .A3(new_n404), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NOR3_X1   g208(.A1(new_n377), .A2(new_n378), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT37), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n411), .A3(new_n398), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n404), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n411), .B1(new_n394), .B2(new_n398), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT38), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT88), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT88), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n417), .B(KEYINPUT38), .C1(new_n413), .C2(new_n414), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT38), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n412), .A2(new_n419), .A3(new_n404), .ZN(new_n420));
  XOR2_X1   g219(.A(KEYINPUT66), .B(KEYINPUT28), .Z(new_n421));
  NAND3_X1  g220(.A1(new_n228), .A2(new_n230), .A3(new_n224), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n423), .A2(new_n207), .A3(new_n232), .ZN(new_n424));
  INV_X1    g223(.A(new_n242), .ZN(new_n425));
  OAI22_X1  g224(.A1(new_n424), .A2(new_n425), .B1(new_n212), .B2(new_n221), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n426), .B1(KEYINPUT25), .B2(new_n252), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n389), .B1(new_n427), .B2(KEYINPUT29), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n396), .B1(new_n428), .B2(new_n395), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n392), .A2(new_n388), .A3(new_n393), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT37), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT87), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n414), .A2(KEYINPUT87), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n420), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n416), .A2(new_n406), .A3(new_n418), .A4(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n304), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n374), .A2(KEYINPUT6), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n366), .A2(new_n368), .B1(new_n370), .B2(new_n372), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT6), .B1(new_n441), .B2(new_n304), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n376), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT86), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT86), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n442), .A2(new_n376), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n440), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n410), .B1(new_n437), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n396), .B1(new_n339), .B2(new_n391), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n345), .B1(new_n388), .B2(KEYINPUT29), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n348), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT83), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n451), .A2(new_n348), .A3(KEYINPUT83), .ZN(new_n455));
  INV_X1    g254(.A(G228gat), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n456), .A2(new_n276), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n450), .A2(new_n454), .A3(new_n455), .A4(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n457), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT80), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n386), .A2(new_n387), .A3(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n391), .B1(new_n385), .B2(KEYINPUT80), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n322), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n348), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT81), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n464), .B1(new_n449), .B2(new_n465), .ZN(new_n466));
  AOI211_X1 g265(.A(KEYINPUT81), .B(new_n396), .C1(new_n339), .C2(new_n391), .ZN(new_n467));
  OAI211_X1 g266(.A(KEYINPUT82), .B(new_n459), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT29), .B1(new_n344), .B2(new_n322), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT81), .B1(new_n470), .B2(new_n396), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n449), .A2(new_n465), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(new_n472), .A3(new_n464), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT82), .B1(new_n473), .B2(new_n459), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n458), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(G22gat), .ZN(new_n476));
  INV_X1    g275(.A(G22gat), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n477), .B(new_n458), .C1(new_n469), .C2(new_n474), .ZN(new_n478));
  XNOR2_X1  g277(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n479), .B(G50gat), .ZN(new_n480));
  XOR2_X1   g279(.A(G78gat), .B(G106gat), .Z(new_n481));
  XOR2_X1   g280(.A(new_n480), .B(new_n481), .Z(new_n482));
  NAND4_X1  g281(.A1(new_n476), .A2(KEYINPUT84), .A3(new_n478), .A4(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT84), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n478), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n486), .A2(new_n482), .B1(new_n476), .B2(new_n478), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n299), .B1(new_n448), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n442), .B1(new_n304), .B2(new_n441), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n490), .A2(new_n439), .B1(new_n408), .B2(new_n407), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n492), .B1(new_n484), .B2(new_n487), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n447), .A2(KEYINPUT35), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n291), .A2(new_n295), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n488), .A2(new_n494), .A3(new_n409), .A4(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n458), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n459), .B1(new_n466), .B2(new_n467), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT82), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n497), .B1(new_n500), .B2(new_n468), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT84), .B1(new_n501), .B2(new_n477), .ZN(new_n502));
  INV_X1    g301(.A(new_n482), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n500), .A2(new_n468), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n477), .B1(new_n504), .B2(new_n458), .ZN(new_n505));
  AOI211_X1 g304(.A(G22gat), .B(new_n497), .C1(new_n500), .C2(new_n468), .ZN(new_n506));
  OAI22_X1  g305(.A1(new_n502), .A2(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n507), .A2(new_n491), .A3(new_n483), .A4(new_n495), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT35), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n489), .A2(new_n493), .B1(new_n496), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G113gat), .B(G141gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(G197gat), .ZN(new_n512));
  XOR2_X1   g311(.A(KEYINPUT11), .B(G169gat), .Z(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  XOR2_X1   g313(.A(new_n514), .B(KEYINPUT12), .Z(new_n515));
  XNOR2_X1  g314(.A(G15gat), .B(G22gat), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT90), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(G1gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT16), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n516), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n516), .A2(new_n517), .A3(G1gat), .ZN(new_n522));
  INV_X1    g321(.A(G8gat), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n521), .A2(new_n522), .B1(KEYINPUT91), .B2(new_n523), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n523), .A2(KEYINPUT91), .ZN(new_n525));
  OR2_X1    g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n525), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G29gat), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n529), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(KEYINPUT14), .B(G29gat), .ZN(new_n531));
  INV_X1    g330(.A(G36gat), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(G43gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(G50gat), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT89), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT15), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G43gat), .B(G50gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT15), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n533), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n543), .B1(new_n538), .B2(new_n539), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n528), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n526), .A2(new_n545), .A3(new_n527), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(KEYINPUT92), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n550), .B(KEYINPUT13), .Z(new_n551));
  INV_X1    g350(.A(KEYINPUT92), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n528), .A2(new_n552), .A3(new_n546), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n549), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n545), .A2(KEYINPUT17), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n556), .B1(new_n541), .B2(new_n544), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n555), .A2(new_n557), .B1(new_n527), .B2(new_n526), .ZN(new_n558));
  INV_X1    g357(.A(new_n548), .ZN(new_n559));
  INV_X1    g358(.A(new_n550), .ZN(new_n560));
  NOR3_X1   g359(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n554), .B1(new_n561), .B2(KEYINPUT18), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(KEYINPUT18), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n515), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n561), .A2(KEYINPUT18), .ZN(new_n566));
  INV_X1    g365(.A(new_n515), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n566), .A2(new_n567), .A3(new_n563), .A4(new_n554), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n510), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G71gat), .B(G78gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT95), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT94), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(G57gat), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n575), .B(G64gat), .Z(new_n576));
  AOI21_X1  g375(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n577));
  OR3_X1    g376(.A1(new_n573), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(G57gat), .B(G64gat), .Z(new_n579));
  INV_X1    g378(.A(new_n577), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT93), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n579), .A2(new_n580), .B1(new_n572), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n582), .B1(new_n581), .B2(new_n572), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT21), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G231gat), .A2(G233gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(G127gat), .B(G155gat), .Z(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT96), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n588), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G183gat), .B(G211gat), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n528), .B1(new_n585), .B2(new_n584), .ZN(new_n596));
  XOR2_X1   g395(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n593), .A2(new_n598), .A3(new_n594), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT100), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT101), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT41), .ZN(new_n607));
  NAND2_X1  g406(.A1(G232gat), .A2(G233gat), .ZN(new_n608));
  OAI22_X1  g407(.A1(new_n605), .A2(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(KEYINPUT97), .B(G92gat), .Z(new_n610));
  INV_X1    g409(.A(G85gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(G99gat), .A2(G106gat), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n610), .A2(new_n611), .B1(KEYINPUT8), .B2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT98), .ZN(new_n614));
  XOR2_X1   g413(.A(G99gat), .B(G106gat), .Z(new_n615));
  NAND2_X1  g414(.A1(G85gat), .A2(G92gat), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n616), .A2(KEYINPUT7), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(KEYINPUT7), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n615), .A2(KEYINPUT99), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n615), .A2(KEYINPUT99), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n621), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n614), .A2(new_n623), .A3(new_n619), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n609), .B1(new_n625), .B2(new_n545), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n555), .A2(new_n557), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n627), .A2(new_n622), .A3(new_n624), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n605), .A2(new_n606), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n626), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G134gat), .B(G162gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n608), .A2(new_n607), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n632), .B(new_n633), .Z(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n629), .B1(new_n626), .B2(new_n628), .ZN(new_n636));
  OR3_X1    g435(.A1(new_n631), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n635), .B1(new_n631), .B2(new_n636), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n603), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G120gat), .B(G148gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(G176gat), .B(G204gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n642), .B(new_n643), .Z(new_n644));
  INV_X1    g443(.A(new_n584), .ZN(new_n645));
  INV_X1    g444(.A(new_n624), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n623), .B1(new_n614), .B2(new_n619), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n622), .A2(new_n584), .A3(new_n624), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n625), .A2(KEYINPUT10), .A3(new_n645), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(G230gat), .A2(G233gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n648), .A2(new_n649), .ZN(new_n656));
  INV_X1    g455(.A(new_n654), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n644), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n655), .A2(new_n658), .A3(new_n644), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n641), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n571), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n490), .A2(new_n439), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(new_n519), .ZN(G1324gat));
  INV_X1    g466(.A(new_n664), .ZN(new_n668));
  INV_X1    g467(.A(new_n409), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n520), .A2(new_n523), .ZN(new_n671));
  NOR2_X1   g470(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n523), .B1(new_n668), .B2(new_n669), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT42), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n676), .B1(KEYINPUT42), .B2(new_n674), .ZN(G1325gat));
  AOI21_X1  g476(.A(G15gat), .B1(new_n668), .B2(new_n495), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n299), .A2(G15gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT102), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n678), .B1(new_n668), .B2(new_n680), .ZN(G1326gat));
  NOR3_X1   g480(.A1(new_n510), .A2(new_n488), .A3(new_n570), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n663), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT43), .B(G22gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1327gat));
  INV_X1    g484(.A(new_n665), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n603), .A2(new_n640), .A3(new_n662), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n571), .A2(new_n529), .A3(new_n686), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT45), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n662), .B(KEYINPUT103), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n690), .A2(new_n569), .A3(new_n602), .ZN(new_n691));
  OAI21_X1  g490(.A(KEYINPUT44), .B1(new_n510), .B2(new_n640), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n507), .A2(new_n409), .A3(new_n483), .A4(new_n495), .ZN(new_n693));
  INV_X1    g492(.A(new_n494), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n509), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n495), .A2(KEYINPUT36), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n296), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n507), .A2(new_n483), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n356), .A2(new_n361), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT40), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n669), .A2(new_n376), .A3(new_n701), .A4(new_n363), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n442), .A2(new_n376), .A3(new_n445), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n445), .B1(new_n442), .B2(new_n376), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n439), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n702), .B1(new_n705), .B2(new_n436), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n493), .B(new_n697), .C1(new_n698), .C2(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n640), .B1(new_n695), .B2(new_n707), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n691), .B1(new_n692), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n686), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n689), .B1(new_n529), .B2(new_n713), .ZN(G1328gat));
  NAND2_X1  g513(.A1(new_n571), .A2(new_n687), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n715), .A2(G36gat), .A3(new_n409), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT46), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n711), .A2(new_n669), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n717), .B1(new_n532), .B2(new_n719), .ZN(G1329gat));
  NAND3_X1  g519(.A1(new_n711), .A2(G43gat), .A3(new_n299), .ZN(new_n721));
  INV_X1    g520(.A(new_n495), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n534), .B1(new_n715), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1330gat));
  INV_X1    g525(.A(new_n691), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n695), .A2(new_n707), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n728), .B1(new_n729), .B2(new_n639), .ZN(new_n730));
  INV_X1    g529(.A(new_n709), .ZN(new_n731));
  AOI211_X1 g530(.A(new_n640), .B(new_n731), .C1(new_n695), .C2(new_n707), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n698), .B(new_n727), .C1(new_n730), .C2(new_n732), .ZN(new_n733));
  NOR4_X1   g532(.A1(new_n603), .A2(G50gat), .A3(new_n640), .A4(new_n662), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n733), .A2(G50gat), .B1(new_n682), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT48), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT106), .A2(KEYINPUT48), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n735), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n738), .A2(new_n741), .ZN(G1331gat));
  NOR3_X1   g541(.A1(new_n641), .A2(new_n569), .A3(new_n690), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n729), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(new_n665), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g545(.A1(new_n744), .A2(new_n409), .ZN(new_n747));
  NOR2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  AND2_X1   g547(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(new_n747), .B2(new_n748), .ZN(G1333gat));
  OAI21_X1  g550(.A(G71gat), .B1(new_n744), .B2(new_n697), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n722), .A2(G71gat), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n744), .B2(new_n753), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n754), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g554(.A1(new_n744), .A2(new_n488), .ZN(new_n756));
  XNOR2_X1  g555(.A(KEYINPUT107), .B(G78gat), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1335gat));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n697), .B1(new_n706), .B2(new_n698), .ZN(new_n761));
  INV_X1    g560(.A(new_n493), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n693), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n764), .A2(new_n494), .B1(KEYINPUT35), .B2(new_n508), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n760), .B(new_n639), .C1(new_n763), .C2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n602), .A2(new_n570), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n760), .B1(new_n729), .B2(new_n639), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n759), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n767), .B1(new_n708), .B2(new_n760), .ZN(new_n772));
  OAI21_X1  g571(.A(KEYINPUT108), .B1(new_n510), .B2(new_n640), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n772), .A2(new_n773), .A3(KEYINPUT51), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n686), .A2(new_n662), .A3(new_n611), .ZN(new_n776));
  XOR2_X1   g575(.A(new_n776), .B(KEYINPUT109), .Z(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n662), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n767), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n692), .B2(new_n710), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(G85gat), .B1(new_n783), .B2(new_n665), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n778), .A2(new_n784), .ZN(G1336gat));
  OAI211_X1 g584(.A(new_n669), .B(new_n780), .C1(new_n730), .C2(new_n732), .ZN(new_n786));
  INV_X1    g585(.A(new_n610), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT110), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n690), .A2(G92gat), .A3(new_n409), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n793), .B1(new_n771), .B2(new_n774), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n610), .B1(new_n782), .B2(new_n669), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n790), .B(new_n791), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n769), .A2(new_n759), .A3(new_n770), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT51), .B1(new_n772), .B2(new_n773), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n792), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n799), .B(new_n788), .C1(new_n789), .C2(KEYINPUT52), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n796), .A2(new_n800), .ZN(G1337gat));
  NOR3_X1   g600(.A1(new_n779), .A2(new_n722), .A3(G99gat), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n775), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(G99gat), .B1(new_n783), .B2(new_n697), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(G1338gat));
  OR3_X1    g604(.A1(new_n690), .A2(G106gat), .A3(new_n488), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n771), .B2(new_n774), .ZN(new_n807));
  INV_X1    g606(.A(G106gat), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n808), .B1(new_n782), .B2(new_n698), .ZN(new_n809));
  OR3_X1    g608(.A1(new_n807), .A2(new_n809), .A3(KEYINPUT53), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT53), .B1(new_n807), .B2(new_n809), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(G1339gat));
  NAND3_X1  g611(.A1(new_n651), .A2(new_n652), .A3(new_n657), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n655), .A2(KEYINPUT54), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n657), .B1(new_n651), .B2(new_n652), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n644), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n814), .A2(KEYINPUT55), .A3(new_n817), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n820), .A2(new_n569), .A3(new_n661), .A4(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n558), .A2(new_n559), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(new_n550), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n551), .B1(new_n549), .B2(new_n553), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n514), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n662), .A2(new_n568), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n639), .B1(new_n822), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n820), .A2(new_n661), .A3(new_n821), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n637), .A2(new_n568), .A3(new_n638), .A4(new_n826), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n602), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n603), .A2(new_n570), .A3(new_n640), .A4(new_n779), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n698), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n665), .A2(new_n669), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n835), .A2(new_n495), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(G113gat), .B1(new_n838), .B2(new_n570), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n832), .A2(new_n833), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n686), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n693), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(new_n265), .A3(new_n569), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(KEYINPUT111), .ZN(G1340gat));
  AOI21_X1  g644(.A(G120gat), .B1(new_n842), .B2(new_n662), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n690), .A2(new_n263), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n837), .B2(new_n847), .ZN(G1341gat));
  NOR3_X1   g647(.A1(new_n841), .A2(new_n693), .A3(new_n602), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n849), .A2(KEYINPUT112), .ZN(new_n850));
  AOI21_X1  g649(.A(G127gat), .B1(new_n849), .B2(KEYINPUT112), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n602), .A2(new_n258), .ZN(new_n852));
  AOI22_X1  g651(.A1(new_n850), .A2(new_n851), .B1(new_n837), .B2(new_n852), .ZN(G1342gat));
  OAI21_X1  g652(.A(G134gat), .B1(new_n838), .B2(new_n640), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n842), .A2(new_n260), .A3(new_n639), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n855), .A2(KEYINPUT113), .A3(KEYINPUT56), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT113), .B1(new_n855), .B2(KEYINPUT56), .ZN(new_n857));
  OAI221_X1 g656(.A(new_n854), .B1(KEYINPUT56), .B2(new_n855), .C1(new_n856), .C2(new_n857), .ZN(G1343gat));
  NAND2_X1  g657(.A1(new_n840), .A2(new_n698), .ZN(new_n859));
  XOR2_X1   g658(.A(KEYINPUT114), .B(KEYINPUT57), .Z(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n488), .B1(new_n832), .B2(new_n833), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n697), .A2(new_n835), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n862), .A2(new_n569), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n324), .A2(new_n325), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n299), .A2(new_n488), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n871), .A2(KEYINPUT115), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n669), .B1(new_n871), .B2(KEYINPUT115), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n840), .A2(new_n872), .A3(new_n686), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n569), .A2(new_n316), .ZN(new_n875));
  XOR2_X1   g674(.A(new_n875), .B(KEYINPUT116), .Z(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n870), .A2(KEYINPUT118), .A3(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n880), .A2(new_n881), .A3(KEYINPUT58), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n878), .B1(new_n867), .B2(new_n869), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT117), .B1(new_n883), .B2(KEYINPUT118), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT58), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n885), .B1(new_n883), .B2(KEYINPUT117), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n882), .B1(new_n884), .B2(new_n886), .ZN(G1344gat));
  XOR2_X1   g686(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n888));
  NAND2_X1  g687(.A1(new_n866), .A2(new_n662), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n863), .A2(KEYINPUT57), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n863), .A2(new_n861), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n888), .B1(new_n893), .B2(new_n314), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n862), .A2(new_n662), .A3(new_n865), .A4(new_n866), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n314), .A2(KEYINPUT59), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n895), .A2(KEYINPUT119), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(KEYINPUT119), .B1(new_n895), .B2(new_n896), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n874), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n314), .A3(new_n662), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(G1345gat));
  NAND3_X1  g701(.A1(new_n862), .A2(new_n865), .A3(new_n866), .ZN(new_n903));
  OAI21_X1  g702(.A(G155gat), .B1(new_n903), .B2(new_n602), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n900), .A2(new_n306), .A3(new_n603), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n904), .A2(KEYINPUT121), .A3(new_n905), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1346gat));
  OAI21_X1  g709(.A(new_n307), .B1(new_n874), .B2(new_n640), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n639), .A2(G162gat), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n911), .B1(new_n903), .B2(new_n912), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT122), .ZN(G1347gat));
  NOR3_X1   g713(.A1(new_n722), .A2(new_n686), .A3(new_n409), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n834), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(G169gat), .B1(new_n916), .B2(new_n570), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n917), .A2(KEYINPUT124), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n917), .A2(KEYINPUT124), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n686), .B1(new_n832), .B2(new_n833), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n698), .A2(new_n409), .A3(new_n722), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(KEYINPUT123), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT123), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n569), .A2(new_n215), .ZN(new_n928));
  OAI22_X1  g727(.A1(new_n918), .A2(new_n919), .B1(new_n927), .B2(new_n928), .ZN(G1348gat));
  NOR3_X1   g728(.A1(new_n916), .A2(new_n216), .A3(new_n690), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n924), .A2(new_n662), .A3(new_n926), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(new_n216), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT125), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT125), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n931), .A2(new_n934), .A3(new_n216), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n930), .B1(new_n933), .B2(new_n935), .ZN(G1349gat));
  OAI21_X1  g735(.A(G183gat), .B1(new_n916), .B2(new_n602), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n603), .A2(new_n225), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n922), .B2(new_n938), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g739(.A(G190gat), .B1(new_n916), .B2(new_n640), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n941), .A2(KEYINPUT126), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(KEYINPUT126), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n942), .A2(KEYINPUT61), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n639), .A2(new_n224), .ZN(new_n945));
  OAI221_X1 g744(.A(new_n944), .B1(KEYINPUT61), .B2(new_n943), .C1(new_n927), .C2(new_n945), .ZN(G1351gat));
  INV_X1    g745(.A(G197gat), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n299), .A2(new_n686), .A3(new_n409), .ZN(new_n948));
  INV_X1    g747(.A(new_n892), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n569), .B(new_n948), .C1(new_n949), .C2(new_n890), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n947), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n952), .B1(new_n951), .B2(new_n950), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n299), .A2(new_n488), .A3(new_n409), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n920), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n569), .A2(new_n947), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(G1352gat));
  NOR3_X1   g756(.A1(new_n955), .A2(G204gat), .A3(new_n779), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n958), .B(KEYINPUT62), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n948), .B1(new_n949), .B2(new_n890), .ZN(new_n960));
  OAI21_X1  g759(.A(G204gat), .B1(new_n960), .B2(new_n690), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n961), .ZN(G1353gat));
  OR3_X1    g761(.A1(new_n955), .A2(G211gat), .A3(new_n602), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n603), .B(new_n948), .C1(new_n949), .C2(new_n890), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n964), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT63), .B1(new_n964), .B2(G211gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(G1354gat));
  OAI21_X1  g766(.A(G218gat), .B1(new_n960), .B2(new_n640), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n640), .A2(G218gat), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n968), .B1(new_n955), .B2(new_n969), .ZN(G1355gat));
endmodule


