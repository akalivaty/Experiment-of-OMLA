//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n569, new_n570, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197, new_n1198;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  AND3_X1   g037(.A1(new_n460), .A2(new_n462), .A3(KEYINPUT65), .ZN(new_n463));
  AOI21_X1  g038(.A(KEYINPUT65), .B1(new_n460), .B2(new_n462), .ZN(new_n464));
  OAI21_X1  g039(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n458), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n461), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n468), .A2(new_n460), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n470), .B1(new_n459), .B2(KEYINPUT3), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n469), .A2(G137), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G101), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n467), .A2(new_n474), .ZN(G160));
  AND2_X1   g050(.A1(new_n469), .A2(new_n471), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(new_n458), .B2(G112), .ZN(new_n480));
  OAI22_X1  g055(.A1(new_n477), .A2(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n476), .A2(new_n458), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n481), .B1(G136), .B2(new_n483), .ZN(G162));
  OAI211_X1 g059(.A(G138), .B(new_n458), .C1(new_n463), .C2(new_n464), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n471), .A2(new_n468), .A3(G126), .A4(new_n460), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(new_n459), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  AND2_X1   g066(.A1(KEYINPUT4), .A2(G138), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n471), .A2(new_n468), .A3(new_n460), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(G102), .A2(G2104), .ZN(new_n494));
  AOI21_X1  g069(.A(G2105), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n487), .A2(new_n491), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT67), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n495), .B1(new_n485), .B2(new_n486), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(KEYINPUT67), .A3(new_n491), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  OR2_X1    g078(.A1(KEYINPUT69), .A2(KEYINPUT6), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT69), .A2(KEYINPUT6), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n504), .A2(G651), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT68), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT68), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G651), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n508), .A2(new_n510), .A3(KEYINPUT6), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT5), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(KEYINPUT70), .A3(G543), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n506), .A2(new_n511), .A3(G543), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n508), .A2(new_n510), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n518), .A2(G62), .ZN(new_n526));
  NAND2_X1  g101(.A1(G75), .A2(G543), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n523), .A2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NAND2_X1  g105(.A1(new_n506), .A2(new_n511), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n515), .A2(new_n517), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G89), .ZN(new_n534));
  AND2_X1   g109(.A1(G63), .A2(G651), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n518), .A2(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT71), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n522), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n506), .A2(new_n511), .A3(KEYINPUT71), .A4(G543), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n542), .A2(G51), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n540), .A2(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  NAND2_X1  g121(.A1(new_n542), .A2(new_n543), .ZN(new_n547));
  INV_X1    g122(.A(G52), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(G77), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G64), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n532), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n533), .A2(G90), .B1(new_n553), .B2(new_n524), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n550), .A2(new_n554), .ZN(G301));
  INV_X1    g130(.A(G301), .ZN(G171));
  NAND3_X1  g131(.A1(new_n542), .A2(G43), .A3(new_n543), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n533), .A2(G81), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT72), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT72), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n557), .A2(new_n561), .A3(new_n558), .ZN(new_n562));
  NAND2_X1  g137(.A1(G68), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G56), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n532), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n560), .A2(new_n562), .B1(new_n524), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n532), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G651), .ZN(new_n575));
  INV_X1    g150(.A(G91), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n519), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(G53), .ZN(new_n578));
  OAI21_X1  g153(.A(KEYINPUT9), .B1(new_n522), .B2(new_n578), .ZN(new_n579));
  OR3_X1    g154(.A1(new_n522), .A2(KEYINPUT9), .A3(new_n578), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n577), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G299));
  NAND2_X1  g157(.A1(new_n533), .A2(G87), .ZN(new_n583));
  INV_X1    g158(.A(new_n522), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(G49), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n583), .A2(new_n585), .A3(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(new_n533), .A2(G86), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(G48), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n532), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(new_n524), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n588), .A2(new_n589), .A3(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT73), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n594), .B(new_n595), .ZN(G305));
  NAND2_X1  g171(.A1(new_n533), .A2(G85), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G47), .ZN(new_n599));
  OAI221_X1 g174(.A(new_n597), .B1(new_n525), .B2(new_n598), .C1(new_n547), .C2(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n518), .A2(G92), .A3(new_n511), .A4(new_n506), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n602), .B(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n542), .A2(G54), .A3(new_n543), .ZN(new_n605));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  XOR2_X1   g181(.A(KEYINPUT74), .B(G66), .Z(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n532), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G651), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n604), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n601), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n601), .B1(new_n611), .B2(G868), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G868), .B2(new_n581), .ZN(G297));
  OAI21_X1  g190(.A(new_n614), .B1(G868), .B2(new_n581), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n611), .B1(new_n617), .B2(G860), .ZN(G148));
  INV_X1    g193(.A(new_n566), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n610), .A2(G559), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT75), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n621), .B1(new_n623), .B2(G868), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g200(.A(new_n464), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n460), .A2(new_n462), .A3(KEYINPUT65), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n628), .A2(G2104), .A3(new_n458), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT76), .B(KEYINPUT12), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n629), .B(new_n630), .Z(new_n631));
  XOR2_X1   g206(.A(KEYINPUT77), .B(KEYINPUT13), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G2100), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT78), .Z(new_n635));
  INV_X1    g210(.A(G123), .ZN(new_n636));
  NOR2_X1   g211(.A1(G99), .A2(G2105), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(new_n458), .B2(G111), .ZN(new_n638));
  OAI22_X1  g213(.A1(new_n477), .A2(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n639), .B1(G135), .B2(new_n483), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2096), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n635), .B(new_n641), .C1(G2100), .C2(new_n633), .ZN(G156));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(KEYINPUT14), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n648), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2443), .B(G2446), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT79), .ZN(new_n657));
  OAI211_X1 g232(.A(new_n657), .B(G14), .C1(new_n655), .C2(new_n653), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G401));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT18), .Z(new_n665));
  INV_X1    g240(.A(new_n663), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n662), .B1(new_n666), .B2(new_n660), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n667), .A2(KEYINPUT80), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(KEYINPUT80), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n660), .B(KEYINPUT17), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n668), .B(new_n669), .C1(new_n666), .C2(new_n670), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(new_n662), .A3(new_n666), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n665), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(G2096), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G2100), .ZN(G227));
  XOR2_X1   g250(.A(G1971), .B(G1976), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT81), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1956), .B(G2474), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1961), .B(G1966), .ZN(new_n680));
  NOR3_X1   g255(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT20), .Z(new_n682));
  AND2_X1   g257(.A1(new_n679), .A2(new_n680), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(new_n680), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n683), .B1(new_n678), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n678), .A2(KEYINPUT82), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n682), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT83), .B(G1981), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n688), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G229));
  XNOR2_X1  g271(.A(KEYINPUT93), .B(KEYINPUT25), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  AOI22_X1  g274(.A1(new_n628), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n700), .A2(new_n458), .ZN(new_n701));
  AOI211_X1 g276(.A(new_n699), .B(new_n701), .C1(G139), .C2(new_n483), .ZN(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(new_n703), .B2(G33), .ZN(new_n705));
  INV_X1    g280(.A(G2072), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT94), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G5), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G171), .B2(new_n709), .ZN(new_n711));
  INV_X1    g286(.A(G1961), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n703), .A2(G32), .ZN(new_n714));
  NAND3_X1  g289(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT95), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT26), .ZN(new_n717));
  INV_X1    g292(.A(G129), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n717), .B1(new_n718), .B2(new_n477), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n476), .A2(G141), .ZN(new_n720));
  NAND2_X1  g295(.A1(G105), .A2(G2104), .ZN(new_n721));
  AOI21_X1  g296(.A(G2105), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n714), .B1(new_n723), .B2(new_n703), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT96), .Z(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT27), .B(G1996), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n703), .A2(G26), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT28), .ZN(new_n730));
  OR2_X1    g305(.A1(G104), .A2(G2105), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n731), .B(G2104), .C1(G116), .C2(new_n458), .ZN(new_n732));
  INV_X1    g307(.A(G140), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n482), .B2(new_n733), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n476), .A2(G2105), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT92), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n735), .A2(new_n736), .A3(G128), .ZN(new_n737));
  INV_X1    g312(.A(G128), .ZN(new_n738));
  OAI21_X1  g313(.A(KEYINPUT92), .B1(new_n477), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n734), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n730), .B1(new_n740), .B2(new_n703), .ZN(new_n741));
  INV_X1    g316(.A(G2067), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n708), .A2(new_n713), .A3(new_n728), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n640), .A2(G29), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT31), .B(G11), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT98), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT30), .ZN(new_n748));
  AOI21_X1  g323(.A(G29), .B1(new_n748), .B2(G28), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n748), .B2(G28), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n745), .A2(new_n747), .A3(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT24), .ZN(new_n752));
  INV_X1    g327(.A(G34), .ZN(new_n753));
  AOI21_X1  g328(.A(G29), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n752), .B2(new_n753), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G160), .B2(new_n703), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n751), .B1(G2084), .B2(new_n756), .ZN(new_n757));
  OAI221_X1 g332(.A(new_n757), .B1(G2084), .B2(new_n756), .C1(new_n705), .C2(new_n706), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n709), .A2(G21), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G168), .B2(new_n709), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1966), .ZN(new_n761));
  NOR3_X1   g336(.A1(new_n744), .A2(new_n758), .A3(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n725), .A2(new_n727), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT97), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n703), .A2(G27), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G164), .B2(new_n703), .ZN(new_n766));
  INV_X1    g341(.A(G2078), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n566), .A2(new_n709), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n709), .B2(G19), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n764), .B(new_n768), .C1(G1341), .C2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n709), .A2(G4), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n611), .B2(new_n709), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT91), .ZN(new_n776));
  INV_X1    g351(.A(G1348), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n703), .A2(G35), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G162), .B2(new_n703), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT29), .Z(new_n781));
  INV_X1    g356(.A(G2090), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n709), .A2(G20), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT23), .Z(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G299), .B2(G16), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G1956), .ZN(new_n787));
  INV_X1    g362(.A(new_n781), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(G2090), .ZN(new_n789));
  AOI211_X1 g364(.A(new_n783), .B(new_n789), .C1(G1341), .C2(new_n771), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n762), .A2(new_n773), .A3(new_n778), .A4(new_n790), .ZN(new_n791));
  MUX2_X1   g366(.A(G6), .B(G305), .S(G16), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT87), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT32), .B(G1981), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(KEYINPUT88), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(KEYINPUT88), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n709), .A2(G22), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G166), .B2(new_n709), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT90), .ZN(new_n800));
  INV_X1    g375(.A(G1971), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  MUX2_X1   g377(.A(G23), .B(G288), .S(G16), .Z(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT33), .B(G1976), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT89), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n803), .B(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n796), .A2(new_n797), .A3(new_n807), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT86), .B(KEYINPUT34), .Z(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n796), .A2(new_n797), .A3(new_n809), .A4(new_n807), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n703), .A2(G25), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(KEYINPUT84), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(KEYINPUT84), .ZN(new_n815));
  INV_X1    g390(.A(G119), .ZN(new_n816));
  NOR2_X1   g391(.A1(G95), .A2(G2105), .ZN(new_n817));
  OAI21_X1  g392(.A(G2104), .B1(new_n458), .B2(G107), .ZN(new_n818));
  OAI22_X1  g393(.A1(new_n477), .A2(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(G131), .B2(new_n483), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT85), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n814), .B(new_n815), .C1(new_n821), .C2(new_n703), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT35), .B(G1991), .Z(new_n824));
  OR2_X1    g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n709), .A2(G24), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(G290), .B2(G16), .ZN(new_n828));
  INV_X1    g403(.A(G1986), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n825), .A2(new_n826), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n811), .A2(new_n812), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(KEYINPUT36), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n832), .B1(new_n808), .B2(new_n810), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT36), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n836), .A2(new_n837), .A3(new_n812), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n791), .B1(new_n835), .B2(new_n838), .ZN(G311));
  INV_X1    g414(.A(new_n791), .ZN(new_n840));
  INV_X1    g415(.A(new_n838), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n837), .B1(new_n836), .B2(new_n812), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(G150));
  NAND2_X1  g418(.A1(G80), .A2(G543), .ZN(new_n844));
  INV_X1    g419(.A(G67), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n844), .B1(new_n532), .B2(new_n845), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n533), .A2(G93), .B1(new_n846), .B2(new_n524), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n542), .A2(G55), .A3(new_n543), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(KEYINPUT100), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT100), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n847), .A2(new_n851), .A3(new_n848), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n566), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n565), .A2(new_n524), .ZN(new_n854));
  INV_X1    g429(.A(new_n562), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n561), .B1(new_n557), .B2(new_n558), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n852), .B(new_n854), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n850), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n853), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n611), .A2(G559), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n862), .B(new_n863), .Z(new_n864));
  AND2_X1   g439(.A1(new_n864), .A2(KEYINPUT39), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n864), .A2(KEYINPUT39), .ZN(new_n866));
  NOR3_X1   g441(.A1(new_n865), .A2(new_n866), .A3(G860), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n849), .A2(G860), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT101), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(KEYINPUT37), .Z(new_n870));
  OR2_X1    g445(.A1(new_n867), .A2(new_n870), .ZN(G145));
  XNOR2_X1  g446(.A(new_n740), .B(new_n497), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n702), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n631), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n476), .A2(G142), .A3(new_n458), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT102), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n735), .A2(G130), .ZN(new_n877));
  NOR2_X1   g452(.A1(G106), .A2(G2105), .ZN(new_n878));
  OAI21_X1  g453(.A(G2104), .B1(new_n458), .B2(G118), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n876), .B(new_n877), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n820), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n723), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n874), .B(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n640), .B(G160), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n884), .B(G162), .Z(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(G37), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  NOR3_X1   g462(.A1(new_n883), .A2(KEYINPUT103), .A3(new_n886), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n889));
  INV_X1    g464(.A(new_n882), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n874), .B(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n889), .B1(new_n891), .B2(new_n885), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n887), .B1(new_n888), .B2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g469(.A(new_n623), .B(new_n860), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n610), .A2(new_n581), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n610), .A2(new_n581), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n895), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n610), .A2(new_n902), .A3(new_n581), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n902), .B1(new_n610), .B2(new_n581), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n903), .A2(new_n904), .A3(new_n896), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT105), .B1(new_n905), .B2(KEYINPUT41), .ZN(new_n906));
  INV_X1    g481(.A(new_n904), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n610), .A2(new_n581), .A3(new_n902), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(new_n897), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT105), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n896), .A2(new_n911), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n898), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n906), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n895), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n901), .A2(new_n916), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n917), .A2(KEYINPUT42), .ZN(new_n918));
  XNOR2_X1  g493(.A(G290), .B(G288), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT106), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n919), .B(KEYINPUT106), .ZN(new_n921));
  XNOR2_X1  g496(.A(G305), .B(G303), .ZN(new_n922));
  MUX2_X1   g497(.A(new_n920), .B(new_n921), .S(new_n922), .Z(new_n923));
  NAND2_X1  g498(.A1(new_n917), .A2(KEYINPUT42), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n918), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n923), .B1(new_n918), .B2(new_n924), .ZN(new_n926));
  OAI21_X1  g501(.A(G868), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n849), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n927), .B1(G868), .B2(new_n928), .ZN(G295));
  OAI21_X1  g504(.A(new_n927), .B1(G868), .B2(new_n928), .ZN(G331));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n554), .A2(KEYINPUT107), .A3(new_n550), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n933));
  INV_X1    g508(.A(new_n554), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n933), .B1(new_n934), .B2(new_n549), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n932), .A2(G168), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(G301), .A2(G286), .A3(new_n933), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n860), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n853), .A2(new_n859), .A3(new_n937), .A4(new_n936), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n915), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n939), .A2(KEYINPUT108), .A3(new_n940), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n860), .A2(new_n944), .A3(new_n938), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n900), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n942), .B1(new_n946), .B2(KEYINPUT109), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n948));
  AOI211_X1 g523(.A(new_n948), .B(new_n900), .C1(new_n943), .C2(new_n945), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT110), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n943), .A2(new_n945), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n899), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n948), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT110), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n946), .A2(KEYINPUT109), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n953), .A2(new_n954), .A3(new_n955), .A4(new_n942), .ZN(new_n956));
  INV_X1    g531(.A(new_n923), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n950), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n947), .A2(new_n949), .ZN(new_n959));
  AOI21_X1  g534(.A(G37), .B1(new_n959), .B2(new_n923), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n931), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n947), .A2(new_n957), .A3(new_n949), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n903), .A2(new_n904), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n963), .A2(new_n913), .B1(new_n899), .B2(new_n911), .ZN(new_n964));
  OAI22_X1  g539(.A1(new_n951), .A2(new_n964), .B1(new_n900), .B2(new_n941), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n965), .A2(new_n957), .ZN(new_n966));
  NOR4_X1   g541(.A1(new_n962), .A2(new_n966), .A3(KEYINPUT43), .A4(G37), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n961), .A2(KEYINPUT44), .A3(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n958), .A2(new_n960), .A3(new_n931), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OR2_X1    g546(.A1(new_n962), .A2(G37), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT43), .B1(new_n972), .B2(new_n966), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n958), .A2(new_n960), .A3(KEYINPUT111), .A4(new_n931), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n971), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n968), .B1(new_n975), .B2(KEYINPUT44), .ZN(G397));
  AOI21_X1  g551(.A(G1384), .B1(new_n500), .B2(new_n491), .ZN(new_n977));
  INV_X1    g552(.A(G40), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n467), .A2(new_n474), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n980), .A2(G8), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n594), .B(KEYINPUT49), .ZN(new_n982));
  INV_X1    g557(.A(G1981), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT117), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n983), .B1(new_n593), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n982), .B(new_n985), .ZN(new_n986));
  AOI211_X1 g561(.A(G1976), .B(G288), .C1(new_n986), .C2(new_n981), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n594), .A2(G1981), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n981), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(G303), .A2(G8), .ZN(new_n990));
  XOR2_X1   g565(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n991));
  NOR2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n992), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n996));
  AOI21_X1  g571(.A(G1384), .B1(new_n499), .B2(new_n501), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n996), .B1(new_n997), .B2(KEYINPUT45), .ZN(new_n998));
  INV_X1    g573(.A(G1384), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n500), .A2(KEYINPUT67), .A3(new_n491), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT67), .B1(new_n500), .B2(new_n491), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n999), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(KEYINPUT113), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n497), .A2(new_n999), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n979), .B1(new_n1005), .B2(new_n1003), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n998), .A2(new_n1004), .A3(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1008), .A2(KEYINPUT114), .A3(new_n801), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n979), .B1(new_n1005), .B2(KEYINPUT50), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1010), .B1(new_n1002), .B2(KEYINPUT50), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n782), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT114), .B1(new_n1008), .B2(new_n801), .ZN(new_n1014));
  OAI211_X1 g589(.A(G8), .B(new_n995), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n986), .A2(new_n981), .ZN(new_n1016));
  INV_X1    g591(.A(G1976), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n980), .B(G8), .C1(new_n1017), .C2(G288), .ZN(new_n1018));
  NAND2_X1  g593(.A1(KEYINPUT116), .A2(KEYINPUT52), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n1022));
  NAND3_X1  g597(.A1(G288), .A2(new_n1022), .A3(new_n1017), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1016), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n989), .B1(new_n1015), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT63), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT45), .B1(new_n502), .B2(new_n999), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1006), .B1(new_n1028), .B2(KEYINPUT113), .ZN(new_n1029));
  AOI21_X1  g604(.A(G1971), .B1(new_n1029), .B2(new_n998), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT50), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1032), .B1(new_n497), .B2(new_n999), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n472), .A2(new_n473), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n458), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n465), .A2(new_n466), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1035), .B(G40), .C1(new_n1036), .C2(new_n458), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1031), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1032), .B(new_n999), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1039));
  OAI211_X1 g614(.A(KEYINPUT118), .B(new_n979), .C1(new_n977), .C2(new_n1032), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(G2090), .ZN(new_n1042));
  OAI21_X1  g617(.A(G8), .B1(new_n1030), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1025), .B1(new_n1043), .B2(new_n994), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n1015), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1037), .B1(new_n977), .B2(new_n1032), .ZN(new_n1046));
  INV_X1    g621(.A(G2084), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1046), .B(new_n1047), .C1(new_n997), .C2(new_n1032), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n979), .B1(new_n977), .B2(KEYINPUT45), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1049), .B1(new_n997), .B2(KEYINPUT45), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1048), .B1(new_n1050), .B2(G1966), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1051), .A2(G8), .A3(G168), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1027), .B1(new_n1045), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(G8), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n994), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1025), .A2(new_n1027), .A3(new_n1052), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1055), .A2(new_n1015), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1026), .B1(new_n1053), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1046), .B1(new_n997), .B2(new_n1032), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n777), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT119), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n977), .A2(new_n979), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1061), .B1(new_n977), .B2(new_n979), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n742), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n610), .A2(KEYINPUT60), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1060), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1002), .A2(KEYINPUT50), .ZN(new_n1069));
  AOI21_X1  g644(.A(G1348), .B1(new_n1069), .B2(new_n1046), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1064), .ZN(new_n1071));
  AOI21_X1  g646(.A(G2067), .B1(new_n1071), .B2(new_n1062), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n611), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1060), .A2(new_n610), .A3(new_n1065), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1068), .B1(new_n1075), .B2(KEYINPUT60), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT56), .B(G2072), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n998), .A2(new_n1004), .A3(new_n1007), .A4(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n581), .B(KEYINPUT57), .ZN(new_n1079));
  INV_X1    g654(.A(G1956), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1041), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1078), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT61), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1078), .A2(new_n1081), .A3(KEYINPUT61), .A4(new_n1079), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G1996), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n998), .A2(new_n1004), .A3(new_n1087), .A4(new_n1007), .ZN(new_n1088));
  XOR2_X1   g663(.A(KEYINPUT58), .B(G1341), .Z(new_n1089));
  NAND3_X1  g664(.A1(new_n1071), .A2(new_n1062), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1091), .A2(KEYINPUT59), .A3(new_n566), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n566), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1076), .A2(new_n1086), .A3(new_n1092), .A4(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1079), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1073), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1097), .B1(new_n1098), .B2(new_n1082), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g675(.A(G301), .B(KEYINPUT54), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n1011), .B2(G1961), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1059), .A2(KEYINPUT122), .A3(new_n712), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1037), .B1(new_n1005), .B2(new_n1003), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1105), .B(KEYINPUT123), .ZN(new_n1106));
  NOR2_X1   g681(.A1(KEYINPUT124), .A2(G2078), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT124), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT53), .B1(new_n1108), .B2(new_n767), .ZN(new_n1109));
  AOI211_X1 g684(.A(new_n1107), .B(new_n1109), .C1(new_n977), .C2(KEYINPUT45), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1103), .A2(new_n1104), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(new_n1008), .B2(G2078), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1101), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1112), .A2(G2078), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1050), .A2(new_n1115), .B1(new_n1059), .B2(new_n712), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1113), .A2(new_n1116), .A3(new_n1101), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1048), .B(G168), .C1(new_n1050), .C2(G1966), .ZN(new_n1120));
  OAI211_X1 g695(.A(KEYINPUT45), .B(new_n999), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n1105), .ZN(new_n1122));
  INV_X1    g697(.A(G1966), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(G168), .B1(new_n1124), .B2(new_n1048), .ZN(new_n1125));
  NOR2_X1   g700(.A1(KEYINPUT120), .A2(KEYINPUT51), .ZN(new_n1126));
  OAI211_X1 g701(.A(G8), .B(new_n1120), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1120), .A2(G8), .ZN(new_n1128));
  XOR2_X1   g703(.A(KEYINPUT120), .B(KEYINPUT51), .Z(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1127), .A2(KEYINPUT121), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT121), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT62), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(G301), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1100), .A2(new_n1119), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1126), .B1(new_n1051), .B2(G286), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1137), .A2(new_n1128), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1129), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1139), .B1(new_n1120), .B2(G8), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1136), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1127), .A2(new_n1130), .A3(KEYINPUT121), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1134), .A2(KEYINPUT62), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT125), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1044), .A2(new_n1015), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1145), .B1(new_n1044), .B2(new_n1015), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1144), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1058), .B1(new_n1135), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1005), .A2(new_n1003), .A3(new_n979), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT112), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n740), .B(G2067), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n723), .B(G1996), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n820), .B(new_n824), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1152), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(G290), .A2(G1986), .ZN(new_n1158));
  AND2_X1   g733(.A1(G290), .A2(G1986), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1152), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1150), .A2(new_n1162), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1152), .A2(new_n1087), .ZN(new_n1164));
  OR2_X1    g739(.A1(new_n1164), .A2(KEYINPUT46), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1152), .A2(KEYINPUT46), .A3(new_n1087), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1153), .A2(new_n723), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(new_n1152), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1165), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1169), .B(KEYINPUT47), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n821), .A2(new_n824), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1171), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n740), .A2(new_n742), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1152), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  XOR2_X1   g749(.A(new_n1174), .B(KEYINPUT126), .Z(new_n1175));
  AND2_X1   g750(.A1(new_n1152), .A2(new_n1158), .ZN(new_n1176));
  OR2_X1    g751(.A1(new_n1176), .A2(KEYINPUT48), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(KEYINPUT48), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1177), .A2(new_n1157), .A3(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1170), .A2(new_n1175), .A3(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1163), .A2(KEYINPUT127), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT127), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1045), .A2(KEYINPUT125), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1184), .A2(new_n1146), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1134), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1186), .B1(new_n1187), .B2(KEYINPUT62), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1118), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1189));
  OAI211_X1 g764(.A(new_n1185), .B(new_n1144), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1161), .B1(new_n1190), .B2(new_n1058), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1183), .B1(new_n1191), .B2(new_n1180), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1182), .A2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g768(.A(G319), .ZN(new_n1195));
  NOR4_X1   g769(.A1(G229), .A2(G401), .A3(new_n1195), .A4(G227), .ZN(new_n1196));
  NAND2_X1  g770(.A1(new_n893), .A2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g771(.A1(new_n961), .A2(new_n967), .ZN(new_n1198));
  NOR2_X1   g772(.A1(new_n1197), .A2(new_n1198), .ZN(G308));
  OR2_X1    g773(.A1(new_n1197), .A2(new_n1198), .ZN(G225));
endmodule


