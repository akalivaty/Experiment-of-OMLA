//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1273, new_n1274, new_n1275, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n209));
  INV_X1    g0009(.A(G50), .ZN(new_n210));
  INV_X1    g0010(.A(G226), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n208), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n208), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XOR2_X1   g0021(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n222));
  XNOR2_X1  g0022(.A(new_n221), .B(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n225), .A2(new_n206), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT65), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(G58), .A2(G68), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  AND4_X1   g0033(.A1(new_n219), .A2(new_n223), .A3(new_n224), .A4(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT66), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(G97), .B(G107), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NAND3_X1  g0050(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G50), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n225), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n254), .B1(new_n205), .B2(G20), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n252), .B1(new_n255), .B2(G50), .ZN(new_n256));
  INV_X1    g0056(.A(G150), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  OAI22_X1  g0059(.A1(new_n257), .A2(new_n259), .B1(new_n201), .B2(new_n206), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n206), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT67), .ZN(new_n262));
  XNOR2_X1  g0062(.A(new_n261), .B(new_n262), .ZN(new_n263));
  XOR2_X1   g0063(.A(KEYINPUT8), .B(G58), .Z(new_n264));
  AOI21_X1  g0064(.A(new_n260), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n254), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n256), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT9), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g0069(.A(KEYINPUT9), .B(new_n256), .C1(new_n265), .C2(new_n266), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT68), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT10), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n269), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n271), .A2(KEYINPUT10), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G41), .ZN(new_n277));
  INV_X1    g0077(.A(G45), .ZN(new_n278));
  AOI21_X1  g0078(.A(G1), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G274), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(G1), .A3(G13), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n280), .B1(new_n284), .B2(new_n211), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT3), .B(G33), .ZN(new_n286));
  INV_X1    g0086(.A(G1698), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(G222), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(G1698), .ZN(new_n289));
  INV_X1    g0089(.A(G223), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n288), .B1(new_n202), .B2(new_n286), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n285), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G200), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(G190), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n274), .A2(new_n276), .A3(new_n295), .A4(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n296), .B1(new_n294), .B2(new_n293), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n275), .B1(new_n298), .B2(new_n273), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n293), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n267), .B1(new_n293), .B2(G169), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AND3_X1   g0103(.A1(new_n297), .A2(new_n299), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT14), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT70), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT13), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n286), .A2(G232), .A3(G1698), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n286), .A2(G226), .A3(new_n287), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G97), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n292), .ZN(new_n312));
  INV_X1    g0112(.A(G238), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n280), .B1(new_n284), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n307), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  AOI211_X1 g0116(.A(KEYINPUT13), .B(new_n314), .C1(new_n311), .C2(new_n292), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G169), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n306), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n305), .A2(KEYINPUT70), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(new_n318), .B2(G179), .ZN(new_n322));
  INV_X1    g0122(.A(new_n306), .ZN(new_n323));
  OAI211_X1 g0123(.A(G169), .B(new_n323), .C1(new_n316), .C2(new_n317), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n320), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n261), .B(KEYINPUT67), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(new_n202), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n259), .A2(new_n210), .B1(new_n206), .B2(G68), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n254), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT11), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI211_X1 g0131(.A(KEYINPUT11), .B(new_n254), .C1(new_n327), .C2(new_n328), .ZN(new_n332));
  OR3_X1    g0132(.A1(new_n251), .A2(KEYINPUT12), .A3(G68), .ZN(new_n333));
  OAI21_X1  g0133(.A(KEYINPUT12), .B1(new_n251), .B2(G68), .ZN(new_n334));
  AOI22_X1  g0134(.A1(G68), .A2(new_n255), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n331), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT69), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n331), .A2(KEYINPUT69), .A3(new_n332), .A4(new_n335), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n325), .A2(new_n340), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n338), .A2(new_n339), .B1(G190), .B2(new_n318), .ZN(new_n342));
  OAI21_X1  g0142(.A(G200), .B1(new_n316), .B2(new_n317), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n264), .A2(new_n258), .B1(G20), .B2(G77), .ZN(new_n345));
  XNOR2_X1  g0145(.A(KEYINPUT15), .B(G87), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n345), .B1(new_n261), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n254), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n255), .A2(G77), .ZN(new_n349));
  INV_X1    g0149(.A(new_n251), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n202), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n348), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G244), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n280), .B1(new_n284), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n286), .A2(G232), .A3(new_n287), .ZN(new_n355));
  INV_X1    g0155(.A(G107), .ZN(new_n356));
  OAI221_X1 g0156(.A(new_n355), .B1(new_n356), .B2(new_n286), .C1(new_n289), .C2(new_n313), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n354), .B1(new_n357), .B2(new_n292), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n352), .B1(G169), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n300), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n357), .A2(new_n292), .ZN(new_n363));
  INV_X1    g0163(.A(new_n354), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(G200), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n352), .B1(G190), .B2(new_n358), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n362), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n304), .A2(new_n341), .A3(new_n344), .A4(new_n368), .ZN(new_n369));
  AND2_X1   g0169(.A1(G58), .A2(G68), .ZN(new_n370));
  OAI21_X1  g0170(.A(G20), .B1(new_n370), .B2(new_n229), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT71), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n258), .A2(G159), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n372), .B1(new_n371), .B2(new_n373), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  NOR3_X1   g0177(.A1(new_n286), .A2(new_n377), .A3(G20), .ZN(new_n378));
  INV_X1    g0178(.A(G33), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT3), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT3), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(G33), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT7), .B1(new_n383), .B2(new_n206), .ZN(new_n384));
  OAI21_X1  g0184(.A(G68), .B1(new_n378), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n376), .A2(new_n385), .A3(KEYINPUT16), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  INV_X1    g0187(.A(G68), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n377), .B1(new_n286), .B2(G20), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n383), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n371), .A2(new_n373), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n387), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n386), .A2(new_n393), .A3(new_n254), .ZN(new_n394));
  INV_X1    g0194(.A(new_n264), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n251), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n255), .B2(new_n395), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n380), .A2(new_n382), .A3(G226), .A4(G1698), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n380), .A2(new_n382), .A3(G223), .A4(new_n287), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n399), .B(new_n400), .C1(new_n379), .C2(new_n212), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n292), .ZN(new_n402));
  INV_X1    g0202(.A(new_n280), .ZN(new_n403));
  INV_X1    g0203(.A(new_n284), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n403), .B1(new_n404), .B2(G232), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(G169), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n300), .B2(new_n406), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n398), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT18), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n409), .B(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n402), .A2(new_n405), .A3(G190), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n406), .A2(G200), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n394), .A2(new_n412), .A3(new_n397), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT17), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n413), .A2(new_n412), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT17), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n416), .A2(new_n394), .A3(new_n417), .A4(new_n397), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n415), .A2(new_n418), .A3(KEYINPUT72), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT72), .B1(new_n415), .B2(new_n418), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n411), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OR3_X1    g0221(.A1(new_n369), .A2(new_n421), .A3(KEYINPUT73), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT73), .B1(new_n369), .B2(new_n421), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n205), .A2(G45), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT5), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n425), .B1(new_n426), .B2(G41), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(KEYINPUT76), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT76), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT5), .ZN(new_n430));
  AOI21_X1  g0230(.A(G41), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT77), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n427), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  XNOR2_X1  g0233(.A(KEYINPUT76), .B(KEYINPUT5), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n434), .A2(KEYINPUT77), .A3(G41), .ZN(new_n435));
  OAI211_X1 g0235(.A(G264), .B(new_n282), .C1(new_n433), .C2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n286), .A2(G250), .A3(new_n287), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n286), .A2(G257), .A3(G1698), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G33), .A2(G294), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n292), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(KEYINPUT77), .B1(new_n434), .B2(G41), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n429), .A2(KEYINPUT5), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n426), .A2(KEYINPUT76), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n432), .B(new_n277), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n443), .A2(G274), .A3(new_n446), .A4(new_n427), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT78), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n278), .A2(G1), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(KEYINPUT5), .B2(new_n277), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n277), .B1(new_n444), .B2(new_n445), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n451), .B1(new_n452), .B2(KEYINPUT77), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n453), .A2(KEYINPUT78), .A3(G274), .A4(new_n446), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n442), .A2(G190), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT74), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(new_n379), .B2(G1), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n205), .A2(KEYINPUT74), .A3(G33), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(new_n251), .A3(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(new_n254), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT25), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n462), .B1(new_n251), .B2(G107), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n350), .A2(KEYINPUT25), .A3(new_n356), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n461), .A2(G107), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n380), .A2(new_n382), .A3(new_n206), .A4(G87), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT22), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT22), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n286), .A2(new_n469), .A3(new_n206), .A4(G87), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT23), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(new_n206), .B2(G107), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n356), .A2(KEYINPUT23), .A3(G20), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(G116), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n379), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n206), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n471), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT24), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n266), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n479), .B1(new_n468), .B2(new_n470), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT24), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n466), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n436), .A2(new_n441), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n487), .B1(new_n449), .B2(new_n454), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n456), .B(new_n486), .C1(new_n488), .C2(new_n294), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n449), .A2(new_n454), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G283), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n380), .A2(new_n382), .A3(G250), .A4(G1698), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n380), .A2(new_n382), .A3(G244), .A4(new_n287), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT75), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n491), .B(new_n492), .C1(new_n493), .C2(new_n495), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n493), .A2(new_n495), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n292), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g0298(.A(G257), .B(new_n282), .C1(new_n433), .C2(new_n435), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n319), .B1(new_n490), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n461), .A2(G97), .ZN(new_n502));
  INV_X1    g0302(.A(G97), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n350), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(G107), .B1(new_n378), .B2(new_n384), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n356), .A2(KEYINPUT6), .A3(G97), .ZN(new_n507));
  INV_X1    g0307(.A(new_n248), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G20), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n258), .A2(G77), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n506), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n505), .B1(new_n512), .B2(new_n254), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n455), .A2(new_n300), .A3(new_n498), .A4(new_n499), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n501), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(G200), .B1(new_n490), .B2(new_n500), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n455), .A2(G190), .A3(new_n498), .A4(new_n499), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(new_n513), .A3(new_n518), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n489), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n319), .B1(new_n490), .B2(new_n487), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n254), .B1(new_n484), .B2(KEYINPUT24), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n471), .A2(KEYINPUT24), .A3(new_n480), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n465), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n442), .A2(new_n300), .A3(new_n455), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n521), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n491), .B(new_n206), .C1(G33), .C2(new_n503), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n476), .A2(G20), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n527), .A2(new_n254), .A3(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT20), .ZN(new_n530));
  XNOR2_X1  g0330(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n251), .A2(G116), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n461), .B2(G116), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n319), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n286), .A2(G257), .A3(new_n287), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n383), .A2(G303), .ZN(new_n536));
  INV_X1    g0336(.A(G264), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n535), .B(new_n536), .C1(new_n289), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n292), .ZN(new_n539));
  OAI211_X1 g0339(.A(G270), .B(new_n282), .C1(new_n433), .C2(new_n435), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n534), .B1(new_n490), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(KEYINPUT79), .A2(KEYINPUT21), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n539), .A2(new_n540), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n531), .A2(new_n533), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n545), .A2(G179), .A3(new_n455), .A4(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n543), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n548), .B(new_n534), .C1(new_n490), .C2(new_n541), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n526), .A2(new_n544), .A3(new_n547), .A4(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n380), .A2(new_n382), .A3(G238), .A4(new_n287), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n380), .A2(new_n382), .A3(G244), .A4(G1698), .ZN(new_n553));
  INV_X1    g0353(.A(new_n477), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n292), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n450), .A2(G274), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n425), .A2(G250), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n557), .B1(new_n292), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n319), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n346), .A2(new_n350), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT19), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n206), .B1(new_n310), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n212), .A2(new_n503), .A3(new_n356), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n380), .A2(new_n382), .A3(new_n206), .A4(G68), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n565), .B1(new_n261), .B2(new_n503), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n564), .B1(new_n571), .B2(new_n254), .ZN(new_n572));
  INV_X1    g0372(.A(new_n461), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n572), .B1(new_n346), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n559), .B1(new_n555), .B2(new_n292), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n300), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n562), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(G190), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n461), .A2(G87), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n572), .B(new_n580), .C1(new_n575), .C2(new_n294), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n577), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n545), .A2(new_n455), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n546), .B1(new_n584), .B2(G190), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n583), .A2(G200), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n582), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n424), .A2(new_n520), .A3(new_n551), .A4(new_n587), .ZN(new_n588));
  XNOR2_X1  g0388(.A(new_n588), .B(KEYINPUT80), .ZN(G372));
  AND2_X1   g0389(.A1(new_n516), .A2(new_n519), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT81), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n578), .B1(new_n581), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n561), .A2(G200), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n571), .A2(new_n254), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n594), .A2(new_n580), .A3(new_n563), .ZN(new_n595));
  AOI21_X1  g0395(.A(KEYINPUT81), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n577), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n590), .A2(new_n550), .A3(new_n489), .A4(new_n598), .ZN(new_n599));
  XOR2_X1   g0399(.A(new_n577), .B(KEYINPUT82), .Z(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT83), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT26), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n602), .B(new_n603), .C1(new_n516), .C2(new_n597), .ZN(new_n604));
  INV_X1    g0404(.A(new_n582), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n455), .A2(new_n498), .A3(new_n499), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n513), .B1(new_n606), .B2(new_n319), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n605), .A2(KEYINPUT26), .A3(new_n515), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n593), .A2(new_n595), .A3(KEYINPUT81), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n581), .A2(new_n591), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(new_n611), .A3(new_n578), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n607), .A2(new_n612), .A3(new_n515), .A4(new_n577), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n602), .B1(new_n613), .B2(new_n603), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n599), .B(new_n601), .C1(new_n609), .C2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n424), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n303), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT84), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n398), .A2(new_n618), .A3(new_n408), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n618), .B1(new_n398), .B2(new_n408), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n410), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n409), .A2(KEYINPUT84), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n398), .A2(new_n618), .A3(new_n408), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n622), .A2(KEYINPUT18), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n344), .A2(new_n362), .B1(new_n340), .B2(new_n325), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n419), .A2(new_n420), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n297), .A2(new_n299), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n617), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n616), .A2(new_n630), .ZN(G369));
  NAND2_X1  g0431(.A1(new_n549), .A2(new_n547), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n548), .B1(new_n583), .B2(new_n534), .ZN(new_n633));
  XNOR2_X1  g0433(.A(KEYINPUT85), .B(KEYINPUT27), .ZN(new_n634));
  INV_X1    g0434(.A(G13), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(G20), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  OR3_X1    g0437(.A1(new_n634), .A2(new_n637), .A3(G1), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n634), .B1(new_n637), .B2(G1), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(G213), .A3(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(G343), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n546), .ZN(new_n643));
  OR3_X1    g0443(.A1(new_n632), .A2(new_n633), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n544), .A2(new_n547), .A3(new_n549), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n643), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n585), .A2(new_n586), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n644), .A2(new_n646), .A3(G330), .A4(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n642), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n521), .A2(new_n524), .A3(new_n525), .A4(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n486), .A2(new_n649), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n524), .B1(new_n488), .B2(G190), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n442), .A2(new_n455), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(G200), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n651), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n526), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n650), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n648), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n650), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n649), .B1(new_n632), .B2(new_n633), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(KEYINPUT86), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT86), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n663), .B(new_n649), .C1(new_n632), .C2(new_n633), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n524), .A2(new_n642), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n489), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n660), .B1(new_n526), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n660), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n659), .A2(new_n669), .ZN(G399));
  INV_X1    g0470(.A(new_n220), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G41), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n567), .A2(G116), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G1), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n231), .B2(new_n673), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT28), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n550), .A2(new_n598), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n516), .A2(new_n489), .A3(new_n519), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n601), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n613), .A2(KEYINPUT26), .ZN(new_n681));
  INV_X1    g0481(.A(new_n516), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n682), .A2(new_n603), .A3(new_n605), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n649), .B1(new_n680), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(KEYINPUT29), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n545), .A2(G179), .A3(new_n455), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT87), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n545), .A2(KEYINPUT87), .A3(G179), .A4(new_n455), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n436), .A2(new_n441), .A3(new_n575), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n606), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT30), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n689), .A2(new_n692), .A3(KEYINPUT30), .A4(new_n690), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n575), .A2(G179), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n583), .A2(new_n653), .A3(new_n606), .A4(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n642), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n551), .A2(new_n520), .A3(new_n587), .A4(new_n649), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT31), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n699), .A2(new_n703), .A3(new_n642), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n702), .A2(G330), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT29), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n615), .A2(new_n706), .A3(new_n649), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n686), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n677), .B1(new_n709), .B2(G1), .ZN(G364));
  AOI21_X1  g0510(.A(new_n205), .B1(new_n636), .B2(G45), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n672), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n671), .A2(new_n383), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G355), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(G116), .B2(new_n220), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n671), .A2(new_n286), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n718), .B1(new_n278), .B2(new_n232), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n245), .A2(new_n278), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n716), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(G13), .A2(G33), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G20), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n225), .B1(G20), .B2(new_n319), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n713), .B1(new_n721), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(G190), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n206), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n300), .A2(G200), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(G58), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n286), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n206), .A2(G190), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G179), .A2(G200), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(G159), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XOR2_X1   g0539(.A(new_n739), .B(KEYINPUT32), .Z(new_n740));
  AOI21_X1  g0540(.A(new_n206), .B1(new_n736), .B2(G190), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI211_X1 g0542(.A(new_n734), .B(new_n740), .C1(G97), .C2(new_n742), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n206), .A2(new_n300), .A3(new_n294), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n744), .A2(KEYINPUT89), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(KEYINPUT89), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n745), .A2(G190), .A3(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n745), .A2(new_n729), .A3(new_n746), .ZN(new_n748));
  OAI221_X1 g0548(.A(new_n743), .B1(new_n210), .B2(new_n747), .C1(new_n388), .C2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT88), .ZN(new_n750));
  AND3_X1   g0550(.A1(new_n731), .A2(new_n735), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n750), .B1(new_n731), .B2(new_n735), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n300), .A2(KEYINPUT90), .A3(G200), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(KEYINPUT90), .B1(new_n300), .B2(G200), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n735), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n753), .A2(G77), .B1(new_n759), .B2(G107), .ZN(new_n760));
  INV_X1    g0560(.A(new_n757), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n730), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n760), .B1(new_n212), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G303), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n383), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT91), .Z(new_n766));
  INV_X1    g0566(.A(new_n747), .ZN(new_n767));
  INV_X1    g0567(.A(new_n748), .ZN(new_n768));
  XNOR2_X1  g0568(.A(KEYINPUT33), .B(G317), .ZN(new_n769));
  AOI22_X1  g0569(.A1(G326), .A2(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n753), .A2(G311), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n759), .A2(G283), .ZN(new_n772));
  INV_X1    g0572(.A(G322), .ZN(new_n773));
  INV_X1    g0573(.A(G329), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n732), .A2(new_n773), .B1(new_n737), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(G294), .B2(new_n742), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n770), .A2(new_n771), .A3(new_n772), .A4(new_n776), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n749), .A2(new_n763), .B1(new_n766), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n728), .B1(new_n778), .B2(new_n725), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n644), .A2(new_n647), .A3(new_n646), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(new_n724), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT92), .Z(new_n783));
  INV_X1    g0583(.A(G330), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n713), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n785), .A2(new_n648), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n783), .A2(new_n787), .ZN(G396));
  NAND2_X1  g0588(.A1(new_n358), .A2(G190), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n349), .A2(new_n351), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(new_n347), .B2(new_n254), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n366), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n352), .A2(new_n642), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n791), .B1(new_n365), .B2(new_n319), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n792), .A2(new_n793), .B1(new_n360), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n794), .A2(new_n360), .A3(new_n649), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(KEYINPUT96), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT96), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n649), .A2(new_n791), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(new_n367), .B2(new_n366), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n799), .B(new_n796), .C1(new_n801), .C2(new_n362), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n609), .A2(new_n614), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n649), .B(new_n803), .C1(new_n804), .C2(new_n680), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT97), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n615), .A2(KEYINPUT97), .A3(new_n649), .A4(new_n803), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n632), .A2(new_n633), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n597), .B1(new_n810), .B2(new_n526), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n600), .B1(new_n811), .B2(new_n520), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n603), .B1(new_n516), .B2(new_n597), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(KEYINPUT83), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n814), .A2(new_n608), .A3(new_n604), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n642), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n809), .B1(new_n816), .B2(new_n803), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(new_n705), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n713), .B1(new_n817), .B2(new_n705), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n798), .A2(new_n802), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n722), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n725), .A2(new_n722), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n713), .B1(new_n824), .B2(G77), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n767), .A2(G303), .B1(G116), .B2(new_n753), .ZN(new_n826));
  XOR2_X1   g0626(.A(KEYINPUT93), .B(G283), .Z(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n826), .B1(new_n748), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT94), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n732), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n286), .B1(new_n832), .B2(G294), .ZN(new_n833));
  INV_X1    g0633(.A(G311), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n833), .B1(new_n503), .B2(new_n741), .C1(new_n834), .C2(new_n737), .ZN(new_n835));
  INV_X1    g0635(.A(new_n759), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n836), .A2(new_n212), .B1(new_n762), .B2(new_n356), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n831), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n830), .B2(new_n829), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n753), .A2(G159), .B1(G143), .B2(new_n832), .ZN(new_n840));
  INV_X1    g0640(.A(G137), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n840), .B1(new_n841), .B2(new_n747), .C1(new_n257), .C2(new_n748), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT95), .Z(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(KEYINPUT34), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n836), .A2(new_n388), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(G132), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n286), .B1(new_n741), .B2(new_n733), .C1(new_n847), .C2(new_n737), .ZN(new_n848));
  INV_X1    g0648(.A(new_n762), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n848), .B1(new_n849), .B2(G50), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n844), .A2(new_n846), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n843), .A2(KEYINPUT34), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n839), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n825), .B1(new_n853), .B2(new_n725), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n819), .A2(new_n820), .B1(new_n822), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(G384));
  OAI211_X1 g0656(.A(new_n228), .B(G116), .C1(KEYINPUT35), .C2(new_n509), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(KEYINPUT35), .B2(new_n509), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n858), .B(KEYINPUT36), .Z(new_n859));
  OAI21_X1  g0659(.A(G77), .B1(new_n733), .B2(new_n388), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n231), .A2(new_n860), .B1(G50), .B2(new_n388), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n861), .A2(G1), .A3(new_n635), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT98), .ZN(new_n863));
  INV_X1    g0663(.A(new_n640), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n625), .A2(new_n864), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n343), .A2(new_n342), .B1(new_n340), .B2(new_n642), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n325), .A2(new_n340), .A3(KEYINPUT99), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT99), .B1(new_n325), .B2(new_n340), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n325), .A2(new_n340), .A3(new_n642), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n809), .B2(new_n796), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n391), .A2(new_n374), .A3(new_n375), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n266), .B1(new_n874), .B2(KEYINPUT16), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(KEYINPUT16), .B2(new_n874), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n640), .B1(new_n876), .B2(new_n397), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n421), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n408), .A2(new_n864), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n397), .B2(new_n876), .ZN(new_n880));
  INV_X1    g0680(.A(new_n414), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT37), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n398), .A2(new_n864), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n883), .A2(new_n414), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT37), .B1(new_n398), .B2(new_n408), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT100), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n885), .A2(new_n414), .A3(new_n883), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT100), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n882), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n878), .A2(KEYINPUT38), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT38), .B1(new_n878), .B2(new_n890), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n865), .B1(new_n873), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT101), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n867), .A2(new_n868), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n897), .A2(new_n642), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT38), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n415), .A2(new_n418), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n883), .B1(new_n625), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n884), .A2(KEYINPUT100), .A3(new_n885), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n887), .A2(new_n888), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n414), .B(new_n883), .C1(new_n619), .C2(new_n620), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n902), .A2(new_n903), .B1(new_n904), .B2(KEYINPUT37), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n899), .B1(new_n901), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n878), .A2(new_n890), .A3(KEYINPUT38), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n908), .A2(KEYINPUT39), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT39), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n878), .A2(new_n890), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n899), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n910), .B1(new_n912), .B2(new_n907), .ZN(new_n913));
  OR2_X1    g0713(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n895), .A2(new_n896), .B1(new_n898), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT97), .B1(new_n816), .B2(new_n803), .ZN(new_n916));
  AND4_X1   g0716(.A1(KEYINPUT97), .A2(new_n615), .A3(new_n649), .A4(new_n803), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n796), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n918), .A2(new_n894), .A3(new_n871), .ZN(new_n919));
  INV_X1    g0719(.A(new_n865), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n896), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n915), .A2(new_n922), .ZN(new_n923));
  AND3_X1   g0723(.A1(new_n699), .A2(new_n703), .A3(new_n642), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n703), .B1(new_n699), .B2(new_n642), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n924), .B1(new_n701), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n821), .B1(new_n869), .B2(new_n870), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n926), .B(new_n927), .C1(new_n891), .C2(new_n892), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT40), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n927), .A2(new_n702), .A3(new_n704), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n929), .B1(new_n906), .B2(new_n907), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n930), .A2(G330), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n424), .A2(G330), .A3(new_n926), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n928), .A2(new_n929), .B1(new_n931), .B2(new_n932), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n937), .A2(new_n424), .A3(new_n926), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n923), .B(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n686), .A2(new_n707), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT102), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n941), .A2(new_n942), .A3(new_n424), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n942), .B1(new_n941), .B2(new_n424), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n630), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT103), .Z(new_n947));
  NAND2_X1  g0747(.A1(new_n940), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n205), .B2(new_n636), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n940), .A2(new_n947), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n859), .B(new_n863), .C1(new_n949), .C2(new_n950), .ZN(G367));
  NOR2_X1   g0751(.A1(new_n718), .A2(new_n241), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n726), .B1(new_n220), .B2(new_n346), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n713), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n836), .A2(new_n503), .ZN(new_n955));
  INV_X1    g0755(.A(new_n737), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n286), .B(new_n955), .C1(G317), .C2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT112), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n762), .A2(new_n476), .ZN(new_n960));
  INV_X1    g0760(.A(G294), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n960), .A2(KEYINPUT46), .B1(new_n961), .B2(new_n748), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(KEYINPUT46), .B2(new_n960), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n957), .A2(new_n958), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n732), .A2(new_n764), .B1(new_n741), .B2(new_n356), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n747), .A2(new_n834), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n965), .B(new_n966), .C1(new_n753), .C2(new_n827), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n959), .A2(new_n963), .A3(new_n964), .A4(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n753), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n969), .A2(new_n210), .B1(new_n748), .B2(new_n738), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n970), .A2(KEYINPUT113), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(KEYINPUT113), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n767), .A2(G143), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n836), .A2(new_n202), .B1(new_n762), .B2(new_n733), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n383), .B1(new_n832), .B2(G150), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n742), .A2(G68), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n975), .B(new_n976), .C1(new_n841), .C2(new_n737), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n971), .A2(new_n972), .A3(new_n973), .A4(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(KEYINPUT47), .B1(new_n968), .B2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n725), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n968), .A2(KEYINPUT47), .A3(new_n979), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n954), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n724), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n649), .A2(new_n595), .ZN(new_n986));
  MUX2_X1   g0786(.A(new_n598), .B(new_n600), .S(new_n986), .Z(new_n987));
  OAI21_X1  g0787(.A(new_n984), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT111), .ZN(new_n989));
  INV_X1    g0789(.A(new_n664), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n663), .B1(new_n645), .B2(new_n649), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n668), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AND3_X1   g0792(.A1(new_n992), .A2(KEYINPUT110), .A3(new_n648), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n648), .B1(new_n992), .B2(KEYINPUT110), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n665), .A2(new_n668), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  NOR3_X1   g0796(.A1(new_n993), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n648), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n657), .B1(new_n664), .B2(new_n662), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT110), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n992), .A2(KEYINPUT110), .A3(new_n648), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n995), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n997), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n989), .B1(new_n1004), .B2(new_n708), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n514), .A2(new_n642), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n516), .A2(new_n519), .A3(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n607), .A2(new_n515), .A3(new_n642), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n992), .A2(new_n650), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(KEYINPUT109), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT109), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n669), .A2(new_n1012), .A3(new_n1009), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1011), .A2(KEYINPUT45), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT44), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n669), .B2(new_n1009), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1009), .ZN(new_n1017));
  OAI211_X1 g0817(.A(KEYINPUT44), .B(new_n1017), .C1(new_n999), .C2(new_n660), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1014), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(KEYINPUT45), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n658), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT45), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1025), .A2(new_n659), .A3(new_n1019), .A4(new_n1014), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n996), .B1(new_n993), .B2(new_n994), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1001), .A2(new_n995), .A3(new_n1002), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n709), .A2(new_n1029), .A3(KEYINPUT111), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1005), .A2(new_n1022), .A3(new_n1026), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n709), .ZN(new_n1032));
  XOR2_X1   g0832(.A(KEYINPUT108), .B(KEYINPUT41), .Z(new_n1033));
  XOR2_X1   g0833(.A(new_n672), .B(new_n1033), .Z(new_n1034));
  AOI21_X1  g0834(.A(new_n712), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT42), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n999), .B2(new_n1009), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n665), .A2(new_n1036), .A3(new_n668), .A4(new_n1009), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT106), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n999), .A2(KEYINPUT106), .A3(new_n1036), .A4(new_n1009), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1037), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT104), .ZN(new_n1043));
  AND3_X1   g0843(.A1(new_n1007), .A2(new_n1043), .A3(new_n1008), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1043), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1045));
  NOR3_X1   g0845(.A1(new_n1044), .A2(new_n1045), .A3(new_n526), .ZN(new_n1046));
  OAI21_X1  g0846(.A(KEYINPUT105), .B1(new_n1046), .B2(new_n682), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1045), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1007), .A2(new_n1043), .A3(new_n1008), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1048), .A2(new_n656), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT105), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1050), .A2(new_n1051), .A3(new_n516), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1047), .A2(new_n649), .A3(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n987), .A2(KEYINPUT43), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1042), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT107), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1042), .A2(new_n1053), .A3(KEYINPUT107), .A4(new_n1054), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1042), .A2(new_n1053), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n987), .B(KEYINPUT43), .Z(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1057), .A2(new_n1058), .A3(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n659), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1062), .B(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n988), .B1(new_n1035), .B2(new_n1067), .ZN(G387));
  NAND2_X1  g0868(.A1(new_n1004), .A2(new_n708), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n709), .A2(new_n1029), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1069), .A2(new_n672), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n718), .B1(new_n238), .B2(G45), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n674), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1072), .B1(new_n1073), .B2(new_n714), .ZN(new_n1074));
  AOI21_X1  g0874(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n264), .A2(new_n210), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n674), .B(new_n1075), .C1(new_n1076), .C2(KEYINPUT50), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(KEYINPUT50), .B2(new_n1076), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n1074), .A2(new_n1078), .B1(G107), .B2(new_n220), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n786), .B1(new_n1079), .B2(new_n726), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT114), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n762), .A2(new_n202), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1082), .B(new_n955), .C1(G68), .C2(new_n753), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n741), .A2(new_n346), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n286), .B1(new_n737), .B2(new_n257), .C1(new_n732), .C2(new_n210), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1084), .B(new_n1085), .C1(new_n768), .C2(new_n264), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1083), .B(new_n1086), .C1(new_n738), .C2(new_n747), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT115), .Z(new_n1088));
  AOI21_X1  g0888(.A(new_n286), .B1(new_n956), .B2(G326), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n753), .A2(G303), .B1(G317), .B2(new_n832), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1090), .B1(new_n834), .B2(new_n748), .C1(new_n773), .C2(new_n747), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT48), .Z(new_n1092));
  OAI22_X1  g0892(.A1(new_n762), .A2(new_n961), .B1(new_n741), .B2(new_n828), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1089), .B1(new_n476), .B2(new_n836), .C1(new_n1094), .C2(KEYINPUT49), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n1094), .A2(KEYINPUT49), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1088), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1081), .B1(new_n1097), .B2(new_n725), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n668), .B2(new_n985), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1071), .B(new_n1099), .C1(new_n711), .C2(new_n1004), .ZN(G393));
  NAND3_X1  g0900(.A1(new_n1022), .A2(new_n1026), .A3(new_n712), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n718), .A2(new_n249), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n726), .B1(new_n503), .B2(new_n220), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n713), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n767), .A2(G317), .B1(G311), .B2(new_n832), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(KEYINPUT117), .B(KEYINPUT52), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n768), .A2(G303), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n383), .B1(new_n741), .B2(new_n476), .C1(new_n773), .C2(new_n737), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G107), .B2(new_n759), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n849), .A2(new_n827), .B1(G294), .B2(new_n753), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1107), .A2(new_n1108), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n747), .A2(new_n257), .B1(new_n732), .B2(new_n738), .ZN(new_n1114));
  XOR2_X1   g0914(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n1115));
  NOR2_X1   g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n768), .A2(G50), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n741), .A2(new_n202), .ZN(new_n1119));
  INV_X1    g0919(.A(G143), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n286), .B1(new_n737), .B2(new_n1120), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1119), .B(new_n1121), .C1(new_n759), .C2(G87), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n849), .A2(G68), .B1(new_n264), .B2(new_n753), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1117), .A2(new_n1118), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n1112), .A2(new_n1113), .B1(new_n1116), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1104), .B1(new_n1125), .B2(new_n725), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n1063), .B2(new_n985), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1031), .A2(new_n672), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1022), .A2(new_n1026), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1129), .A2(new_n1070), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1101), .B(new_n1127), .C1(new_n1128), .C2(new_n1130), .ZN(G390));
  OAI21_X1  g0931(.A(new_n713), .B1(new_n824), .B2(new_n264), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n849), .A2(G150), .ZN(new_n1133));
  OR2_X1    g0933(.A1(new_n1133), .A2(KEYINPUT53), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1133), .A2(KEYINPUT53), .B1(G137), .B2(new_n768), .ZN(new_n1135));
  XOR2_X1   g0935(.A(KEYINPUT54), .B(G143), .Z(new_n1136));
  NAND2_X1  g0936(.A1(new_n753), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n383), .B1(new_n956), .B2(G125), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n738), .B2(new_n741), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(G50), .B2(new_n759), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1134), .A2(new_n1135), .A3(new_n1137), .A4(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(G128), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n747), .A2(new_n1142), .B1(new_n732), .B2(new_n847), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT118), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n383), .B1(new_n737), .B2(new_n961), .C1(new_n732), .C2(new_n476), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1119), .B(new_n1145), .C1(new_n767), .C2(G283), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n356), .B2(new_n748), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n846), .B1(new_n212), .B2(new_n762), .C1(new_n503), .C2(new_n969), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n1141), .A2(new_n1144), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1132), .B1(new_n1149), .B2(new_n725), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n914), .B2(new_n723), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n898), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n908), .A2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n649), .B(new_n803), .C1(new_n680), .C2(new_n684), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n872), .B1(new_n796), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n898), .B1(new_n918), .B2(new_n871), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1157), .B1(new_n1158), .B2(new_n914), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n926), .A2(G330), .A3(new_n927), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n797), .B1(new_n807), .B2(new_n808), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1152), .B1(new_n1163), .B2(new_n872), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n909), .A2(new_n913), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1166), .A2(new_n1160), .A3(new_n1157), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1162), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1151), .B1(new_n1168), .B2(new_n711), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n872), .B1(new_n705), .B2(new_n821), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n796), .A2(new_n809), .B1(new_n1170), .B2(new_n1160), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1154), .A2(new_n796), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1170), .A2(new_n1160), .A3(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n630), .B(new_n935), .C1(new_n943), .C2(new_n944), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n673), .B1(new_n1168), .B2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1162), .A2(new_n1167), .A3(new_n1176), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1169), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(G378));
  INV_X1    g0981(.A(KEYINPUT57), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1160), .B1(new_n1166), .B2(new_n1157), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1161), .B(new_n1156), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1175), .B1(new_n1185), .B2(new_n1176), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT120), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n304), .B(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n267), .A2(new_n864), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n304), .B(KEYINPUT120), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1191), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1188), .B1(new_n1192), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1197), .A2(new_n1198), .A3(new_n1187), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1196), .A2(new_n1199), .ZN(new_n1200));
  AND4_X1   g1000(.A1(G330), .A2(new_n930), .A3(new_n1200), .A4(new_n933), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1200), .B1(new_n937), .B2(G330), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1203), .A2(new_n915), .A3(new_n922), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1200), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n934), .A2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n937), .A2(G330), .A3(new_n1200), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n919), .A2(new_n896), .A3(new_n920), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n914), .A2(new_n898), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1208), .B1(new_n1211), .B2(new_n921), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1204), .A2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1182), .B1(new_n1186), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1175), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1179), .A2(new_n1215), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1216), .A2(KEYINPUT57), .A3(new_n1204), .A4(new_n1212), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1214), .A2(new_n672), .A3(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n786), .B1(new_n210), .B2(new_n823), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n976), .B1(new_n747), .B2(new_n476), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT119), .Z(new_n1221));
  NOR2_X1   g1021(.A1(new_n969), .A2(new_n346), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n836), .A2(new_n733), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n286), .A2(G41), .ZN(new_n1224));
  INV_X1    g1024(.A(G283), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1224), .B1(new_n1225), .B2(new_n737), .C1(new_n356), .C2(new_n732), .ZN(new_n1226));
  NOR4_X1   g1026(.A1(new_n1222), .A2(new_n1223), .A3(new_n1082), .A4(new_n1226), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1221), .B(new_n1227), .C1(new_n503), .C2(new_n748), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT58), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(G125), .A2(new_n767), .B1(new_n768), .B2(G132), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n732), .A2(new_n1142), .B1(new_n741), .B2(new_n257), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n849), .B2(new_n1136), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1231), .B(new_n1233), .C1(new_n841), .C2(new_n969), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1234), .A2(KEYINPUT59), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(KEYINPUT59), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n759), .A2(G159), .ZN(new_n1237));
  AOI211_X1 g1037(.A(G33), .B(G41), .C1(new_n956), .C2(G124), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1230), .B1(new_n1235), .B2(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1241));
  AOI211_X1 g1041(.A(G50), .B(new_n1224), .C1(new_n379), .C2(new_n277), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n1219), .B1(new_n981), .B2(new_n1243), .C1(new_n1205), .C2(new_n723), .ZN(new_n1244));
  XOR2_X1   g1044(.A(new_n1244), .B(KEYINPUT121), .Z(new_n1245));
  INV_X1    g1045(.A(new_n1213), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1245), .B1(new_n1246), .B2(new_n712), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1218), .A2(new_n1247), .ZN(G375));
  INV_X1    g1048(.A(new_n1174), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n872), .A2(new_n722), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n713), .B1(new_n824), .B2(G68), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT122), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n286), .B1(new_n732), .B2(new_n841), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n1253), .B(new_n1223), .C1(G50), .C2(new_n742), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(G132), .A2(new_n767), .B1(new_n768), .B2(new_n1136), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1254), .B(new_n1255), .C1(new_n257), .C2(new_n969), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n762), .A2(new_n738), .B1(new_n1142), .B2(new_n737), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1257), .B(KEYINPUT124), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n969), .A2(new_n356), .B1(new_n748), .B2(new_n476), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT123), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n836), .A2(new_n202), .B1(new_n762), .B2(new_n503), .ZN(new_n1262));
  OAI221_X1 g1062(.A(new_n383), .B1(new_n737), .B2(new_n764), .C1(new_n732), .C2(new_n1225), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(new_n1262), .A2(new_n1263), .A3(new_n1084), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1264), .B(new_n1265), .C1(new_n961), .C2(new_n747), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n1256), .A2(new_n1258), .B1(new_n1261), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1252), .B1(new_n1267), .B2(new_n725), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1249), .A2(new_n712), .B1(new_n1250), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1177), .A2(new_n1034), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1249), .A2(new_n1215), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1269), .B1(new_n1270), .B2(new_n1271), .ZN(G381));
  NAND3_X1  g1072(.A1(new_n1218), .A2(new_n1180), .A3(new_n1247), .ZN(new_n1273));
  OR2_X1    g1073(.A1(G393), .A2(G396), .ZN(new_n1274));
  OR4_X1    g1074(.A1(G384), .A2(G381), .A3(G390), .A4(new_n1274), .ZN(new_n1275));
  OR3_X1    g1075(.A1(new_n1273), .A2(new_n1275), .A3(G387), .ZN(G407));
  OAI211_X1 g1076(.A(G407), .B(G213), .C1(G343), .C2(new_n1273), .ZN(G409));
  INV_X1    g1077(.A(KEYINPUT61), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n641), .A2(G213), .A3(G2897), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1271), .A2(KEYINPUT60), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT60), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n1249), .B2(new_n1215), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1281), .A2(new_n672), .A3(new_n1177), .A4(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1269), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n855), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1285), .A2(new_n855), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1280), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1288), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1290), .A2(new_n1286), .A3(new_n1279), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1218), .A2(G378), .A3(new_n1247), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1246), .A2(new_n1034), .A3(new_n1216), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1247), .A2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1180), .ZN(new_n1296));
  AOI22_X1  g1096(.A1(new_n1293), .A2(new_n1296), .B1(G213), .B2(new_n641), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1278), .B1(new_n1292), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1297), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT63), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(G393), .B(G396), .ZN(new_n1304));
  AOI22_X1  g1104(.A1(new_n1055), .A2(new_n1056), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1065), .B1(new_n1305), .B2(new_n1058), .ZN(new_n1306));
  AND4_X1   g1106(.A1(new_n1065), .A2(new_n1057), .A3(new_n1058), .A4(new_n1061), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1034), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1309), .B1(new_n1031), .B2(new_n709), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1308), .B1(new_n1310), .B2(new_n712), .ZN(new_n1311));
  AOI21_X1  g1111(.A(G390), .B1(new_n1311), .B2(new_n988), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1304), .B1(new_n1312), .B2(KEYINPUT125), .ZN(new_n1313));
  INV_X1    g1113(.A(G390), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(G387), .A2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1311), .A2(new_n988), .A3(G390), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1313), .B1(new_n1317), .B2(KEYINPUT125), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT126), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1311), .A2(new_n988), .A3(G390), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1320), .A2(new_n1312), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1319), .B1(new_n1321), .B2(new_n1304), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1315), .A2(new_n1319), .A3(new_n1316), .A4(new_n1304), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1318), .B1(new_n1322), .B2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1297), .A2(KEYINPUT63), .A3(new_n1300), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1299), .A2(new_n1303), .A3(new_n1325), .A4(new_n1326), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1301), .A2(KEYINPUT62), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT62), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1329), .B1(new_n1297), .B2(new_n1300), .ZN(new_n1330));
  NOR3_X1   g1130(.A1(new_n1328), .A2(new_n1298), .A3(new_n1330), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1327), .B1(new_n1331), .B2(new_n1325), .ZN(G405));
  INV_X1    g1132(.A(new_n1293), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1333), .A2(KEYINPUT127), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1315), .A2(new_n1316), .A3(new_n1304), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(KEYINPUT126), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n1323), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(G375), .A2(new_n1180), .ZN(new_n1338));
  AND3_X1   g1138(.A1(new_n1337), .A2(new_n1318), .A3(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1338), .B1(new_n1337), .B2(new_n1318), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1334), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1338), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1325), .A2(new_n1342), .ZN(new_n1343));
  OR2_X1    g1143(.A1(new_n1333), .A2(KEYINPUT127), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1337), .A2(new_n1338), .A3(new_n1318), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1343), .A2(new_n1344), .A3(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1300), .ZN(new_n1347));
  AND3_X1   g1147(.A1(new_n1341), .A2(new_n1346), .A3(new_n1347), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1347), .B1(new_n1341), .B2(new_n1346), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n1348), .A2(new_n1349), .ZN(G402));
endmodule


