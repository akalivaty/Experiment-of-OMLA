//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n449, new_n450, new_n452, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n570, new_n572, new_n573, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n631, new_n632,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1180;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT68), .ZN(new_n449));
  AND2_X1   g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n449), .B(new_n450), .ZN(G223));
  NAND2_X1  g026(.A1(new_n450), .A2(G567), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT69), .Z(G234));
  NAND2_X1  g028(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n456), .A2(G2106), .ZN(new_n461));
  INV_X1    g036(.A(G567), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(new_n457), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  AND3_X1   g043(.A1(KEYINPUT71), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(KEYINPUT3), .B1(KEYINPUT71), .B2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n467), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT72), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT72), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n475), .B(new_n467), .C1(new_n471), .C2(new_n472), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT70), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n479), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n478), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g061(.A1(G113), .A2(G2104), .ZN(new_n487));
  OAI21_X1  g062(.A(G2105), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n477), .A2(new_n488), .ZN(G160));
  NOR2_X1   g064(.A1(new_n469), .A2(new_n470), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(new_n468), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G124), .ZN(new_n492));
  INV_X1    g067(.A(new_n471), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G136), .ZN(new_n494));
  NOR2_X1   g069(.A1(G100), .A2(G2105), .ZN(new_n495));
  XOR2_X1   g070(.A(new_n495), .B(KEYINPUT73), .Z(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(new_n468), .B2(G112), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n492), .B(new_n494), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  XNOR2_X1  g073(.A(new_n498), .B(KEYINPUT74), .ZN(G162));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR3_X1   g075(.A1(new_n500), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n501));
  AND3_X1   g076(.A1(new_n479), .A2(new_n481), .A3(new_n484), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n484), .B1(new_n479), .B2(new_n481), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT76), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT4), .B1(new_n471), .B2(new_n500), .ZN(new_n507));
  OAI211_X1 g082(.A(KEYINPUT76), .B(new_n501), .C1(new_n502), .C2(new_n503), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n468), .A2(G114), .ZN(new_n510));
  XOR2_X1   g085(.A(new_n510), .B(KEYINPUT75), .Z(new_n511));
  OAI21_X1  g086(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n511), .A2(new_n513), .B1(G126), .B2(new_n491), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(G164));
  OR2_X1    g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n519), .A2(G50), .A3(G543), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT77), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n520), .B(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT5), .ZN(new_n523));
  OAI21_X1  g098(.A(KEYINPUT78), .B1(new_n523), .B2(G543), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT78), .ZN(new_n525));
  INV_X1    g100(.A(G543), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n525), .A2(new_n526), .A3(KEYINPUT5), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n523), .A2(G543), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n519), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  XOR2_X1   g107(.A(KEYINPUT79), .B(G88), .Z(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n528), .A2(new_n529), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n535), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G651), .ZN(new_n537));
  OAI211_X1 g112(.A(new_n522), .B(new_n534), .C1(new_n536), .C2(new_n537), .ZN(G303));
  INV_X1    g113(.A(G303), .ZN(G166));
  INV_X1    g114(.A(KEYINPUT80), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n519), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n517), .A2(KEYINPUT80), .A3(new_n518), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n541), .A2(G543), .A3(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G51), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n532), .A2(G89), .ZN(new_n546));
  NAND3_X1  g121(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT7), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n535), .A2(G63), .A3(G651), .ZN(new_n549));
  NAND4_X1  g124(.A1(new_n545), .A2(new_n546), .A3(new_n548), .A4(new_n549), .ZN(G286));
  INV_X1    g125(.A(G286), .ZN(G168));
  AOI22_X1  g126(.A1(new_n535), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n537), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n535), .A2(new_n519), .ZN(new_n554));
  INV_X1    g129(.A(G90), .ZN(new_n555));
  INV_X1    g130(.A(G52), .ZN(new_n556));
  OAI22_X1  g131(.A1(new_n554), .A2(new_n555), .B1(new_n556), .B2(new_n543), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n553), .A2(new_n557), .ZN(G301));
  INV_X1    g133(.A(G301), .ZN(G171));
  NAND4_X1  g134(.A1(new_n541), .A2(G43), .A3(G543), .A4(new_n542), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n528), .A2(G81), .A3(new_n529), .A4(new_n519), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n560), .A2(KEYINPUT81), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(KEYINPUT81), .B1(new_n560), .B2(new_n561), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(G68), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G56), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n530), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G651), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n564), .A2(G860), .A3(new_n568), .ZN(G153));
  AND3_X1   g144(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G36), .ZN(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n570), .A2(new_n573), .ZN(G188));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  XOR2_X1   g150(.A(new_n575), .B(KEYINPUT84), .Z(new_n576));
  INV_X1    g151(.A(G65), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n530), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(KEYINPUT85), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT85), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n580), .B(new_n576), .C1(new_n530), .C2(new_n577), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(G651), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g157(.A(KEYINPUT83), .B1(KEYINPUT82), .B2(KEYINPUT9), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n583), .B1(KEYINPUT83), .B2(KEYINPUT9), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n544), .A2(G53), .A3(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(G53), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n583), .B1(new_n543), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n532), .A2(G91), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n582), .A2(new_n585), .A3(new_n587), .A4(new_n588), .ZN(G299));
  NAND4_X1  g164(.A1(new_n528), .A2(G87), .A3(new_n529), .A4(new_n519), .ZN(new_n590));
  INV_X1    g165(.A(G49), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n543), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(G74), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n537), .B1(new_n530), .B2(new_n593), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n592), .A2(new_n594), .ZN(G288));
  NAND3_X1  g170(.A1(new_n528), .A2(G61), .A3(new_n529), .ZN(new_n596));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n537), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n528), .A2(G86), .A3(new_n529), .ZN(new_n600));
  NAND2_X1  g175(.A1(G48), .A2(G543), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n531), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n599), .A2(new_n603), .ZN(G305));
  AOI22_X1  g179(.A1(new_n544), .A2(G47), .B1(new_n532), .B2(G85), .ZN(new_n605));
  NAND2_X1  g180(.A1(G72), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G60), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n530), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT86), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n608), .A2(new_n609), .A3(G651), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n609), .B1(new_n608), .B2(G651), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n611), .B2(new_n612), .ZN(G290));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n614));
  INV_X1    g189(.A(G92), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n554), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n532), .A2(KEYINPUT10), .A3(G92), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  INV_X1    g194(.A(G66), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n530), .B2(new_n620), .ZN(new_n621));
  AOI22_X1  g196(.A1(G54), .A2(new_n544), .B1(new_n621), .B2(G651), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(G868), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G171), .B2(new_n624), .ZN(G321));
  XOR2_X1   g201(.A(G321), .B(KEYINPUT87), .Z(G284));
  NAND2_X1  g202(.A1(G299), .A2(new_n624), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(new_n624), .B2(G168), .ZN(G297));
  OAI21_X1  g204(.A(new_n628), .B1(new_n624), .B2(G168), .ZN(G280));
  INV_X1    g205(.A(new_n623), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT88), .B(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(G860), .B2(new_n632), .ZN(G148));
  OAI21_X1  g208(.A(new_n568), .B1(new_n562), .B2(new_n563), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n631), .A2(new_n632), .ZN(new_n635));
  MUX2_X1   g210(.A(new_n634), .B(new_n635), .S(G868), .Z(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g212(.A1(new_n483), .A2(new_n485), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(new_n466), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT12), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2100), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n640), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n491), .A2(G123), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n493), .A2(G135), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n468), .A2(G111), .ZN(new_n646));
  OAI21_X1  g221(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n644), .B(new_n645), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT90), .B(G2096), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n643), .A2(new_n650), .ZN(G156));
  XNOR2_X1  g226(.A(G2427), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2430), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(KEYINPUT14), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT91), .Z(new_n665));
  INV_X1    g240(.A(G14), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n662), .B2(new_n663), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(G401));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n670), .ZN(new_n673));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(KEYINPUT17), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n670), .A2(new_n671), .ZN(new_n677));
  OAI221_X1 g252(.A(new_n672), .B1(new_n671), .B2(new_n675), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n672), .A2(new_n674), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT92), .B(KEYINPUT18), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT93), .ZN(new_n683));
  XOR2_X1   g258(.A(G2096), .B(G2100), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(G1971), .B(G1976), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  XOR2_X1   g262(.A(G1956), .B(G2474), .Z(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  AND2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT95), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT94), .B(KEYINPUT20), .Z(new_n693));
  OR2_X1    g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n692), .A2(new_n693), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n688), .A2(new_n689), .ZN(new_n696));
  NOR3_X1   g271(.A1(new_n687), .A2(new_n690), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n687), .B2(new_n696), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n694), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(G1991), .B(G1996), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1981), .B(G1986), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n701), .A2(new_n703), .ZN(new_n708));
  OR3_X1    g283(.A1(new_n705), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n707), .B1(new_n705), .B2(new_n708), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(G229));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G21), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G168), .B2(new_n713), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT106), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G1966), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT107), .Z(new_n718));
  XOR2_X1   g293(.A(KEYINPUT96), .B(G29), .Z(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G26), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT28), .Z(new_n721));
  NAND2_X1  g296(.A1(new_n493), .A2(G140), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT104), .Z(new_n723));
  OAI21_X1  g298(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n724));
  INV_X1    g299(.A(G116), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(G2105), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT105), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G128), .B2(new_n491), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n723), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n721), .B1(new_n729), .B2(G29), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G2067), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT31), .B(G11), .Z(new_n732));
  INV_X1    g307(.A(G28), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n733), .A2(KEYINPUT30), .ZN(new_n734));
  AOI21_X1  g309(.A(G29), .B1(new_n733), .B2(KEYINPUT30), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n732), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G32), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(G29), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n491), .A2(G129), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n493), .A2(G141), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT26), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n743), .A2(new_n744), .B1(G105), .B2(new_n466), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n739), .A2(new_n740), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n738), .B1(new_n746), .B2(G29), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT27), .B(G1996), .ZN(new_n748));
  OAI221_X1 g323(.A(new_n736), .B1(new_n648), .B2(new_n719), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n747), .B2(new_n748), .ZN(new_n750));
  NAND2_X1  g325(.A1(G160), .A2(G29), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT24), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n752), .A2(G34), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(G34), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n719), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2084), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n731), .A2(new_n750), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n713), .A2(G5), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G171), .B2(new_n713), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n760), .A2(G1961), .ZN(new_n761));
  INV_X1    g336(.A(G33), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(G29), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT25), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n493), .A2(G139), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n638), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n769), .B2(new_n468), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n763), .B1(new_n770), .B2(G29), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n772), .A2(G2072), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n760), .A2(G1961), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n772), .A2(G2072), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n761), .A2(new_n773), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n713), .A2(G20), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT23), .Z(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G299), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT108), .B(G1956), .ZN(new_n780));
  AOI211_X1 g355(.A(new_n758), .B(new_n776), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  MUX2_X1   g356(.A(G19), .B(new_n634), .S(G16), .Z(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(G1341), .Z(new_n783));
  INV_X1    g358(.A(new_n719), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n784), .A2(G35), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G162), .B2(new_n784), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT29), .Z(new_n787));
  INV_X1    g362(.A(G2090), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n783), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n788), .B2(new_n787), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n716), .A2(G1966), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n713), .A2(G4), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n631), .B2(new_n713), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT103), .B(G1348), .Z(new_n794));
  XOR2_X1   g369(.A(new_n793), .B(new_n794), .Z(new_n795));
  NOR2_X1   g370(.A1(new_n784), .A2(G27), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G164), .B2(new_n784), .ZN(new_n797));
  INV_X1    g372(.A(G2078), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n779), .B2(new_n780), .ZN(new_n800));
  NOR3_X1   g375(.A1(new_n791), .A2(new_n795), .A3(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n718), .A2(new_n781), .A3(new_n790), .A4(new_n801), .ZN(new_n802));
  OR2_X1    g377(.A1(G16), .A2(G24), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G290), .B2(new_n713), .ZN(new_n804));
  INV_X1    g379(.A(G1986), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n784), .A2(G25), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n491), .A2(G119), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n493), .A2(G131), .ZN(new_n810));
  OR2_X1    g385(.A1(G95), .A2(G2105), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n811), .B(G2104), .C1(G107), .C2(new_n468), .ZN(new_n812));
  AND3_X1   g387(.A1(new_n809), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n808), .B1(new_n813), .B2(new_n784), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT98), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT35), .B(G1991), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT97), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n815), .B(new_n817), .Z(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n805), .B2(new_n804), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n713), .A2(G23), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n592), .A2(new_n594), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(new_n713), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT101), .Z(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT33), .B(G1976), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n713), .A2(G22), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(G166), .B2(new_n713), .ZN(new_n828));
  INV_X1    g403(.A(G1971), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  MUX2_X1   g405(.A(G6), .B(G305), .S(G16), .Z(new_n831));
  XOR2_X1   g406(.A(KEYINPUT32), .B(G1981), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT100), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n831), .B(new_n833), .ZN(new_n834));
  AND4_X1   g409(.A1(new_n825), .A2(new_n826), .A3(new_n830), .A4(new_n834), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT99), .B(KEYINPUT34), .Z(new_n836));
  AOI211_X1 g411(.A(new_n807), .B(new_n819), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT102), .B(KEYINPUT36), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n837), .A2(new_n838), .A3(new_n840), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n802), .B1(new_n842), .B2(new_n843), .ZN(G311));
  INV_X1    g419(.A(G311), .ZN(G150));
  NAND2_X1  g420(.A1(new_n631), .A2(G559), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT38), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n528), .A2(G93), .A3(new_n529), .A4(new_n519), .ZN(new_n848));
  INV_X1    g423(.A(G55), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n543), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n528), .A2(G67), .A3(new_n529), .ZN(new_n851));
  NAND2_X1  g426(.A1(G80), .A2(G543), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n537), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n634), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n850), .A2(new_n853), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n856), .B(new_n568), .C1(new_n563), .C2(new_n562), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n847), .B(new_n858), .Z(new_n859));
  OR2_X1    g434(.A1(new_n859), .A2(KEYINPUT39), .ZN(new_n860));
  INV_X1    g435(.A(G860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(KEYINPUT39), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n856), .A2(new_n861), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT37), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(G145));
  INV_X1    g441(.A(KEYINPUT110), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n491), .A2(G130), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n493), .A2(G142), .ZN(new_n869));
  OR2_X1    g444(.A1(G106), .A2(G2105), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n870), .B(G2104), .C1(G118), .C2(new_n468), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n868), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT109), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n874), .A2(new_n640), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n640), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(new_n876), .A3(new_n813), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n813), .B1(new_n875), .B2(new_n876), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n867), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n879), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n881), .A2(KEYINPUT110), .A3(new_n877), .ZN(new_n882));
  NAND3_X1  g457(.A1(G164), .A2(new_n723), .A3(new_n728), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n729), .A2(new_n515), .ZN(new_n884));
  INV_X1    g459(.A(new_n770), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n746), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n885), .B1(new_n883), .B2(new_n884), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n883), .A2(new_n884), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n770), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n746), .B1(new_n892), .B2(new_n886), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n880), .B(new_n882), .C1(new_n890), .C2(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(KEYINPUT110), .B1(new_n881), .B2(new_n877), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n892), .A2(new_n746), .A3(new_n886), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n888), .B1(new_n887), .B2(new_n889), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(G162), .B(G160), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(new_n648), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n894), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(KEYINPUT111), .B(G37), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT112), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n894), .A2(new_n898), .ZN(new_n905));
  INV_X1    g480(.A(new_n900), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AOI211_X1 g482(.A(KEYINPUT112), .B(new_n900), .C1(new_n894), .C2(new_n898), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n903), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(KEYINPUT113), .B(KEYINPUT40), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n909), .B(new_n910), .ZN(G395));
  INV_X1    g486(.A(KEYINPUT114), .ZN(new_n912));
  NOR2_X1   g487(.A1(G290), .A2(G288), .ZN(new_n913));
  INV_X1    g488(.A(new_n612), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n610), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n821), .B1(new_n915), .B2(new_n605), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n912), .B1(new_n913), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(G290), .A2(G288), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n915), .A2(new_n821), .A3(new_n605), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(KEYINPUT114), .ZN(new_n920));
  XNOR2_X1  g495(.A(G303), .B(G305), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n917), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n921), .A2(KEYINPUT114), .A3(new_n918), .A4(new_n919), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g500(.A(KEYINPUT115), .B(KEYINPUT42), .Z(new_n926));
  OR2_X1    g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n635), .B(new_n858), .ZN(new_n928));
  NAND2_X1  g503(.A1(G299), .A2(new_n623), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n930), .A2(new_n582), .A3(new_n618), .A4(new_n622), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(KEYINPUT41), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT41), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n929), .A2(new_n931), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n933), .B1(new_n928), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n925), .A2(new_n926), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n927), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n938), .B1(new_n927), .B2(new_n939), .ZN(new_n941));
  OAI21_X1  g516(.A(G868), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n854), .A2(new_n624), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(G295));
  INV_X1    g519(.A(KEYINPUT116), .ZN(new_n945));
  XNOR2_X1  g520(.A(G295), .B(new_n945), .ZN(G331));
  INV_X1    g521(.A(KEYINPUT120), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n855), .A2(new_n857), .A3(G301), .ZN(new_n948));
  AOI21_X1  g523(.A(G301), .B1(new_n855), .B2(new_n857), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n948), .A2(new_n949), .A3(G286), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n858), .A2(G171), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n855), .A2(new_n857), .A3(G301), .ZN(new_n952));
  AOI21_X1  g527(.A(G168), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT119), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n936), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n929), .A2(new_n931), .A3(KEYINPUT119), .A4(new_n935), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n956), .A2(new_n934), .A3(new_n957), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(G286), .B1(new_n948), .B2(new_n949), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n951), .A2(G168), .A3(new_n952), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n932), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n947), .B(new_n925), .C1(new_n959), .C2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n962), .B1(new_n954), .B2(new_n958), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n923), .A2(new_n924), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT120), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n902), .ZN(new_n968));
  INV_X1    g543(.A(new_n932), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(new_n950), .B2(new_n953), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n937), .A2(new_n961), .A3(new_n960), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n965), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT118), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT118), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n965), .A2(new_n970), .A3(new_n971), .A4(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n968), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n967), .A2(new_n976), .A3(KEYINPUT43), .ZN(new_n977));
  AOI21_X1  g552(.A(G37), .B1(new_n973), .B2(new_n975), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n970), .A2(new_n971), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT117), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n965), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(new_n980), .B2(new_n979), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT43), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT44), .B1(new_n977), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT44), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n967), .A2(new_n976), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n986), .B1(new_n978), .B2(new_n982), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n984), .A2(new_n989), .ZN(G397));
  NOR2_X1   g565(.A1(G299), .A2(KEYINPUT57), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT57), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n992), .B1(new_n930), .B2(new_n582), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G1956), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n477), .A2(new_n488), .A3(G40), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(G1384), .B1(new_n509), .B2(new_n514), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AOI211_X1 g575(.A(KEYINPUT50), .B(G1384), .C1(new_n509), .C2(new_n514), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n995), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1384), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n515), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n998), .A2(KEYINPUT45), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT56), .B(G2072), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1006), .A2(new_n1007), .A3(new_n997), .A4(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n994), .B1(new_n1002), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n994), .A2(new_n1002), .A3(new_n1009), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n794), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1004), .A2(new_n996), .ZN(new_n1013));
  INV_X1    g588(.A(G2067), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n623), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1010), .B1(new_n1011), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1002), .A2(new_n1009), .ZN(new_n1018));
  INV_X1    g593(.A(new_n994), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1020), .A2(KEYINPUT61), .A3(new_n1011), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT126), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT126), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1020), .A2(new_n1023), .A3(KEYINPUT61), .A4(new_n1011), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(KEYINPUT125), .A2(KEYINPUT59), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n564), .A2(new_n568), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n997), .B1(new_n998), .B2(KEYINPUT45), .ZN(new_n1029));
  AOI211_X1 g604(.A(new_n1005), .B(G1384), .C1(new_n509), .C2(new_n514), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n1029), .A2(G1996), .A3(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g606(.A(KEYINPUT58), .B(G1341), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1013), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1028), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(KEYINPUT125), .A2(KEYINPUT59), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1035), .B(new_n1028), .C1(new_n1031), .C2(new_n1033), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT61), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n994), .A2(new_n1002), .A3(new_n1009), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1040), .B1(new_n1041), .B2(new_n1010), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n623), .A2(KEYINPUT60), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1012), .A2(new_n1015), .A3(new_n1043), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1012), .A2(new_n1015), .A3(new_n623), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT60), .B1(new_n1045), .B2(new_n1016), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1039), .A2(new_n1042), .A3(new_n1044), .A4(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1017), .B1(new_n1025), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1006), .A2(new_n798), .A3(new_n1007), .A4(new_n997), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1004), .A2(KEYINPUT50), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n998), .A2(new_n999), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(new_n997), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1961), .ZN(new_n1055));
  AOI22_X1  g630(.A1(new_n1050), .A2(new_n1051), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1051), .A2(KEYINPUT127), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT53), .B1(new_n1051), .B2(KEYINPUT127), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1059), .A2(G171), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1055), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n1029), .A2(G2078), .A3(new_n1030), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1061), .B1(new_n1062), .B2(KEYINPUT53), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1051), .A2(new_n1050), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1063), .A2(new_n1064), .A3(G171), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1049), .B1(new_n1060), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G1966), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1068));
  INV_X1    g643(.A(G2084), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1052), .A2(new_n1069), .A3(new_n997), .A4(new_n1053), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1068), .A2(new_n1070), .A3(G168), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(G8), .ZN(new_n1072));
  AOI21_X1  g647(.A(G168), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT51), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1071), .A2(new_n1075), .A3(G8), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n997), .A2(new_n998), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT49), .ZN(new_n1079));
  OAI21_X1  g654(.A(G1981), .B1(new_n598), .B2(new_n602), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n598), .A2(new_n602), .A3(G1981), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OR3_X1    g658(.A1(new_n598), .A2(new_n602), .A3(G1981), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1084), .A2(new_n1080), .A3(KEYINPUT49), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1078), .A2(new_n1083), .A3(G8), .A4(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G1976), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT52), .B1(G288), .B2(new_n1087), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n592), .A2(new_n1087), .A3(new_n594), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1078), .A2(new_n1088), .A3(G8), .A4(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G8), .ZN(new_n1092));
  AOI211_X1 g667(.A(new_n1092), .B(new_n1089), .C1(new_n997), .C2(new_n998), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT52), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1086), .B(new_n1091), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1000), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1097), .A2(new_n788), .A3(new_n1053), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n829), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1092), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT122), .B(KEYINPUT55), .ZN(new_n1101));
  NAND3_X1  g676(.A1(G303), .A2(G8), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  AOI22_X1  g678(.A1(G303), .A2(G8), .B1(KEYINPUT122), .B2(KEYINPUT55), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1096), .B1(new_n1100), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n996), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1108));
  AOI21_X1  g683(.A(G1971), .B1(new_n1108), .B2(new_n1007), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1000), .A2(G2090), .A3(new_n1001), .ZN(new_n1110));
  OAI21_X1  g685(.A(G8), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(new_n1105), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1056), .B(G301), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1114));
  OAI21_X1  g689(.A(G171), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1114), .A2(KEYINPUT54), .A3(new_n1115), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1077), .A2(new_n1113), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1048), .A2(new_n1066), .A3(new_n1117), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1086), .A2(new_n1087), .A3(new_n821), .ZN(new_n1119));
  OAI211_X1 g694(.A(G8), .B(new_n1078), .C1(new_n1119), .C2(new_n1082), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1100), .A2(new_n1106), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1120), .B1(new_n1121), .B2(new_n1095), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1123), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1095), .B1(new_n1111), .B2(new_n1105), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1125), .A2(new_n1059), .A3(G171), .A4(new_n1121), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1074), .A2(new_n1123), .A3(new_n1076), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1122), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  AOI211_X1 g704(.A(new_n1092), .B(G286), .C1(new_n1068), .C2(new_n1070), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1125), .A2(new_n1130), .A3(new_n1121), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT63), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1131), .A2(KEYINPUT123), .A3(new_n1132), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1105), .A2(KEYINPUT124), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n1111), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1095), .A2(new_n1132), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1111), .A2(new_n1137), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1138), .A2(new_n1130), .A3(new_n1139), .A4(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1135), .A2(new_n1136), .A3(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1118), .A2(new_n1129), .A3(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1006), .A2(new_n996), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n729), .A2(G2067), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n723), .A2(new_n728), .A3(new_n1014), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT121), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n746), .B(G1996), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1149), .B1(new_n1144), .B2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n813), .A2(new_n816), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n813), .A2(new_n816), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1144), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(G290), .B(G1986), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1155), .B1(new_n1144), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1143), .A2(new_n1157), .ZN(new_n1158));
  OR3_X1    g733(.A1(new_n1006), .A2(G1996), .A3(new_n996), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT46), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1145), .A2(new_n888), .A3(new_n1146), .ZN(new_n1161));
  AOI22_X1  g736(.A1(new_n1159), .A2(new_n1160), .B1(new_n1144), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1162), .B1(new_n1160), .B2(new_n1159), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1163), .B(KEYINPUT47), .ZN(new_n1164));
  NOR4_X1   g739(.A1(new_n1006), .A2(G1986), .A3(G290), .A4(new_n996), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1165), .B(KEYINPUT48), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1164), .B1(new_n1155), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n1146), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1167), .B1(new_n1144), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1158), .A2(new_n1170), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g746(.A1(G227), .A2(new_n463), .ZN(new_n1173));
  AOI21_X1  g747(.A(new_n1173), .B1(new_n665), .B2(new_n667), .ZN(new_n1174));
  NAND3_X1  g748(.A1(new_n909), .A2(new_n711), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g749(.A1(new_n978), .A2(new_n982), .ZN(new_n1176));
  NAND2_X1  g750(.A1(new_n1176), .A2(KEYINPUT43), .ZN(new_n1177));
  NAND3_X1  g751(.A1(new_n967), .A2(new_n976), .A3(new_n986), .ZN(new_n1178));
  AOI21_X1  g752(.A(new_n1175), .B1(new_n1177), .B2(new_n1178), .ZN(G308));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1180));
  NAND4_X1  g754(.A1(new_n1180), .A2(new_n711), .A3(new_n909), .A4(new_n1174), .ZN(G225));
endmodule


