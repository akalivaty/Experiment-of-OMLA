//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n795, new_n797, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929;
  NOR2_X1   g000(.A1(G29gat), .A2(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT14), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT96), .B(G36gat), .ZN(new_n204));
  AOI21_X1  g003(.A(new_n203), .B1(G29gat), .B2(new_n204), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n205), .A2(KEYINPUT15), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(KEYINPUT15), .ZN(new_n207));
  XNOR2_X1  g006(.A(G43gat), .B(G50gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n207), .A2(new_n208), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT97), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT17), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G15gat), .B(G22gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT16), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(G1gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G1gat), .B2(new_n215), .ZN(new_n218));
  INV_X1    g017(.A(G8gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G229gat), .A2(G233gat), .ZN(new_n222));
  INV_X1    g021(.A(new_n220), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n211), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n221), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT18), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G113gat), .B(G141gat), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n228), .B(G197gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT11), .B(G169gat), .ZN(new_n230));
  XOR2_X1   g029(.A(new_n229), .B(new_n230), .Z(new_n231));
  XOR2_X1   g030(.A(new_n231), .B(KEYINPUT12), .Z(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n221), .A2(KEYINPUT18), .A3(new_n222), .A4(new_n224), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n211), .B(new_n223), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n222), .B(KEYINPUT13), .Z(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n227), .A2(new_n233), .A3(new_n234), .A4(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT98), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n225), .A2(new_n226), .B1(new_n235), .B2(new_n236), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT98), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n240), .A2(new_n241), .A3(new_n233), .A4(new_n234), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n234), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n239), .A2(new_n242), .B1(new_n243), .B2(new_n232), .ZN(new_n244));
  NAND2_X1  g043(.A1(G85gat), .A2(G92gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT7), .ZN(new_n246));
  NAND2_X1  g045(.A1(G99gat), .A2(G106gat), .ZN(new_n247));
  INV_X1    g046(.A(G85gat), .ZN(new_n248));
  INV_X1    g047(.A(G92gat), .ZN(new_n249));
  AOI22_X1  g048(.A1(KEYINPUT8), .A2(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G99gat), .B(G106gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n253), .B(KEYINPUT101), .Z(new_n254));
  NAND2_X1  g053(.A1(new_n214), .A2(new_n254), .ZN(new_n255));
  AND2_X1   g054(.A1(G232gat), .A2(G233gat), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n211), .A2(new_n253), .B1(KEYINPUT41), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G190gat), .B(G218gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT102), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n256), .A2(KEYINPUT41), .ZN(new_n262));
  XOR2_X1   g061(.A(new_n262), .B(KEYINPUT100), .Z(new_n263));
  XNOR2_X1  g062(.A(G134gat), .B(G162gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n260), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n255), .A2(new_n266), .A3(new_n257), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n261), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n265), .B1(new_n261), .B2(new_n267), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(G71gat), .B(G78gat), .Z(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT9), .ZN(new_n274));
  INV_X1    g073(.A(G71gat), .ZN(new_n275));
  INV_X1    g074(.A(G78gat), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(G57gat), .B(G64gat), .Z(new_n278));
  NAND3_X1  g077(.A1(new_n273), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n277), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(new_n272), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT21), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(G231gat), .A2(G233gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G127gat), .B(G155gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(KEYINPUT20), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n286), .B(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G183gat), .B(G211gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n220), .B1(new_n283), .B2(new_n282), .ZN(new_n292));
  XOR2_X1   g091(.A(KEYINPUT99), .B(KEYINPUT19), .Z(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n291), .B(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n271), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n252), .A2(KEYINPUT103), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n282), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n298), .B(new_n253), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n253), .A2(KEYINPUT10), .A3(new_n281), .A4(new_n279), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G230gat), .A2(G233gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n299), .A2(G230gat), .A3(G233gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(G120gat), .B(G148gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(G176gat), .B(G204gat), .ZN(new_n307));
  XOR2_X1   g106(.A(new_n306), .B(new_n307), .Z(new_n308));
  NAND3_X1  g107(.A1(new_n304), .A2(new_n305), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  XOR2_X1   g109(.A(new_n303), .B(KEYINPUT104), .Z(new_n311));
  AOI21_X1  g110(.A(new_n311), .B1(new_n300), .B2(new_n301), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n308), .B1(new_n313), .B2(new_n305), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n296), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G15gat), .B(G43gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(KEYINPUT77), .ZN(new_n318));
  XNOR2_X1  g117(.A(G71gat), .B(G99gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n319), .B(KEYINPUT78), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n318), .B(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT25), .ZN(new_n322));
  INV_X1    g121(.A(G169gat), .ZN(new_n323));
  INV_X1    g122(.A(G176gat), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT23), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT23), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n326), .B1(G169gat), .B2(G176gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(G169gat), .A2(G176gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT67), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G183gat), .A2(G190gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT24), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT24), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(G183gat), .A3(G190gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  AOI211_X1 g136(.A(new_n322), .B(new_n329), .C1(new_n332), .C2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n339));
  AND3_X1   g138(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n330), .B1(new_n334), .B2(new_n336), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT65), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AOI211_X1 g142(.A(KEYINPUT65), .B(new_n330), .C1(new_n334), .C2(new_n336), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n339), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT66), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n338), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI211_X1 g146(.A(KEYINPUT66), .B(new_n339), .C1(new_n343), .C2(new_n344), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n349));
  NOR4_X1   g148(.A1(KEYINPUT70), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT70), .ZN(new_n351));
  NOR2_X1   g150(.A1(G169gat), .A2(G176gat), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT26), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n328), .B(new_n349), .C1(new_n350), .C2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT71), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n355), .A2(new_n356), .A3(new_n333), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n356), .B1(new_n355), .B2(new_n333), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT28), .ZN(new_n360));
  XNOR2_X1  g159(.A(KEYINPUT27), .B(G183gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(KEYINPUT68), .ZN(new_n362));
  INV_X1    g161(.A(G190gat), .ZN(new_n363));
  INV_X1    g162(.A(G183gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n364), .A2(KEYINPUT27), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT68), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n363), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n360), .B1(new_n362), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT69), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI211_X1 g169(.A(KEYINPUT69), .B(new_n360), .C1(new_n362), .C2(new_n367), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n361), .A2(KEYINPUT28), .A3(new_n363), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n347), .A2(new_n348), .B1(new_n359), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(G127gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(G134gat), .ZN(new_n376));
  INV_X1    g175(.A(G134gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G127gat), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT1), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT75), .ZN(new_n381));
  INV_X1    g180(.A(G120gat), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n381), .B1(new_n382), .B2(G113gat), .ZN(new_n383));
  INV_X1    g182(.A(G113gat), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n384), .A2(KEYINPUT75), .A3(G120gat), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT74), .B(G120gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(G113gat), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n380), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n384), .A2(G120gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n382), .A2(G113gat), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT1), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OR2_X1    g191(.A1(KEYINPUT72), .A2(G134gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(KEYINPUT72), .A2(G134gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(G127gat), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n376), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n392), .B1(new_n396), .B2(KEYINPUT73), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT73), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n395), .A2(new_n398), .A3(new_n376), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n389), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n374), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT76), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n374), .A2(KEYINPUT76), .A3(new_n400), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n345), .A2(new_n346), .ZN(new_n405));
  INV_X1    g204(.A(new_n338), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(new_n348), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n359), .A2(new_n373), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AND2_X1   g208(.A1(KEYINPUT72), .A2(G134gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(KEYINPUT72), .A2(G134gat), .ZN(new_n411));
  NOR3_X1   g210(.A1(new_n410), .A2(new_n411), .A3(new_n375), .ZN(new_n412));
  INV_X1    g211(.A(new_n376), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT73), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n392), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n399), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n386), .A2(new_n388), .ZN(new_n417));
  INV_X1    g216(.A(new_n380), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n409), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n403), .A2(new_n404), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(G227gat), .A2(G233gat), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT33), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n321), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n403), .A2(new_n423), .A3(new_n404), .A4(new_n421), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT34), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n374), .A2(new_n400), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n430), .B1(new_n402), .B2(new_n401), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT34), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n431), .A2(new_n432), .A3(new_n423), .A4(new_n404), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n427), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT33), .B1(new_n422), .B2(new_n424), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n429), .B(new_n433), .C1(new_n436), .C2(new_n321), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n425), .A2(KEYINPUT32), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n439), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n435), .A2(new_n441), .A3(new_n437), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT36), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n440), .A2(KEYINPUT36), .A3(new_n442), .ZN(new_n446));
  XNOR2_X1  g245(.A(G78gat), .B(G106gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(KEYINPUT31), .B(G50gat), .ZN(new_n448));
  XOR2_X1   g247(.A(new_n447), .B(new_n448), .Z(new_n449));
  XNOR2_X1  g248(.A(G197gat), .B(G204gat), .ZN(new_n450));
  INV_X1    g249(.A(G211gat), .ZN(new_n451));
  INV_X1    g250(.A(G218gat), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n450), .B1(KEYINPUT22), .B2(new_n453), .ZN(new_n454));
  XOR2_X1   g253(.A(G211gat), .B(G218gat), .Z(new_n455));
  XNOR2_X1  g254(.A(new_n454), .B(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT29), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT3), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OR2_X1    g257(.A1(KEYINPUT82), .A2(G148gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(KEYINPUT82), .A2(G148gat), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(G141gat), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(G148gat), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT81), .B1(new_n462), .B2(G141gat), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT81), .ZN(new_n464));
  INV_X1    g263(.A(G141gat), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(new_n465), .A3(G148gat), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n461), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(G155gat), .A2(G162gat), .ZN(new_n468));
  NOR2_X1   g267(.A1(G155gat), .A2(G162gat), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n468), .B1(new_n470), .B2(KEYINPUT2), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT2), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n462), .A2(G141gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n465), .A2(G148gat), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AND2_X1   g274(.A1(G155gat), .A2(G162gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n476), .A2(new_n469), .ZN(new_n477));
  AOI22_X1  g276(.A1(new_n467), .A2(new_n471), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  OR2_X1    g277(.A1(new_n458), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(new_n457), .ZN(new_n482));
  INV_X1    g281(.A(new_n456), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n479), .A2(new_n484), .B1(G228gat), .B2(G233gat), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT83), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n476), .B1(new_n472), .B2(new_n469), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n463), .A2(new_n466), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n487), .B1(new_n488), .B2(new_n461), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n470), .A2(new_n468), .ZN(new_n490));
  XOR2_X1   g289(.A(G141gat), .B(G148gat), .Z(new_n491));
  AOI21_X1  g290(.A(new_n490), .B1(new_n491), .B2(new_n472), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n486), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n459), .A2(G141gat), .A3(new_n460), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n463), .A2(new_n466), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n471), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n475), .A2(new_n477), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(KEYINPUT83), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  OR3_X1    g298(.A1(new_n458), .A2(new_n499), .A3(KEYINPUT89), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT89), .B1(new_n458), .B2(new_n499), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n484), .A2(G228gat), .A3(G233gat), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n485), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  XOR2_X1   g303(.A(KEYINPUT90), .B(G22gat), .Z(new_n505));
  AOI21_X1  g304(.A(new_n449), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n502), .A2(new_n503), .ZN(new_n507));
  OAI21_X1  g306(.A(G22gat), .B1(new_n507), .B2(new_n485), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT91), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n506), .A2(new_n508), .A3(KEYINPUT91), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n504), .B(new_n505), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n449), .ZN(new_n514));
  XOR2_X1   g313(.A(G1gat), .B(G29gat), .Z(new_n515));
  XNOR2_X1  g314(.A(G57gat), .B(G85gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT87), .B(KEYINPUT0), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT4), .B1(new_n400), .B2(new_n478), .ZN(new_n520));
  AND4_X1   g319(.A1(KEYINPUT4), .A2(new_n416), .A3(new_n419), .A4(new_n478), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n420), .A2(KEYINPUT84), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n493), .A2(KEYINPUT3), .A3(new_n498), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT84), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n416), .A2(new_n419), .A3(new_n525), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n523), .A2(new_n524), .A3(new_n526), .A4(new_n481), .ZN(new_n527));
  NAND2_X1  g326(.A1(G225gat), .A2(G233gat), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n528), .B(KEYINPUT85), .Z(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n522), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT5), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n532), .A2(KEYINPUT86), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n533), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n522), .A2(new_n527), .A3(new_n530), .A4(new_n535), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n523), .A2(new_n526), .A3(new_n493), .A4(new_n498), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n416), .A2(new_n478), .A3(new_n419), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n530), .A2(new_n532), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g341(.A(KEYINPUT88), .B(new_n519), .C1(new_n537), .C2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT88), .ZN(new_n544));
  AOI22_X1  g343(.A1(new_n534), .A2(new_n536), .B1(new_n540), .B2(new_n541), .ZN(new_n545));
  INV_X1    g344(.A(new_n519), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT6), .B1(new_n545), .B2(new_n546), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n543), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n545), .A2(KEYINPUT6), .A3(new_n546), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(G226gat), .A2(G233gat), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n552), .B(KEYINPUT79), .Z(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n554), .B1(new_n409), .B2(new_n457), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n374), .A2(new_n553), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n483), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G8gat), .B(G36gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT80), .ZN(new_n559));
  XNOR2_X1  g358(.A(G64gat), .B(G92gat), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n559), .B(new_n560), .Z(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n553), .B1(new_n374), .B2(KEYINPUT29), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n409), .A2(new_n554), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n456), .A3(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n557), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT30), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR3_X1   g367(.A1(new_n555), .A2(new_n556), .A3(new_n483), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n456), .B1(new_n563), .B2(new_n564), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n561), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n557), .A2(KEYINPUT30), .A3(new_n565), .A4(new_n562), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n551), .A2(new_n574), .ZN(new_n575));
  AOI22_X1  g374(.A1(new_n445), .A2(new_n446), .B1(new_n514), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT94), .ZN(new_n577));
  AND4_X1   g376(.A1(new_n523), .A2(new_n524), .A3(new_n526), .A4(new_n481), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT4), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n539), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n400), .A2(KEYINPUT4), .A3(new_n478), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n529), .B1(new_n578), .B2(new_n582), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n583), .B(KEYINPUT39), .C1(new_n529), .C2(new_n540), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT92), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n530), .B1(new_n522), .B2(new_n527), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT39), .ZN(new_n587));
  AOI211_X1 g386(.A(new_n585), .B(new_n546), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n587), .B(new_n529), .C1(new_n578), .C2(new_n582), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT92), .B1(new_n589), .B2(new_n519), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n584), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT93), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT40), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT93), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n594), .B(new_n584), .C1(new_n588), .C2(new_n590), .ZN(new_n595));
  AND3_X1   g394(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n545), .A2(new_n546), .ZN(new_n597));
  OAI211_X1 g396(.A(KEYINPUT40), .B(new_n584), .C1(new_n588), .C2(new_n590), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n597), .B(new_n598), .C1(new_n568), .C2(new_n573), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n577), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(new_n597), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n566), .A2(new_n567), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n604), .A2(new_n572), .A3(new_n571), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n601), .A2(new_n603), .A3(KEYINPUT94), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n600), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT37), .B1(new_n569), .B2(new_n570), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT37), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n557), .A2(new_n609), .A3(new_n565), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n561), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT38), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT38), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n608), .A2(new_n613), .A3(new_n561), .A4(new_n610), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n550), .A2(new_n566), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n612), .A2(new_n549), .A3(new_n614), .A4(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n513), .A2(new_n449), .ZN(new_n617));
  INV_X1    g416(.A(new_n512), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT91), .B1(new_n506), .B2(new_n508), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n607), .A2(KEYINPUT95), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT95), .B1(new_n607), .B2(new_n621), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n576), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n442), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n441), .B1(new_n435), .B2(new_n437), .ZN(new_n626));
  NOR3_X1   g425(.A1(new_n625), .A2(new_n514), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT35), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n627), .A2(new_n628), .A3(new_n574), .A4(new_n551), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n440), .A2(new_n574), .A3(new_n620), .A4(new_n442), .ZN(new_n630));
  INV_X1    g429(.A(new_n551), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT35), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  AOI211_X1 g432(.A(new_n244), .B(new_n316), .C1(new_n624), .C2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n551), .B(KEYINPUT105), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(KEYINPUT106), .B(G1gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(G1324gat));
  XOR2_X1   g438(.A(KEYINPUT16), .B(G8gat), .Z(new_n640));
  NAND4_X1  g439(.A1(new_n634), .A2(KEYINPUT42), .A3(new_n605), .A4(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n634), .A2(new_n605), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT108), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n643), .A2(new_n640), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n645));
  OAI221_X1 g444(.A(new_n641), .B1(new_n219), .B2(new_n643), .C1(new_n644), .C2(new_n645), .ZN(G1325gat));
  INV_X1    g445(.A(G15gat), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n634), .A2(new_n647), .A3(new_n442), .A4(new_n440), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n625), .A2(new_n444), .A3(new_n626), .ZN(new_n649));
  AOI21_X1  g448(.A(KEYINPUT36), .B1(new_n440), .B2(new_n442), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n634), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n648), .B1(new_n652), .B2(new_n647), .ZN(G1326gat));
  NAND2_X1  g452(.A1(new_n634), .A2(new_n514), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT109), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT43), .B(G22gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(G1327gat));
  NAND2_X1  g456(.A1(new_n575), .A2(new_n514), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n658), .B1(new_n649), .B2(new_n650), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n574), .A2(new_n602), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT94), .B1(new_n660), .B2(new_n601), .ZN(new_n661));
  AND4_X1   g460(.A1(KEYINPUT94), .A2(new_n601), .A3(new_n605), .A4(new_n603), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n621), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT95), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n607), .A2(KEYINPUT95), .A3(new_n621), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n659), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n633), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n271), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n624), .A2(new_n633), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n672), .A2(KEYINPUT44), .A3(new_n271), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n295), .ZN(new_n675));
  INV_X1    g474(.A(new_n315), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n244), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(G29gat), .B1(new_n678), .B2(new_n635), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n672), .A2(new_n271), .A3(new_n677), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n680), .A2(G29gat), .A3(new_n635), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT110), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n683), .A2(KEYINPUT45), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(KEYINPUT45), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n679), .B1(new_n684), .B2(new_n685), .ZN(G1328gat));
  OAI21_X1  g485(.A(new_n204), .B1(new_n678), .B2(new_n574), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n680), .A2(new_n574), .A3(new_n204), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT111), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n690), .A2(KEYINPUT46), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(KEYINPUT46), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n687), .B1(new_n691), .B2(new_n692), .ZN(G1329gat));
  NAND2_X1  g492(.A1(new_n651), .A2(G43gat), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n680), .A2(new_n443), .ZN(new_n695));
  OAI22_X1  g494(.A1(new_n678), .A2(new_n694), .B1(G43gat), .B2(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g496(.A(KEYINPUT48), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(KEYINPUT112), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n620), .A2(G50gat), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n699), .B1(new_n680), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n674), .A2(new_n514), .A3(new_n677), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n702), .B1(new_n703), .B2(G50gat), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n698), .A2(KEYINPUT112), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1331gat));
  AND4_X1   g505(.A1(new_n672), .A2(new_n244), .A3(new_n296), .A4(new_n676), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n636), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n605), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n710), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT49), .B(G64gat), .Z(new_n712));
  OAI21_X1  g511(.A(new_n711), .B1(new_n710), .B2(new_n712), .ZN(G1333gat));
  AOI21_X1  g512(.A(new_n275), .B1(new_n707), .B2(new_n651), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n443), .A2(G71gat), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n714), .B1(new_n707), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g516(.A1(new_n707), .A2(new_n514), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g518(.A1(new_n239), .A2(new_n242), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n243), .A2(new_n232), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(new_n675), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n676), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT113), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n674), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(G85gat), .B1(new_n726), .B2(new_n635), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n271), .B(new_n723), .C1(new_n667), .C2(new_n668), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT51), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n672), .A2(KEYINPUT51), .A3(new_n271), .A4(new_n723), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n636), .A2(new_n248), .A3(new_n676), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n727), .B1(new_n733), .B2(new_n734), .ZN(G1336gat));
  OAI21_X1  g534(.A(G92gat), .B1(new_n726), .B2(new_n574), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n732), .A2(new_n249), .A3(new_n605), .A4(new_n676), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(KEYINPUT52), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n736), .A2(new_n740), .A3(new_n737), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n741), .ZN(G1337gat));
  INV_X1    g541(.A(new_n651), .ZN(new_n743));
  OAI21_X1  g542(.A(G99gat), .B1(new_n726), .B2(new_n743), .ZN(new_n744));
  OR3_X1    g543(.A1(new_n443), .A2(G99gat), .A3(new_n315), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n733), .B2(new_n745), .ZN(G1338gat));
  NAND4_X1  g545(.A1(new_n671), .A2(new_n514), .A3(new_n673), .A4(new_n725), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G106gat), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT115), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n620), .A2(G106gat), .A3(new_n315), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n732), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n748), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT114), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT53), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  AOI22_X1  g554(.A1(G106gat), .A2(new_n747), .B1(new_n732), .B2(new_n750), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT114), .B1(new_n756), .B2(new_n749), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n748), .A2(KEYINPUT114), .A3(new_n751), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT53), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n755), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(G1339gat));
  INV_X1    g560(.A(new_n311), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n304), .B(KEYINPUT54), .C1(new_n762), .C2(new_n302), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT54), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n308), .B1(new_n312), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n763), .A2(KEYINPUT55), .A3(new_n765), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n768), .A2(new_n309), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n720), .B2(new_n721), .ZN(new_n771));
  INV_X1    g570(.A(new_n231), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n221), .A2(new_n224), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n773), .A2(G229gat), .A3(G233gat), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n235), .A2(new_n236), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n772), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  AOI211_X1 g576(.A(new_n315), .B(new_n777), .C1(new_n239), .C2(new_n242), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n270), .B1(new_n771), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n270), .A2(new_n770), .ZN(new_n780));
  INV_X1    g579(.A(new_n777), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n780), .A2(new_n720), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n295), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n316), .A2(new_n722), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n635), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n630), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(new_n244), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(new_n384), .ZN(G1340gat));
  OAI21_X1  g590(.A(G120gat), .B1(new_n789), .B2(new_n315), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n676), .A2(new_n387), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT116), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n792), .B1(new_n789), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT117), .ZN(G1341gat));
  NOR2_X1   g595(.A1(new_n789), .A2(new_n295), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(new_n375), .ZN(G1342gat));
  NAND3_X1  g597(.A1(new_n787), .A2(new_n788), .A3(new_n271), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n393), .A2(new_n394), .ZN(new_n800));
  OR3_X1    g599(.A1(new_n799), .A2(KEYINPUT56), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT56), .B1(new_n799), .B2(new_n800), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT118), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n799), .A2(new_n803), .A3(G134gat), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n803), .B1(new_n799), .B2(G134gat), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n801), .B(new_n802), .C1(new_n805), .C2(new_n806), .ZN(G1343gat));
  OAI21_X1  g606(.A(KEYINPUT121), .B1(new_n651), .B2(new_n620), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n651), .A2(new_n620), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT121), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n605), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n244), .A2(G141gat), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n787), .A2(new_n808), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT120), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n675), .B1(new_n779), .B2(new_n782), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n514), .B1(new_n816), .B2(new_n785), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n780), .A2(new_n720), .A3(new_n781), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n720), .A2(new_n676), .A3(new_n781), .ZN(new_n820));
  XNOR2_X1  g619(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n766), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n822), .A2(new_n309), .A3(new_n769), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n820), .B1(new_n244), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n819), .B1(new_n824), .B2(new_n270), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n786), .B1(new_n825), .B2(new_n675), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n620), .A2(new_n818), .ZN(new_n827));
  AOI22_X1  g626(.A1(new_n817), .A2(new_n818), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n635), .A2(new_n605), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n743), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n815), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n830), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n820), .B1(new_n244), .B2(new_n770), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n819), .B1(new_n833), .B2(new_n270), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n786), .B1(new_n834), .B2(new_n675), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT57), .B1(new_n835), .B2(new_n514), .ZN(new_n836));
  INV_X1    g635(.A(new_n827), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n244), .A2(new_n823), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n271), .B1(new_n838), .B2(new_n820), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n295), .B1(new_n839), .B2(new_n819), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n837), .B1(new_n840), .B2(new_n786), .ZN(new_n841));
  OAI211_X1 g640(.A(KEYINPUT120), .B(new_n832), .C1(new_n836), .C2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n831), .A2(new_n722), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n814), .B1(new_n843), .B2(G141gat), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n722), .B(new_n832), .C1(new_n836), .C2(new_n841), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(G141gat), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n813), .A2(new_n845), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n847), .A2(KEYINPUT122), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT122), .B1(new_n847), .B2(new_n848), .ZN(new_n850));
  OAI22_X1  g649(.A1(new_n844), .A2(new_n845), .B1(new_n849), .B2(new_n850), .ZN(G1344gat));
  NAND2_X1  g650(.A1(new_n826), .A2(new_n514), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n818), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n835), .A2(new_n827), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n676), .A3(new_n832), .ZN(new_n856));
  AND2_X1   g655(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n787), .A2(new_n808), .A3(new_n811), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n459), .A2(new_n460), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n315), .A2(new_n859), .ZN(new_n860));
  AOI22_X1  g659(.A1(new_n856), .A2(new_n857), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n831), .A2(new_n676), .A3(new_n842), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n862), .A2(new_n859), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n861), .B1(new_n863), .B2(KEYINPUT59), .ZN(G1345gat));
  INV_X1    g663(.A(G155gat), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n295), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n831), .A2(new_n842), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n858), .A2(new_n675), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n865), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n867), .A2(new_n869), .A3(KEYINPUT123), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(G1346gat));
  AOI21_X1  g673(.A(G162gat), .B1(new_n858), .B2(new_n271), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n831), .A2(new_n842), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n271), .A2(G162gat), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(G1347gat));
  AOI21_X1  g677(.A(new_n636), .B1(new_n784), .B2(new_n786), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n443), .A2(new_n574), .A3(new_n514), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(new_n244), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(new_n323), .ZN(G1348gat));
  INV_X1    g682(.A(KEYINPUT124), .ZN(new_n884));
  INV_X1    g683(.A(new_n881), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n676), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n884), .B1(new_n886), .B2(new_n324), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n885), .A2(KEYINPUT124), .A3(G176gat), .A4(new_n676), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n324), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(G1349gat));
  OAI21_X1  g689(.A(new_n364), .B1(new_n881), .B2(new_n295), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n885), .A2(new_n675), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n892), .B2(new_n361), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT60), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n893), .B(new_n894), .ZN(G1350gat));
  NOR2_X1   g694(.A1(new_n881), .A2(new_n270), .ZN(new_n896));
  NAND2_X1  g695(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  XOR2_X1   g697(.A(KEYINPUT61), .B(G190gat), .Z(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n896), .B2(new_n899), .ZN(G1351gat));
  AND3_X1   g699(.A1(new_n879), .A2(new_n605), .A3(new_n809), .ZN(new_n901));
  AOI21_X1  g700(.A(G197gat), .B1(new_n901), .B2(new_n722), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n651), .A2(new_n574), .A3(new_n636), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n904), .B1(new_n853), .B2(new_n854), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n722), .A2(G197gat), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(G1352gat));
  AOI21_X1  g706(.A(G204gat), .B1(KEYINPUT125), .B2(KEYINPUT62), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n901), .A2(new_n676), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n909), .B(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n905), .A2(new_n676), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(G204gat), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n912), .A2(new_n913), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n911), .B1(new_n915), .B2(new_n916), .ZN(G1353gat));
  NAND3_X1  g716(.A1(new_n901), .A2(new_n451), .A3(new_n675), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n905), .A2(new_n675), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n919), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n920));
  AOI21_X1  g719(.A(KEYINPUT63), .B1(new_n919), .B2(G211gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(G1354gat));
  INV_X1    g721(.A(KEYINPUT127), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n901), .A2(new_n452), .A3(new_n271), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n905), .A2(new_n271), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n923), .B(new_n924), .C1(new_n925), .C2(new_n452), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n452), .B1(new_n905), .B2(new_n271), .ZN(new_n927));
  INV_X1    g726(.A(new_n924), .ZN(new_n928));
  OAI21_X1  g727(.A(KEYINPUT127), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n926), .A2(new_n929), .ZN(G1355gat));
endmodule


