//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n817, new_n818, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012;
  INV_X1    g000(.A(KEYINPUT95), .ZN(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  INV_X1    g002(.A(G36gat), .ZN(new_n204));
  NAND4_X1  g003(.A1(new_n202), .A2(new_n203), .A3(new_n204), .A4(KEYINPUT14), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT14), .ZN(new_n206));
  OAI22_X1  g005(.A1(new_n206), .A2(KEYINPUT95), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n202), .A2(KEYINPUT14), .ZN(new_n208));
  OAI221_X1 g007(.A(new_n205), .B1(new_n203), .B2(new_n204), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT15), .ZN(new_n210));
  XOR2_X1   g009(.A(G43gat), .B(G50gat), .Z(new_n211));
  AOI21_X1  g010(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n211), .A2(new_n210), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n213), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G15gat), .B(G22gat), .ZN(new_n217));
  INV_X1    g016(.A(G1gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT16), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(G1gat), .B2(new_n217), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n221), .A2(G8gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(G8gat), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n216), .B(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G229gat), .A2(G233gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n227), .B(KEYINPUT13), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT17), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n216), .A2(new_n231), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n224), .A2(KEYINPUT96), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n214), .A2(KEYINPUT17), .A3(new_n215), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n224), .A2(KEYINPUT96), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n232), .A2(new_n233), .A3(new_n234), .A4(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n216), .A2(new_n225), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(new_n227), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT18), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n230), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n239), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n240), .B1(new_n242), .B2(KEYINPUT98), .ZN(new_n243));
  XNOR2_X1  g042(.A(G113gat), .B(G141gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT93), .B(KEYINPUT11), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G169gat), .B(G197gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n248), .B(KEYINPUT12), .Z(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT98), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n250), .B1(new_n241), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n243), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n241), .A2(KEYINPUT97), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT97), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n255), .B1(new_n238), .B2(new_n239), .ZN(new_n256));
  NOR3_X1   g055(.A1(new_n254), .A2(new_n240), .A3(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n249), .B(KEYINPUT94), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n253), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT101), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT7), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(KEYINPUT101), .A2(KEYINPUT7), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n262), .A2(G85gat), .A3(G92gat), .A4(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(KEYINPUT101), .A2(KEYINPUT7), .ZN(new_n265));
  NAND2_X1  g064(.A1(G85gat), .A2(G92gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(G99gat), .A2(G106gat), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n265), .A2(new_n266), .B1(new_n267), .B2(KEYINPUT8), .ZN(new_n268));
  OR2_X1    g067(.A1(G85gat), .A2(G92gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n264), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G99gat), .B(G106gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  OR3_X1    g071(.A1(new_n270), .A2(KEYINPUT102), .A3(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT102), .B1(new_n270), .B2(new_n272), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G57gat), .B(G64gat), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n277));
  OR2_X1    g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G71gat), .B(G78gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n270), .B(KEYINPUT106), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n275), .B(new_n280), .C1(new_n271), .C2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT103), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n275), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n273), .A2(KEYINPUT103), .A3(new_n274), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n284), .A2(new_n285), .B1(new_n272), .B2(new_n270), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n282), .B1(new_n286), .B2(new_n280), .ZN(new_n287));
  OR2_X1    g086(.A1(new_n287), .A2(KEYINPUT10), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n286), .A2(KEYINPUT104), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n270), .A2(new_n272), .ZN(new_n290));
  INV_X1    g089(.A(new_n285), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT103), .B1(new_n273), .B2(new_n274), .ZN(new_n292));
  OAI211_X1 g091(.A(KEYINPUT104), .B(new_n290), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  OAI211_X1 g093(.A(KEYINPUT10), .B(new_n280), .C1(new_n289), .C2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n288), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G230gat), .A2(G233gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n297), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n287), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G120gat), .B(G148gat), .ZN(new_n302));
  INV_X1    g101(.A(G176gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G204gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n306), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n298), .A2(new_n300), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n280), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT21), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n314));
  XOR2_X1   g113(.A(new_n313), .B(new_n314), .Z(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n224), .B1(new_n312), .B2(new_n311), .ZN(new_n317));
  INV_X1    g116(.A(G183gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT99), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n320), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n322), .A2(new_n323), .A3(G231gat), .A4(G233gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n317), .B(G183gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n325), .A2(KEYINPUT99), .ZN(new_n326));
  INV_X1    g125(.A(G231gat), .ZN(new_n327));
  INV_X1    g126(.A(G233gat), .ZN(new_n328));
  OAI22_X1  g127(.A1(new_n321), .A2(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G127gat), .B(G155gat), .ZN(new_n330));
  INV_X1    g129(.A(G211gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n324), .A2(new_n329), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n333), .B1(new_n324), .B2(new_n329), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n316), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n336), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n338), .A2(new_n315), .A3(new_n334), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT105), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n341), .B1(new_n289), .B2(new_n294), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n232), .A2(new_n234), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT104), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n346), .A2(KEYINPUT105), .A3(new_n293), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n342), .A2(new_n343), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n216), .B1(new_n289), .B2(new_n294), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G190gat), .ZN(new_n352));
  INV_X1    g151(.A(G190gat), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n348), .A2(new_n353), .A3(new_n349), .A4(new_n350), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(G218gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n352), .A2(G218gat), .A3(new_n354), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(KEYINPUT100), .A3(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G134gat), .B(G162gat), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n357), .A2(KEYINPUT100), .A3(new_n358), .A4(new_n362), .ZN(new_n365));
  AOI211_X1 g164(.A(new_n310), .B(new_n340), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G227gat), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n367), .A2(new_n328), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT1), .ZN(new_n370));
  XNOR2_X1  g169(.A(G127gat), .B(G134gat), .ZN(new_n371));
  XOR2_X1   g170(.A(KEYINPUT71), .B(G113gat), .Z(new_n372));
  INV_X1    g171(.A(G120gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT70), .B(G120gat), .ZN(new_n375));
  INV_X1    g174(.A(G113gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n370), .B(new_n371), .C1(new_n374), .C2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n370), .B1(new_n376), .B2(new_n373), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n379), .B1(new_n376), .B2(new_n373), .ZN(new_n380));
  OR2_X1    g179(.A1(new_n380), .A2(new_n371), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT23), .ZN(new_n383));
  INV_X1    g182(.A(G169gat), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n384), .A3(new_n303), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G169gat), .A2(G176gat), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT64), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n387), .A2(new_n392), .A3(KEYINPUT65), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT65), .B1(new_n387), .B2(new_n392), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n318), .A2(new_n353), .ZN(new_n396));
  NAND2_X1  g195(.A1(G183gat), .A2(G190gat), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(KEYINPUT24), .A3(new_n397), .ZN(new_n398));
  OR2_X1    g197(.A1(new_n397), .A2(KEYINPUT24), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT25), .B1(new_n395), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT66), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n403), .A2(new_n384), .A3(new_n303), .A4(KEYINPUT23), .ZN(new_n404));
  OAI22_X1  g203(.A1(new_n383), .A2(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n405), .A3(KEYINPUT25), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n390), .A2(new_n391), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n400), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(KEYINPUT67), .B1(new_n402), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n387), .A2(new_n392), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT65), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n387), .A2(new_n392), .A3(KEYINPUT65), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n412), .A2(new_n401), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT25), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n408), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT67), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n409), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT27), .B(G183gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n353), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(KEYINPUT28), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT68), .ZN(new_n424));
  NOR2_X1   g223(.A1(G169gat), .A2(G176gat), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n424), .B1(new_n425), .B2(KEYINPUT66), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT26), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n403), .B1(new_n427), .B2(KEYINPUT68), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n429), .A2(new_n425), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n392), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT69), .B1(new_n431), .B2(new_n397), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n426), .A2(new_n427), .B1(new_n425), .B2(new_n429), .ZN(new_n433));
  OAI211_X1 g232(.A(KEYINPUT69), .B(new_n397), .C1(new_n433), .C2(new_n407), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n423), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n382), .B1(new_n419), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n414), .A2(new_n415), .ZN(new_n438));
  INV_X1    g237(.A(new_n408), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n417), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AOI211_X1 g239(.A(KEYINPUT67), .B(new_n408), .C1(new_n414), .C2(new_n415), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n382), .B(new_n436), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n369), .B1(new_n437), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT34), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI211_X1 g245(.A(KEYINPUT34), .B(new_n369), .C1(new_n437), .C2(new_n443), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n436), .B1(new_n440), .B2(new_n441), .ZN(new_n449));
  INV_X1    g248(.A(new_n382), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n451), .A2(new_n368), .A3(new_n442), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT32), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT33), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G15gat), .B(G43gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(G71gat), .B(G99gat), .ZN(new_n457));
  XOR2_X1   g256(.A(new_n456), .B(new_n457), .Z(new_n458));
  NAND3_X1  g257(.A1(new_n453), .A2(new_n455), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n458), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n452), .B(KEYINPUT32), .C1(new_n454), .C2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n448), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT73), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n448), .A2(new_n459), .A3(KEYINPUT73), .A4(new_n461), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n459), .A2(new_n461), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT72), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n448), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n459), .A2(KEYINPUT72), .A3(new_n461), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT81), .ZN(new_n473));
  NOR2_X1   g272(.A1(G197gat), .A2(G204gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(G197gat), .A2(G204gat), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(G211gat), .A2(G218gat), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  OAI22_X1  g277(.A1(new_n474), .A2(new_n476), .B1(new_n478), .B2(KEYINPUT22), .ZN(new_n479));
  NOR2_X1   g278(.A1(G211gat), .A2(G218gat), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n478), .A2(new_n480), .A3(KEYINPUT74), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT74), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n331), .A2(new_n356), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n482), .B1(new_n483), .B2(new_n477), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n479), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT29), .ZN(new_n486));
  OR2_X1    g285(.A1(G197gat), .A2(G204gat), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT22), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n487), .A2(new_n475), .B1(new_n488), .B2(new_n477), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT74), .B1(new_n478), .B2(new_n480), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n483), .A2(new_n482), .A3(new_n477), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n485), .A2(new_n486), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT3), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(G162gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(G155gat), .ZN(new_n497));
  INV_X1    g296(.A(G155gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(G162gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G141gat), .B(G148gat), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n500), .B1(new_n501), .B2(KEYINPUT2), .ZN(new_n502));
  INV_X1    g301(.A(G148gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(G141gat), .ZN(new_n504));
  INV_X1    g303(.A(G141gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(G148gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G155gat), .B(G162gat), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT2), .B1(new_n498), .B2(KEYINPUT79), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n502), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n473), .B1(new_n495), .B2(new_n511), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n502), .A2(new_n510), .ZN(new_n513));
  AOI211_X1 g312(.A(KEYINPUT81), .B(new_n513), .C1(new_n493), .C2(new_n494), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n485), .A2(new_n492), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n513), .A2(new_n494), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n516), .B1(new_n486), .B2(new_n517), .ZN(new_n518));
  NOR3_X1   g317(.A1(new_n512), .A2(new_n514), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G228gat), .A2(G233gat), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT82), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n512), .ZN(new_n523));
  INV_X1    g322(.A(new_n518), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n495), .A2(new_n473), .A3(new_n511), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT82), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(new_n527), .A3(new_n520), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n516), .A2(KEYINPUT75), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n517), .A2(new_n486), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT75), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n529), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT83), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n495), .A2(new_n511), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT83), .A4(new_n532), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n535), .A2(new_n521), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n522), .A2(new_n528), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT85), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT85), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n522), .A2(new_n528), .A3(new_n541), .A4(new_n538), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n540), .A2(G22gat), .A3(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(G78gat), .B(G106gat), .Z(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT31), .ZN(new_n545));
  INV_X1    g344(.A(G50gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT84), .B(G22gat), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT86), .B1(new_n539), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n522), .A2(new_n528), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT86), .ZN(new_n551));
  INV_X1    g350(.A(new_n548), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .A4(new_n538), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n543), .A2(new_n547), .A3(new_n549), .A4(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT87), .ZN(new_n555));
  INV_X1    g354(.A(new_n547), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n539), .A2(new_n548), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n539), .A2(new_n548), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n554), .A2(new_n555), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n555), .B1(new_n554), .B2(new_n559), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n466), .B(new_n472), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n511), .A2(KEYINPUT3), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n382), .A2(new_n517), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT80), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n382), .A2(new_n511), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT4), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT4), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n569), .B1(new_n382), .B2(new_n511), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n382), .A2(KEYINPUT80), .A3(new_n517), .A4(new_n563), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n566), .A2(new_n568), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G225gat), .A2(G233gat), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT5), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n382), .B(new_n511), .ZN(new_n577));
  INV_X1    g376(.A(new_n573), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n574), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n567), .A2(new_n573), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n579), .B1(new_n572), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT0), .B(G57gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(G85gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(G1gat), .B(G29gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n584), .B(new_n585), .Z(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT6), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n576), .A2(new_n581), .A3(new_n586), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n589), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n586), .B1(new_n576), .B2(new_n581), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OR2_X1    g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n529), .A2(new_n532), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(G226gat), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n598), .A2(new_n328), .ZN(new_n599));
  OAI211_X1 g398(.A(new_n436), .B(new_n599), .C1(new_n402), .C2(new_n408), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n397), .B1(new_n433), .B2(new_n407), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT69), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n422), .B1(new_n603), .B2(new_n434), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n604), .B1(new_n409), .B2(new_n418), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n599), .A2(KEYINPUT29), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n597), .B(new_n600), .C1(new_n605), .C2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT76), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n606), .B1(new_n604), .B2(new_n416), .ZN(new_n611));
  INV_X1    g410(.A(new_n599), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n611), .B1(new_n449), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n516), .ZN(new_n614));
  XOR2_X1   g413(.A(G8gat), .B(G36gat), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(G64gat), .ZN(new_n616));
  INV_X1    g415(.A(G92gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n449), .A2(new_n606), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n620), .A2(KEYINPUT76), .A3(new_n597), .A4(new_n600), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n610), .A2(new_n614), .A3(new_n619), .A4(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT30), .ZN(new_n623));
  AOI21_X1  g422(.A(KEYINPUT78), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n622), .A2(KEYINPUT78), .A3(new_n623), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n610), .A2(new_n614), .A3(new_n621), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n618), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n629), .B1(new_n623), .B2(new_n622), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT77), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n622), .A2(new_n623), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT77), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n632), .A2(new_n633), .A3(new_n629), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n595), .A2(new_n627), .A3(new_n631), .A4(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT35), .B1(new_n562), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n626), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n632), .B(new_n629), .C1(new_n637), .C2(new_n624), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n591), .A2(new_n594), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n638), .A2(KEYINPUT35), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n554), .A2(new_n559), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT87), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n554), .A2(new_n555), .A3(new_n559), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n448), .B1(new_n461), .B2(new_n459), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n645), .B1(new_n464), .B2(new_n465), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n640), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n636), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT92), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT36), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n650), .B1(new_n466), .B2(new_n472), .ZN(new_n651));
  AOI211_X1 g450(.A(KEYINPUT36), .B(new_n645), .C1(new_n464), .C2(new_n465), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n635), .A2(new_n642), .A3(new_n643), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT88), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n605), .A2(new_n607), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n604), .A2(new_n612), .A3(new_n416), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n655), .B(new_n596), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n657), .B1(new_n449), .B2(new_n606), .ZN(new_n659));
  OAI21_X1  g458(.A(KEYINPUT88), .B1(new_n659), .B2(new_n597), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n515), .B(new_n611), .C1(new_n449), .C2(new_n612), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(KEYINPUT37), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT89), .B(KEYINPUT38), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT90), .B(KEYINPUT37), .Z(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n610), .A2(new_n614), .A3(new_n621), .A4(new_n667), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n663), .A2(new_n618), .A3(new_n665), .A4(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n622), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n628), .A2(KEYINPUT37), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n618), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT91), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n671), .A2(KEYINPUT91), .A3(new_n618), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n674), .A2(new_n668), .A3(new_n675), .ZN(new_n676));
  AOI211_X1 g475(.A(new_n595), .B(new_n670), .C1(new_n676), .C2(new_n664), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n572), .A2(new_n578), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n678), .A2(KEYINPUT39), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n678), .B(KEYINPUT39), .C1(new_n578), .C2(new_n577), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(new_n680), .A3(new_n586), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT40), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n683), .A2(new_n684), .A3(new_n593), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n638), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n686), .B1(new_n561), .B2(new_n560), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n653), .B(new_n654), .C1(new_n677), .C2(new_n687), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n648), .A2(new_n649), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n649), .B1(new_n648), .B2(new_n688), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n259), .B(new_n366), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n691), .A2(new_n595), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(new_n218), .ZN(G1324gat));
  INV_X1    g492(.A(new_n638), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT16), .B(G8gat), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT42), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n691), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n698), .A2(KEYINPUT110), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(KEYINPUT110), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(new_n691), .B2(new_n694), .ZN(new_n702));
  INV_X1    g501(.A(new_n259), .ZN(new_n703));
  AOI22_X1  g502(.A1(new_n642), .A2(new_n643), .B1(new_n638), .B2(new_n685), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n669), .A2(new_n622), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT91), .B1(new_n671), .B2(new_n618), .ZN(new_n706));
  AOI211_X1 g505(.A(new_n673), .B(new_n619), .C1(new_n628), .C2(KEYINPUT37), .ZN(new_n707));
  INV_X1    g506(.A(new_n668), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n639), .B(new_n705), .C1(new_n709), .C2(new_n665), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n704), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n466), .A2(new_n472), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT36), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n646), .A2(new_n650), .ZN(new_n714));
  AND4_X1   g513(.A1(new_n595), .A2(new_n627), .A3(new_n634), .A4(new_n631), .ZN(new_n715));
  OAI211_X1 g514(.A(new_n713), .B(new_n714), .C1(new_n715), .C2(new_n644), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n712), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n715), .A2(new_n718), .A3(new_n644), .ZN(new_n719));
  INV_X1    g518(.A(new_n645), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n466), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n721), .B1(new_n642), .B2(new_n643), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n719), .A2(KEYINPUT35), .B1(new_n722), .B2(new_n640), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT92), .B1(new_n717), .B2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n648), .A2(new_n688), .A3(new_n649), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n703), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n726), .A2(KEYINPUT108), .A3(new_n638), .A4(new_n366), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n702), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  AOI22_X1  g528(.A1(new_n699), .A2(new_n700), .B1(new_n729), .B2(G8gat), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n696), .ZN(new_n731));
  XOR2_X1   g530(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(KEYINPUT109), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n735));
  AOI211_X1 g534(.A(new_n735), .B(new_n732), .C1(new_n728), .C2(new_n696), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n730), .B1(new_n734), .B2(new_n736), .ZN(G1325gat));
  INV_X1    g536(.A(new_n691), .ZN(new_n738));
  AOI21_X1  g537(.A(G15gat), .B1(new_n738), .B2(new_n646), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n691), .A2(new_n653), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n739), .B1(G15gat), .B2(new_n740), .ZN(G1326gat));
  NOR2_X1   g540(.A1(new_n691), .A2(new_n644), .ZN(new_n742));
  XOR2_X1   g541(.A(KEYINPUT43), .B(G22gat), .Z(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1327gat));
  NAND2_X1  g543(.A1(new_n724), .A2(new_n725), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n364), .A2(new_n365), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n340), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(new_n310), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n648), .A2(new_n688), .ZN(new_n752));
  INV_X1    g551(.A(new_n746), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n747), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n749), .A2(new_n259), .A3(new_n751), .A4(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(G29gat), .B1(new_n756), .B2(new_n595), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n259), .B(new_n751), .C1(new_n689), .C2(new_n690), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n759), .A2(new_n595), .A3(new_n746), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n758), .B1(new_n760), .B2(new_n203), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n745), .A2(new_n259), .A3(new_n753), .A4(new_n751), .ZN(new_n762));
  NOR4_X1   g561(.A1(new_n762), .A2(KEYINPUT45), .A3(G29gat), .A4(new_n595), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n757), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT111), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT111), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n757), .B(new_n766), .C1(new_n761), .C2(new_n763), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1328gat));
  NOR3_X1   g567(.A1(new_n762), .A2(G36gat), .A3(new_n694), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT46), .ZN(new_n770));
  OR2_X1    g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(G36gat), .B1(new_n756), .B2(new_n694), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n769), .A2(new_n770), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(G1329gat));
  OAI21_X1  g573(.A(G43gat), .B1(new_n756), .B2(new_n653), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n759), .A2(new_n721), .A3(new_n746), .ZN(new_n777));
  INV_X1    g576(.A(G43gat), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR4_X1   g578(.A1(new_n762), .A2(KEYINPUT112), .A3(G43gat), .A4(new_n721), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n775), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT47), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n775), .B(KEYINPUT47), .C1(new_n779), .C2(new_n780), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(G1330gat));
  INV_X1    g584(.A(KEYINPUT48), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n546), .B1(new_n762), .B2(new_n644), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n756), .A2(new_n546), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n786), .B(new_n787), .C1(new_n788), .C2(new_n644), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n756), .A2(new_n546), .A3(new_n644), .ZN(new_n790));
  INV_X1    g589(.A(new_n787), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT48), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(G1331gat));
  NAND2_X1  g592(.A1(new_n746), .A2(new_n750), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(new_n259), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n752), .A2(new_n310), .A3(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n639), .B(KEYINPUT114), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g603(.A1(new_n800), .A2(new_n694), .ZN(new_n805));
  NOR2_X1   g604(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n806));
  AND2_X1   g605(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n805), .B2(new_n806), .ZN(G1333gat));
  INV_X1    g608(.A(G71gat), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n801), .A2(new_n810), .A3(new_n646), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n812));
  OAI21_X1  g611(.A(G71gat), .B1(new_n800), .B2(new_n653), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n812), .B1(new_n811), .B2(new_n813), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(G1334gat));
  INV_X1    g615(.A(new_n644), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(G78gat), .ZN(G1335gat));
  AOI22_X1  g618(.A1(new_n745), .A2(new_n748), .B1(new_n747), .B2(new_n754), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n750), .A2(new_n259), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n310), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n820), .A2(new_n639), .A3(new_n824), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n825), .A2(KEYINPUT115), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(KEYINPUT115), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(G85gat), .A3(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT51), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n754), .B2(new_n822), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n752), .A2(KEYINPUT51), .A3(new_n753), .A4(new_n821), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n823), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n595), .A2(G85gat), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n828), .B1(new_n833), .B2(new_n834), .ZN(G1336gat));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n820), .A2(G92gat), .A3(new_n638), .A4(new_n824), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(G92gat), .B1(new_n832), .B2(new_n638), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n836), .B(KEYINPUT52), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n832), .A2(new_n638), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n617), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n836), .A2(KEYINPUT52), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n836), .A2(KEYINPUT52), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n842), .A2(new_n843), .A3(new_n844), .A4(new_n837), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n840), .A2(new_n845), .ZN(G1337gat));
  INV_X1    g645(.A(new_n653), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n820), .A2(new_n847), .A3(new_n824), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(G99gat), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n830), .A2(new_n831), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n721), .A2(new_n823), .A3(G99gat), .ZN(new_n851));
  XOR2_X1   g650(.A(new_n851), .B(KEYINPUT117), .Z(new_n852));
  OAI21_X1  g651(.A(new_n849), .B1(new_n850), .B2(new_n852), .ZN(G1338gat));
  NAND3_X1  g652(.A1(new_n820), .A2(new_n817), .A3(new_n824), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(G106gat), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(KEYINPUT118), .ZN(new_n856));
  INV_X1    g655(.A(G106gat), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n832), .A2(new_n857), .A3(new_n817), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n856), .A2(new_n859), .A3(KEYINPUT53), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n855), .B(new_n858), .C1(KEYINPUT118), .C2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(new_n862), .ZN(G1339gat));
  NAND3_X1  g662(.A1(new_n288), .A2(new_n299), .A3(new_n295), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n298), .A2(new_n864), .A3(KEYINPUT54), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n299), .B1(new_n288), .B2(new_n295), .ZN(new_n866));
  XNOR2_X1  g665(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n308), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT55), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n865), .A2(new_n868), .A3(KEYINPUT55), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n871), .A2(new_n259), .A3(new_n309), .A4(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n227), .B1(new_n236), .B2(new_n237), .ZN(new_n874));
  INV_X1    g673(.A(new_n226), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n874), .B1(new_n875), .B2(new_n228), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n310), .B(new_n253), .C1(new_n248), .C2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n358), .ZN(new_n879));
  AOI21_X1  g678(.A(G218gat), .B1(new_n352), .B2(new_n354), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n362), .B1(new_n881), .B2(KEYINPUT100), .ZN(new_n882));
  INV_X1    g681(.A(new_n365), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n878), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n871), .A2(new_n309), .A3(new_n872), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n253), .B1(new_n248), .B2(new_n876), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n364), .A3(new_n365), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  AOI22_X1  g688(.A1(new_n889), .A2(new_n340), .B1(new_n366), .B2(new_n703), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n890), .A2(new_n817), .A3(new_n721), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n638), .A2(new_n595), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(G113gat), .B1(new_n893), .B2(new_n703), .ZN(new_n894));
  INV_X1    g693(.A(new_n890), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n802), .A2(new_n694), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n562), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n703), .A2(new_n372), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n894), .B1(new_n899), .B2(new_n900), .ZN(G1340gat));
  OAI21_X1  g700(.A(G120gat), .B1(new_n893), .B2(new_n823), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n823), .A2(new_n375), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n899), .B2(new_n903), .ZN(G1341gat));
  INV_X1    g703(.A(G127gat), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n893), .A2(new_n905), .A3(new_n340), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n897), .A2(new_n898), .A3(new_n750), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(new_n905), .ZN(G1342gat));
  NOR3_X1   g707(.A1(new_n899), .A2(G134gat), .A3(new_n746), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT56), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  OAI21_X1  g711(.A(G134gat), .B1(new_n893), .B2(new_n746), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(G1343gat));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n871), .A2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n309), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT55), .B1(new_n865), .B2(new_n868), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(KEYINPUT120), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n916), .A2(new_n919), .A3(new_n259), .A4(new_n872), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n877), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n746), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n750), .B1(new_n922), .B2(new_n888), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n794), .A2(new_n259), .A3(new_n310), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n817), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT57), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT57), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n895), .A2(new_n927), .A3(new_n817), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n653), .A2(new_n892), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n926), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(G141gat), .B1(new_n930), .B2(new_n703), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n847), .A2(new_n644), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n895), .A2(new_n896), .A3(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n934), .A2(new_n505), .A3(new_n259), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT58), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n937), .B1(new_n935), .B2(KEYINPUT121), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n931), .B(new_n935), .C1(KEYINPUT121), .C2(new_n937), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1344gat));
  INV_X1    g740(.A(KEYINPUT59), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n942), .B(G148gat), .C1(new_n930), .C2(new_n823), .ZN(new_n943));
  OAI21_X1  g742(.A(KEYINPUT57), .B1(new_n890), .B2(new_n644), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n927), .B(new_n817), .C1(new_n923), .C2(new_n924), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n944), .A2(new_n945), .A3(new_n310), .A4(new_n929), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(G148gat), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT122), .B1(new_n947), .B2(KEYINPUT59), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT122), .ZN(new_n949));
  AOI211_X1 g748(.A(new_n949), .B(new_n942), .C1(new_n946), .C2(G148gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n943), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n934), .A2(new_n503), .A3(new_n310), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1345gat));
  XNOR2_X1  g752(.A(KEYINPUT79), .B(G155gat), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n930), .A2(new_n340), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n934), .A2(new_n750), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n955), .B1(new_n954), .B2(new_n956), .ZN(G1346gat));
  AOI21_X1  g756(.A(G162gat), .B1(new_n934), .B2(new_n753), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n930), .A2(new_n496), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n958), .B1(new_n959), .B2(new_n753), .ZN(G1347gat));
  NOR2_X1   g759(.A1(new_n802), .A2(new_n694), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n891), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(G169gat), .B1(new_n962), .B2(new_n703), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n890), .A2(new_n639), .A3(new_n694), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(new_n898), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n259), .A2(new_n384), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(G1348gat));
  INV_X1    g766(.A(new_n962), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n968), .A2(G176gat), .A3(new_n310), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n969), .A2(KEYINPUT123), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n969), .A2(KEYINPUT123), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n965), .A2(new_n823), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n972), .A2(G176gat), .ZN(new_n973));
  NOR3_X1   g772(.A1(new_n970), .A2(new_n971), .A3(new_n973), .ZN(G1349gat));
  OAI21_X1  g773(.A(G183gat), .B1(new_n962), .B2(new_n340), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n750), .A2(new_n420), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n975), .B1(new_n965), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(KEYINPUT60), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT60), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n975), .B(new_n979), .C1(new_n965), .C2(new_n976), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(G1350gat));
  NAND2_X1  g780(.A1(new_n968), .A2(new_n753), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(G190gat), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT61), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n983), .A2(KEYINPUT124), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(KEYINPUT124), .ZN(new_n986));
  OR2_X1    g785(.A1(new_n984), .A2(KEYINPUT124), .ZN(new_n987));
  NAND4_X1  g786(.A1(new_n982), .A2(G190gat), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n964), .A2(new_n353), .A3(new_n898), .A4(new_n753), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n985), .A2(new_n988), .A3(new_n989), .ZN(G1351gat));
  NAND2_X1  g789(.A1(new_n964), .A2(new_n932), .ZN(new_n991));
  NOR3_X1   g790(.A1(new_n991), .A2(G197gat), .A3(new_n703), .ZN(new_n992));
  XNOR2_X1  g791(.A(new_n992), .B(KEYINPUT125), .ZN(new_n993));
  AND2_X1   g792(.A1(new_n961), .A2(new_n653), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n944), .A2(new_n945), .A3(new_n994), .ZN(new_n995));
  OAI21_X1  g794(.A(G197gat), .B1(new_n995), .B2(new_n703), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n993), .A2(new_n996), .ZN(G1352gat));
  NOR3_X1   g796(.A1(new_n991), .A2(G204gat), .A3(new_n823), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT62), .ZN(new_n999));
  OR2_X1    g798(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n998), .A2(new_n999), .ZN(new_n1001));
  AND4_X1   g800(.A1(new_n310), .A2(new_n944), .A3(new_n945), .A4(new_n994), .ZN(new_n1002));
  OAI211_X1 g801(.A(new_n1000), .B(new_n1001), .C1(new_n305), .C2(new_n1002), .ZN(G1353gat));
  OAI21_X1  g802(.A(G211gat), .B1(new_n995), .B2(new_n340), .ZN(new_n1004));
  NAND2_X1  g803(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n1005));
  OR2_X1    g804(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g806(.A(new_n991), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n1008), .A2(new_n331), .A3(new_n750), .ZN(new_n1009));
  OAI211_X1 g808(.A(new_n1007), .B(new_n1009), .C1(new_n1004), .C2(new_n1006), .ZN(G1354gat));
  OAI21_X1  g809(.A(G218gat), .B1(new_n995), .B2(new_n746), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n753), .A2(new_n356), .ZN(new_n1012));
  OAI21_X1  g811(.A(new_n1011), .B1(new_n991), .B2(new_n1012), .ZN(G1355gat));
endmodule


