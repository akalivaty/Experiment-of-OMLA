//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980;
  INV_X1    g000(.A(G227gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(KEYINPUT27), .B(G183gat), .ZN(new_n208));
  INV_X1    g007(.A(G190gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n207), .B1(new_n210), .B2(KEYINPUT28), .ZN(new_n211));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT26), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT68), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI211_X1 g016(.A(KEYINPUT68), .B(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n213), .A2(new_n214), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT28), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n208), .A2(new_n221), .A3(new_n209), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n211), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n213), .ZN(new_n224));
  NOR2_X1   g023(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n212), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g025(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n227));
  NAND2_X1  g026(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n213), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NOR3_X1   g028(.A1(new_n226), .A2(new_n229), .A3(KEYINPUT25), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT64), .B1(new_n207), .B2(KEYINPUT24), .ZN(new_n231));
  INV_X1    g030(.A(G183gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n232), .A2(new_n209), .A3(KEYINPUT65), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(G183gat), .B2(G190gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT64), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT24), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n206), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n207), .A2(KEYINPUT24), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n231), .A2(new_n236), .A3(new_n239), .A4(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n230), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n228), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(new_n224), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n206), .A2(new_n245), .A3(new_n238), .ZN(new_n246));
  OAI211_X1 g045(.A(G183gat), .B(G190gat), .C1(KEYINPUT67), .C2(KEYINPUT24), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n209), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n227), .A2(new_n213), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n244), .A2(new_n249), .A3(new_n212), .A4(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(KEYINPUT25), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n223), .A2(new_n242), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G113gat), .ZN(new_n254));
  INV_X1    g053(.A(G120gat), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT1), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n256), .B1(new_n254), .B2(new_n255), .ZN(new_n257));
  XNOR2_X1  g056(.A(G127gat), .B(G134gat), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT69), .B(G113gat), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n256), .B(new_n258), .C1(new_n261), .C2(new_n255), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n253), .A2(new_n264), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n230), .A2(new_n241), .B1(new_n251), .B2(KEYINPUT25), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n263), .B1(new_n266), .B2(new_n223), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n205), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT73), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(new_n269), .A3(KEYINPUT34), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT34), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n271), .B(new_n205), .C1(new_n265), .C2(new_n267), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT74), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n253), .A2(new_n264), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n266), .A2(new_n263), .A3(new_n223), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n204), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(KEYINPUT73), .B1(new_n277), .B2(new_n271), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(KEYINPUT74), .A3(new_n271), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n270), .A2(new_n274), .A3(new_n278), .A4(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT72), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n275), .A2(new_n276), .A3(new_n204), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT33), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT70), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n282), .A2(new_n286), .A3(new_n283), .ZN(new_n287));
  XNOR2_X1  g086(.A(G15gat), .B(G43gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(G71gat), .B(G99gat), .ZN(new_n289));
  XOR2_X1   g088(.A(new_n288), .B(new_n289), .Z(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n291), .B1(new_n282), .B2(KEYINPUT32), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n285), .A2(new_n287), .A3(new_n292), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n291), .A2(KEYINPUT71), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n291), .A2(KEYINPUT71), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(KEYINPUT33), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n282), .A2(KEYINPUT32), .A3(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n293), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n293), .A2(new_n297), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n299), .A2(KEYINPUT72), .A3(new_n280), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(G78gat), .B(G106gat), .Z(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT31), .B(G50gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G22gat), .ZN(new_n305));
  INV_X1    g104(.A(G228gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n306), .A2(new_n203), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G211gat), .ZN(new_n309));
  INV_X1    g108(.A(G218gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G211gat), .A2(G218gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G197gat), .B(G204gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT76), .B(KEYINPUT22), .ZN(new_n315));
  INV_X1    g114(.A(new_n312), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n313), .B(new_n314), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(KEYINPUT82), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n318), .A2(KEYINPUT29), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n320));
  INV_X1    g119(.A(new_n313), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n322), .A2(KEYINPUT82), .A3(new_n317), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT3), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G141gat), .B(G148gat), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G155gat), .ZN(new_n327));
  INV_X1    g126(.A(G162gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G155gat), .A2(G162gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(KEYINPUT2), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n326), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n330), .B(new_n329), .C1(new_n325), .C2(KEYINPUT2), .ZN(new_n334));
  AND2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n324), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n322), .A2(new_n317), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT77), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n322), .A2(KEYINPUT77), .A3(new_n317), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n333), .A2(new_n334), .A3(new_n342), .ZN(new_n343));
  AOI22_X1  g142(.A1(new_n339), .A2(new_n340), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n308), .B1(new_n336), .B2(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(new_n308), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n333), .A2(new_n334), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT29), .B1(new_n322), .B2(new_n317), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n347), .B1(new_n348), .B2(KEYINPUT3), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n305), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT83), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n304), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n319), .A2(new_n323), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n347), .B1(new_n354), .B2(KEYINPUT3), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n343), .A2(new_n341), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n307), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n358), .A2(new_n307), .A3(new_n349), .ZN(new_n360));
  OAI21_X1  g159(.A(G22gat), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n350), .A3(new_n305), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n353), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n361), .A2(new_n362), .A3(new_n352), .A4(new_n304), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT86), .B1(new_n301), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n358), .B1(new_n335), .B2(new_n324), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n368), .A2(new_n308), .B1(new_n346), .B2(new_n349), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT83), .B1(new_n369), .B2(new_n305), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n370), .A2(new_n304), .B1(new_n362), .B2(new_n361), .ZN(new_n371));
  INV_X1    g170(.A(new_n365), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT86), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n373), .A2(new_n374), .A3(new_n298), .A4(new_n300), .ZN(new_n375));
  AOI22_X1  g174(.A1(new_n347), .A2(KEYINPUT3), .B1(new_n260), .B2(new_n262), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n343), .ZN(new_n377));
  NAND2_X1  g176(.A1(G225gat), .A2(G233gat), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT4), .B1(new_n347), .B2(new_n263), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NOR3_X1   g179(.A1(new_n347), .A2(new_n263), .A3(KEYINPUT4), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n377), .B(new_n378), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT5), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(G1gat), .B(G29gat), .ZN(new_n385));
  INV_X1    g184(.A(G85gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT0), .B(G57gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n264), .A2(new_n335), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n347), .A2(new_n263), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n378), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT4), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n264), .A2(new_n335), .A3(new_n394), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n395), .A2(new_n379), .B1(new_n376), .B2(new_n343), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n393), .B1(new_n396), .B2(new_n378), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n384), .B(new_n390), .C1(new_n397), .C2(new_n383), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n393), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n383), .B1(new_n382), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT5), .B1(new_n396), .B2(new_n378), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n389), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT6), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n399), .B1(new_n405), .B2(KEYINPUT81), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n384), .B1(new_n397), .B2(new_n383), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT6), .B1(new_n407), .B2(new_n389), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT81), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n398), .A2(new_n404), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(G226gat), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n414), .A2(new_n203), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n253), .A2(new_n341), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n266), .A2(new_n223), .A3(new_n415), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n356), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT78), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT78), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n417), .A2(new_n356), .A3(new_n421), .A4(new_n418), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n356), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n253), .A2(new_n416), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n416), .A2(new_n341), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n426), .B1(new_n266), .B2(new_n223), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n424), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT79), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT79), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n430), .B(new_n424), .C1(new_n425), .C2(new_n427), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n423), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT30), .ZN(new_n434));
  XNOR2_X1  g233(.A(G64gat), .B(G92gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n435), .B(KEYINPUT80), .ZN(new_n436));
  XNOR2_X1  g235(.A(G8gat), .B(G36gat), .ZN(new_n437));
  XOR2_X1   g236(.A(new_n436), .B(new_n437), .Z(new_n438));
  NAND3_X1  g237(.A1(new_n433), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n438), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n440), .B1(new_n423), .B2(new_n432), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n420), .A2(new_n422), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n442), .A2(new_n438), .A3(new_n429), .A4(new_n431), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n441), .A2(KEYINPUT30), .A3(new_n443), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n411), .A2(new_n413), .B1(new_n439), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n367), .A2(new_n375), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT35), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n299), .A2(KEYINPUT75), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT75), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n293), .A2(new_n449), .A3(new_n297), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n280), .A3(new_n450), .ZN(new_n451));
  AND4_X1   g250(.A1(new_n270), .A2(new_n274), .A3(new_n278), .A4(new_n279), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n299), .A2(new_n452), .A3(KEYINPUT75), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n444), .A2(new_n439), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n408), .A2(new_n398), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT35), .B1(new_n457), .B2(new_n413), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n373), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n447), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT84), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n366), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n364), .A2(KEYINPUT84), .A3(new_n365), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n444), .A2(new_n439), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n412), .B1(new_n406), .B2(new_n410), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n464), .B(new_n465), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n391), .A2(new_n378), .A3(new_n392), .ZN(new_n469));
  OAI211_X1 g268(.A(KEYINPUT39), .B(new_n469), .C1(new_n396), .C2(new_n378), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n377), .B1(new_n380), .B2(new_n381), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT39), .ZN(new_n472));
  INV_X1    g271(.A(new_n378), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n470), .A2(new_n474), .A3(new_n389), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT85), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT40), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n398), .B1(new_n475), .B2(new_n477), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n476), .B1(new_n475), .B2(new_n477), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n481), .A2(new_n439), .A3(new_n444), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT38), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT37), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n438), .B1(new_n433), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n442), .A2(new_n429), .A3(new_n431), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT37), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n483), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n428), .A2(new_n419), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT38), .B1(new_n489), .B2(KEYINPUT37), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n440), .B(new_n490), .C1(new_n486), .C2(KEYINPUT37), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n491), .A2(new_n413), .A3(new_n443), .A4(new_n457), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n482), .B(new_n373), .C1(new_n488), .C2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT36), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n451), .A2(new_n494), .A3(new_n453), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n298), .A2(KEYINPUT36), .A3(new_n300), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n468), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n462), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(G50gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(G43gat), .ZN(new_n501));
  INV_X1    g300(.A(G43gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(G50gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n501), .A2(new_n503), .A3(KEYINPUT15), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(KEYINPUT92), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NOR3_X1   g306(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n508));
  OR2_X1    g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT91), .B(G36gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(G29gat), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n501), .A2(new_n503), .A3(KEYINPUT93), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT15), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n512), .B(new_n513), .C1(KEYINPUT93), .C2(new_n501), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n505), .A2(new_n509), .A3(new_n511), .A4(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT90), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n507), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n511), .B(new_n517), .C1(new_n509), .C2(new_n516), .ZN(new_n518));
  INV_X1    g317(.A(new_n504), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT17), .ZN(new_n522));
  XOR2_X1   g321(.A(G15gat), .B(G22gat), .Z(new_n523));
  INV_X1    g322(.A(G1gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT94), .ZN(new_n526));
  AOI21_X1  g325(.A(G8gat), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n524), .A2(KEYINPUT16), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n525), .B1(new_n528), .B2(new_n523), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n527), .B(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n520), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n522), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(G229gat), .A2(G233gat), .ZN(new_n535));
  INV_X1    g334(.A(new_n530), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(new_n531), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n534), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT18), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n534), .A2(KEYINPUT18), .A3(new_n535), .A4(new_n537), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT95), .B1(new_n521), .B2(new_n530), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n537), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n535), .B(KEYINPUT13), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n536), .A2(KEYINPUT95), .A3(new_n531), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n543), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n540), .A2(new_n541), .A3(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G113gat), .B(G141gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT88), .B(KEYINPUT89), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(G169gat), .B(G197gat), .Z(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT12), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n548), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n557), .A2(new_n540), .A3(new_n541), .A4(new_n547), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT96), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n560), .A2(new_n561), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n559), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(G57gat), .B(G64gat), .Z(new_n565));
  INV_X1    g364(.A(KEYINPUT97), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT9), .ZN(new_n567));
  INV_X1    g366(.A(G71gat), .ZN(new_n568));
  INV_X1    g367(.A(G78gat), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n565), .A2(new_n566), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G71gat), .B(G78gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n571), .B(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT102), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT7), .ZN(new_n576));
  OAI211_X1 g375(.A(G85gat), .B(G92gat), .C1(new_n576), .C2(KEYINPUT101), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT101), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n578), .A2(KEYINPUT7), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n575), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(KEYINPUT101), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(KEYINPUT7), .ZN(new_n582));
  AND2_X1   g381(.A1(G85gat), .A2(G92gat), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n581), .A2(new_n582), .A3(new_n583), .A4(KEYINPUT102), .ZN(new_n584));
  INV_X1    g383(.A(G92gat), .ZN(new_n585));
  OAI21_X1  g384(.A(KEYINPUT7), .B1(new_n386), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n580), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G99gat), .B(G106gat), .ZN(new_n588));
  XOR2_X1   g387(.A(KEYINPUT103), .B(G85gat), .Z(new_n589));
  NAND2_X1  g388(.A1(G99gat), .A2(G106gat), .ZN(new_n590));
  AOI22_X1  g389(.A1(new_n589), .A2(new_n585), .B1(KEYINPUT8), .B2(new_n590), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n587), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n588), .B1(new_n587), .B2(new_n591), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n574), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n587), .A2(new_n591), .ZN(new_n595));
  INV_X1    g394(.A(new_n588), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n571), .A2(new_n573), .ZN(new_n598));
  INV_X1    g397(.A(G64gat), .ZN(new_n599));
  OR2_X1    g398(.A1(new_n599), .A2(G57gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(G57gat), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT97), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n572), .B1(new_n602), .B2(new_n570), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n587), .A2(new_n588), .A3(new_n591), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n597), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT10), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n594), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n592), .A2(new_n593), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n609), .A2(KEYINPUT10), .A3(new_n604), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G230gat), .A2(G233gat), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT107), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT107), .ZN(new_n614));
  INV_X1    g413(.A(new_n612), .ZN(new_n615));
  AOI211_X1 g414(.A(new_n614), .B(new_n615), .C1(new_n608), .C2(new_n610), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n594), .A2(new_n606), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n615), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G120gat), .B(G148gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(G176gat), .B(G204gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n623), .B(KEYINPUT106), .Z(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT105), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n615), .B1(new_n611), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n627), .B1(new_n626), .B2(new_n611), .ZN(new_n628));
  INV_X1    g427(.A(new_n623), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n628), .A2(new_n629), .A3(new_n619), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT21), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n574), .B1(new_n530), .B2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G127gat), .B(G155gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G231gat), .A2(G233gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT98), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(new_n232), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(new_n309), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n636), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n530), .A2(new_n633), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n643));
  XOR2_X1   g442(.A(new_n642), .B(new_n643), .Z(new_n644));
  OR2_X1    g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n641), .A2(new_n644), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n522), .B(new_n533), .C1(new_n592), .C2(new_n593), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n609), .A2(new_n531), .ZN(new_n650));
  NAND2_X1  g449(.A1(G232gat), .A2(G233gat), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n651), .B(KEYINPUT99), .Z(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(KEYINPUT41), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n649), .A2(new_n650), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G190gat), .B(G218gat), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n656), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n649), .A2(new_n650), .A3(new_n654), .A4(new_n658), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n653), .A2(KEYINPUT41), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(new_n328), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT100), .B(G134gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(KEYINPUT104), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n664), .B(KEYINPUT104), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n666), .B1(new_n660), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n648), .A2(new_n669), .ZN(new_n670));
  AND4_X1   g469(.A1(new_n499), .A2(new_n564), .A3(new_n632), .A4(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n467), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n466), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT16), .B(G8gat), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n677), .B(KEYINPUT109), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n674), .B(KEYINPUT108), .ZN(new_n679));
  INV_X1    g478(.A(new_n676), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n675), .ZN(new_n682));
  INV_X1    g481(.A(G8gat), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n678), .B(new_n682), .C1(new_n683), .C2(new_n679), .ZN(G1325gat));
  AOI21_X1  g483(.A(G15gat), .B1(new_n671), .B2(new_n454), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n497), .A2(KEYINPUT110), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n497), .A2(KEYINPUT110), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n688), .A2(G15gat), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n685), .B1(new_n671), .B2(new_n689), .ZN(G1326gat));
  AND2_X1   g489(.A1(new_n464), .A2(new_n465), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n671), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT43), .B(G22gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1327gat));
  AOI21_X1  g493(.A(new_n668), .B1(new_n462), .B2(new_n498), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n564), .A2(new_n632), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n696), .A2(new_n647), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(G29gat), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n699), .A2(new_n700), .A3(new_n467), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT45), .ZN(new_n702));
  INV_X1    g501(.A(new_n467), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n668), .A2(KEYINPUT44), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT112), .B1(new_n462), .B2(new_n498), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n460), .B1(new_n446), .B2(KEYINPUT35), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n468), .A2(new_n493), .A3(new_n497), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT112), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n704), .B1(new_n705), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711));
  OAI21_X1  g510(.A(KEYINPUT111), .B1(new_n695), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n669), .B1(new_n706), .B2(new_n707), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT111), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n713), .A2(new_n714), .A3(KEYINPUT44), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n710), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(KEYINPUT113), .B1(new_n716), .B2(new_n697), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n716), .A2(KEYINPUT113), .A3(new_n697), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n703), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n702), .B1(new_n720), .B2(new_n700), .ZN(G1328gat));
  INV_X1    g520(.A(new_n510), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n699), .A2(new_n466), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT46), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT114), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n456), .B1(new_n718), .B2(new_n719), .ZN(new_n726));
  OAI221_X1 g525(.A(new_n725), .B1(KEYINPUT46), .B2(new_n723), .C1(new_n726), .C2(new_n722), .ZN(G1329gat));
  NOR3_X1   g526(.A1(new_n698), .A2(G43gat), .A3(new_n455), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n716), .ZN(new_n731));
  NOR4_X1   g530(.A1(new_n731), .A2(new_n497), .A3(new_n696), .A4(new_n647), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n732), .B2(new_n502), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n716), .A2(KEYINPUT113), .A3(new_n697), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n688), .B1(new_n734), .B2(new_n717), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n728), .B1(new_n735), .B2(G43gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n733), .B1(new_n736), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g536(.A1(new_n716), .A2(new_n366), .A3(new_n697), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n738), .A2(KEYINPUT48), .A3(G50gat), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n699), .A2(new_n500), .A3(new_n691), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT115), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n739), .B(new_n740), .C1(new_n741), .C2(KEYINPUT48), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n691), .B1(new_n734), .B2(new_n717), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n743), .B1(new_n744), .B2(G50gat), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n742), .B1(new_n745), .B2(KEYINPUT48), .ZN(G1331gat));
  OR2_X1    g545(.A1(new_n705), .A2(new_n709), .ZN(new_n747));
  INV_X1    g546(.A(new_n564), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n670), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n749), .A2(new_n632), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n467), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g553(.A1(new_n751), .A2(new_n456), .ZN(new_n755));
  NOR2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  AND2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n755), .B2(new_n756), .ZN(G1333gat));
  INV_X1    g558(.A(new_n688), .ZN(new_n760));
  OAI21_X1  g559(.A(G71gat), .B1(new_n751), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n454), .A2(new_n568), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(new_n751), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n763), .B(new_n764), .ZN(G1334gat));
  NAND2_X1  g564(.A1(new_n752), .A2(new_n691), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g566(.A1(new_n748), .A2(new_n648), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n695), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n772), .A2(new_n631), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n467), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n768), .A2(new_n632), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n731), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n703), .A2(new_n589), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n774), .A2(new_n589), .B1(new_n777), .B2(new_n778), .ZN(G1336gat));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n466), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G92gat), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n632), .A2(new_n456), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n783), .A2(G92gat), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT52), .B1(new_n772), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n770), .A2(KEYINPUT117), .A3(new_n771), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n771), .A2(KEYINPUT117), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n695), .A2(new_n769), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  AOI22_X1  g589(.A1(new_n780), .A2(G92gat), .B1(new_n784), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n786), .B1(new_n791), .B2(new_n792), .ZN(G1337gat));
  XOR2_X1   g592(.A(KEYINPUT118), .B(G99gat), .Z(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n773), .A2(new_n454), .A3(new_n795), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n731), .A2(new_n760), .A3(new_n776), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n797), .B2(new_n795), .ZN(G1338gat));
  NAND2_X1  g597(.A1(new_n777), .A2(new_n366), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(G106gat), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n373), .A2(G106gat), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT53), .B1(new_n773), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n631), .ZN(new_n804));
  AOI211_X1 g603(.A(KEYINPUT119), .B(new_n804), .C1(new_n787), .C2(new_n789), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT119), .ZN(new_n806));
  INV_X1    g605(.A(new_n804), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n806), .B1(new_n790), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n716), .A2(new_n691), .A3(new_n775), .ZN(new_n809));
  AOI211_X1 g608(.A(new_n805), .B(new_n808), .C1(G106gat), .C2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n803), .B1(new_n810), .B2(new_n811), .ZN(G1339gat));
  OAI211_X1 g611(.A(new_n628), .B(KEYINPUT54), .C1(new_n611), .C2(new_n612), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n613), .B2(new_n616), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n815), .A2(KEYINPUT121), .A3(new_n623), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT121), .B1(new_n815), .B2(new_n623), .ZN(new_n817));
  OAI211_X1 g616(.A(KEYINPUT55), .B(new_n813), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n630), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(KEYINPUT122), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT122), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n818), .A2(new_n821), .A3(new_n630), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n815), .A2(new_n623), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT121), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n815), .A2(KEYINPUT121), .A3(new_n623), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n813), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n820), .A2(new_n564), .A3(new_n822), .A4(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n562), .A2(new_n563), .ZN(new_n832));
  INV_X1    g631(.A(new_n555), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n545), .B1(new_n543), .B2(new_n546), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n535), .B1(new_n534), .B2(new_n537), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n631), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n669), .B1(new_n831), .B2(new_n839), .ZN(new_n840));
  AOI22_X1  g639(.A1(new_n819), .A2(KEYINPUT122), .B1(new_n828), .B2(new_n829), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n832), .A2(new_n668), .A3(new_n837), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(new_n822), .A3(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n648), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n670), .A2(new_n748), .A3(new_n632), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT120), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n846), .B(new_n847), .ZN(new_n848));
  AOI211_X1 g647(.A(new_n455), .B(new_n691), .C1(new_n845), .C2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n703), .A2(new_n466), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(G113gat), .B1(new_n851), .B2(new_n748), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n703), .B1(new_n845), .B2(new_n848), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n367), .A2(new_n375), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n853), .A2(new_n855), .A3(new_n456), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n261), .A3(new_n564), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n852), .A2(new_n857), .ZN(G1340gat));
  OAI21_X1  g657(.A(G120gat), .B1(new_n851), .B2(new_n632), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n856), .A2(new_n255), .A3(new_n631), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(G1341gat));
  INV_X1    g660(.A(G127gat), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n851), .A2(new_n862), .A3(new_n648), .ZN(new_n863));
  AOI21_X1  g662(.A(G127gat), .B1(new_n856), .B2(new_n647), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n863), .A2(new_n864), .ZN(G1342gat));
  OAI21_X1  g664(.A(G134gat), .B1(new_n851), .B2(new_n668), .ZN(new_n866));
  INV_X1    g665(.A(G134gat), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n668), .A2(new_n466), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n853), .A2(new_n867), .A3(new_n855), .A4(new_n868), .ZN(new_n869));
  XNOR2_X1  g668(.A(KEYINPUT123), .B(KEYINPUT56), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n866), .A2(new_n871), .A3(new_n872), .ZN(G1343gat));
  AND2_X1   g672(.A1(new_n850), .A2(new_n497), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n845), .A2(new_n848), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT57), .B1(new_n875), .B2(new_n366), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n691), .A2(KEYINPUT57), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n830), .A2(new_n564), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n839), .B1(new_n878), .B2(new_n819), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n668), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n647), .B1(new_n880), .B2(new_n843), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n877), .B1(new_n882), .B2(new_n848), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n564), .B(new_n874), .C1(new_n876), .C2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(G141gat), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n688), .A2(new_n373), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n748), .A2(G141gat), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n853), .A2(new_n456), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT124), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT58), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n885), .A2(new_n888), .A3(new_n892), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1344gat));
  AND2_X1   g695(.A1(new_n853), .A2(new_n886), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n632), .A2(G148gat), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n897), .A2(new_n456), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n874), .B1(new_n876), .B2(new_n883), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n900), .A2(new_n632), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(G148gat), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n875), .A2(new_n366), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT57), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT57), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n749), .A2(new_n631), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n907), .B(new_n691), .C1(new_n881), .C2(new_n908), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n906), .A2(new_n631), .A3(new_n874), .A4(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n902), .B1(new_n910), .B2(G148gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n899), .B1(new_n904), .B2(new_n911), .ZN(G1345gat));
  NOR3_X1   g711(.A1(new_n900), .A2(new_n327), .A3(new_n648), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n897), .A2(new_n456), .A3(new_n647), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n327), .B2(new_n914), .ZN(G1346gat));
  OAI21_X1  g714(.A(G162gat), .B1(new_n900), .B2(new_n668), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n897), .A2(new_n328), .A3(new_n868), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1347gat));
  NOR2_X1   g717(.A1(new_n467), .A2(new_n456), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n849), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(G169gat), .B1(new_n920), .B2(new_n748), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n875), .A2(new_n703), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT125), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n854), .A2(new_n456), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n748), .A2(G169gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n921), .B1(new_n925), .B2(new_n926), .ZN(G1348gat));
  OAI21_X1  g726(.A(G176gat), .B1(new_n920), .B2(new_n632), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n632), .A2(G176gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n928), .B1(new_n925), .B2(new_n929), .ZN(G1349gat));
  AND2_X1   g729(.A1(new_n647), .A2(new_n208), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n922), .A2(KEYINPUT125), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT125), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n933), .B1(new_n875), .B2(new_n703), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n924), .B(new_n931), .C1(new_n932), .C2(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(G183gat), .B1(new_n920), .B2(new_n648), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(KEYINPUT60), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT60), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n935), .A2(new_n936), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(G1350gat));
  NOR2_X1   g740(.A1(new_n668), .A2(G190gat), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n924), .B(new_n942), .C1(new_n932), .C2(new_n934), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n943), .A2(KEYINPUT126), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n943), .A2(KEYINPUT126), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n849), .A2(new_n669), .A3(new_n919), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(G190gat), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n947), .A2(KEYINPUT61), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n947), .A2(KEYINPUT61), .ZN(new_n949));
  OAI22_X1  g748(.A1(new_n944), .A2(new_n945), .B1(new_n948), .B2(new_n949), .ZN(G1351gat));
  NOR3_X1   g749(.A1(new_n688), .A2(new_n467), .A3(new_n456), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n373), .B1(new_n845), .B2(new_n848), .ZN(new_n952));
  OAI211_X1 g751(.A(new_n909), .B(new_n951), .C1(new_n952), .C2(new_n907), .ZN(new_n953));
  OAI21_X1  g752(.A(G197gat), .B1(new_n953), .B2(new_n748), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n923), .A2(new_n466), .A3(new_n886), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n748), .A2(G197gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(G1352gat));
  NOR2_X1   g756(.A1(new_n783), .A2(G204gat), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n923), .A2(new_n886), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT62), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n923), .A2(new_n961), .A3(new_n886), .A4(new_n958), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n906), .A2(new_n631), .A3(new_n909), .ZN(new_n963));
  INV_X1    g762(.A(new_n951), .ZN(new_n964));
  OAI21_X1  g763(.A(G204gat), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n960), .A2(new_n962), .A3(new_n965), .ZN(G1353gat));
  OAI211_X1 g765(.A(KEYINPUT63), .B(G211gat), .C1(new_n953), .C2(new_n648), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(KEYINPUT127), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n906), .A2(new_n647), .A3(new_n909), .A4(new_n951), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n969), .A2(new_n970), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n971));
  OAI21_X1  g770(.A(G211gat), .B1(new_n953), .B2(new_n648), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT63), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n968), .A2(new_n971), .A3(new_n974), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n648), .A2(G211gat), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n923), .A2(new_n466), .A3(new_n886), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n975), .A2(new_n977), .ZN(G1354gat));
  NOR3_X1   g777(.A1(new_n953), .A2(new_n310), .A3(new_n668), .ZN(new_n979));
  NAND4_X1  g778(.A1(new_n923), .A2(new_n466), .A3(new_n669), .A4(new_n886), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n979), .B1(new_n980), .B2(new_n310), .ZN(G1355gat));
endmodule


