

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U554 ( .A(KEYINPUT1), .B(n532), .Z(n790) );
  NOR2_X1 U555 ( .A1(G651), .A2(n547), .ZN(n789) );
  OR2_X1 U556 ( .A1(n663), .A2(n662), .ZN(n698) );
  AND2_X1 U557 ( .A1(n526), .A2(G2104), .ZN(n878) );
  XOR2_X1 U558 ( .A(KEYINPUT64), .B(n689), .Z(n519) );
  XNOR2_X1 U559 ( .A(KEYINPUT110), .B(n754), .ZN(n520) );
  AND2_X1 U560 ( .A1(n741), .A2(n740), .ZN(n521) );
  NAND2_X1 U561 ( .A1(n708), .A2(n707), .ZN(n522) );
  NOR2_X1 U562 ( .A1(n618), .A2(n969), .ZN(n617) );
  INV_X1 U563 ( .A(n668), .ZN(n641) );
  INV_X1 U564 ( .A(KEYINPUT30), .ZN(n651) );
  INV_X1 U565 ( .A(G168), .ZN(n653) );
  AND2_X1 U566 ( .A1(n654), .A2(n653), .ZN(n657) );
  INV_X1 U567 ( .A(KEYINPUT102), .ZN(n647) );
  NAND2_X1 U568 ( .A1(G8), .A2(n668), .ZN(n703) );
  NOR2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n525) );
  NOR2_X1 U570 ( .A1(n602), .A2(n601), .ZN(n604) );
  INV_X1 U571 ( .A(G2105), .ZN(n526) );
  AND2_X1 U572 ( .A1(G2104), .A2(G2105), .ZN(n873) );
  NAND2_X1 U573 ( .A1(G114), .A2(n873), .ZN(n524) );
  NOR2_X1 U574 ( .A1(G2104), .A2(n526), .ZN(n874) );
  NAND2_X1 U575 ( .A1(G126), .A2(n874), .ZN(n523) );
  NAND2_X1 U576 ( .A1(n524), .A2(n523), .ZN(n530) );
  XOR2_X2 U577 ( .A(KEYINPUT17), .B(n525), .Z(n877) );
  NAND2_X1 U578 ( .A1(G138), .A2(n877), .ZN(n528) );
  NAND2_X1 U579 ( .A1(G102), .A2(n878), .ZN(n527) );
  NAND2_X1 U580 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U581 ( .A1(n530), .A2(n529), .ZN(G164) );
  XOR2_X1 U582 ( .A(G543), .B(KEYINPUT0), .Z(n547) );
  NAND2_X1 U583 ( .A1(n789), .A2(G51), .ZN(n531) );
  XOR2_X1 U584 ( .A(KEYINPUT75), .B(n531), .Z(n534) );
  INV_X1 U585 ( .A(G651), .ZN(n536) );
  NOR2_X1 U586 ( .A1(G543), .A2(n536), .ZN(n532) );
  NAND2_X1 U587 ( .A1(n790), .A2(G63), .ZN(n533) );
  NAND2_X1 U588 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U589 ( .A(KEYINPUT6), .B(n535), .ZN(n543) );
  NOR2_X1 U590 ( .A1(n547), .A2(n536), .ZN(n786) );
  NAND2_X1 U591 ( .A1(n786), .A2(G76), .ZN(n537) );
  XNOR2_X1 U592 ( .A(KEYINPUT74), .B(n537), .ZN(n540) );
  NOR2_X1 U593 ( .A1(G543), .A2(G651), .ZN(n785) );
  NAND2_X1 U594 ( .A1(n785), .A2(G89), .ZN(n538) );
  XNOR2_X1 U595 ( .A(KEYINPUT4), .B(n538), .ZN(n539) );
  NAND2_X1 U596 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U597 ( .A(n541), .B(KEYINPUT5), .Z(n542) );
  NOR2_X1 U598 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U599 ( .A(KEYINPUT76), .B(n544), .Z(n545) );
  XNOR2_X1 U600 ( .A(KEYINPUT7), .B(n545), .ZN(G168) );
  NAND2_X1 U601 ( .A1(G49), .A2(n789), .ZN(n546) );
  XNOR2_X1 U602 ( .A(n546), .B(KEYINPUT84), .ZN(n552) );
  NAND2_X1 U603 ( .A1(G87), .A2(n547), .ZN(n549) );
  NAND2_X1 U604 ( .A1(G74), .A2(G651), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U606 ( .A1(n790), .A2(n550), .ZN(n551) );
  NAND2_X1 U607 ( .A1(n552), .A2(n551), .ZN(G288) );
  NAND2_X1 U608 ( .A1(n786), .A2(G77), .ZN(n553) );
  XOR2_X1 U609 ( .A(KEYINPUT67), .B(n553), .Z(n555) );
  NAND2_X1 U610 ( .A1(n785), .A2(G90), .ZN(n554) );
  NAND2_X1 U611 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U612 ( .A(KEYINPUT9), .B(n556), .ZN(n560) );
  NAND2_X1 U613 ( .A1(n789), .A2(G52), .ZN(n558) );
  NAND2_X1 U614 ( .A1(G64), .A2(n790), .ZN(n557) );
  AND2_X1 U615 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U616 ( .A1(n560), .A2(n559), .ZN(G301) );
  INV_X1 U617 ( .A(G301), .ZN(G171) );
  NAND2_X1 U618 ( .A1(G88), .A2(n785), .ZN(n562) );
  NAND2_X1 U619 ( .A1(G62), .A2(n790), .ZN(n561) );
  NAND2_X1 U620 ( .A1(n562), .A2(n561), .ZN(n565) );
  NAND2_X1 U621 ( .A1(G75), .A2(n786), .ZN(n563) );
  XNOR2_X1 U622 ( .A(KEYINPUT85), .B(n563), .ZN(n564) );
  NOR2_X1 U623 ( .A1(n565), .A2(n564), .ZN(n567) );
  NAND2_X1 U624 ( .A1(n789), .A2(G50), .ZN(n566) );
  NAND2_X1 U625 ( .A1(n567), .A2(n566), .ZN(G303) );
  INV_X1 U626 ( .A(G303), .ZN(G166) );
  XOR2_X1 U627 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U628 ( .A1(G86), .A2(n785), .ZN(n569) );
  NAND2_X1 U629 ( .A1(G61), .A2(n790), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n569), .A2(n568), .ZN(n572) );
  NAND2_X1 U631 ( .A1(n786), .A2(G73), .ZN(n570) );
  XOR2_X1 U632 ( .A(KEYINPUT2), .B(n570), .Z(n571) );
  NOR2_X1 U633 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U634 ( .A1(n789), .A2(G48), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n574), .A2(n573), .ZN(G305) );
  NAND2_X1 U636 ( .A1(G85), .A2(n785), .ZN(n576) );
  NAND2_X1 U637 ( .A1(G72), .A2(n786), .ZN(n575) );
  NAND2_X1 U638 ( .A1(n576), .A2(n575), .ZN(n580) );
  NAND2_X1 U639 ( .A1(G47), .A2(n789), .ZN(n578) );
  NAND2_X1 U640 ( .A1(G60), .A2(n790), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n578), .A2(n577), .ZN(n579) );
  OR2_X1 U642 ( .A1(n580), .A2(n579), .ZN(G290) );
  NAND2_X1 U643 ( .A1(G101), .A2(n878), .ZN(n581) );
  XOR2_X1 U644 ( .A(n581), .B(KEYINPUT23), .Z(n583) );
  NAND2_X1 U645 ( .A1(n874), .A2(G125), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U647 ( .A1(G113), .A2(n873), .ZN(n584) );
  XNOR2_X1 U648 ( .A(KEYINPUT65), .B(n584), .ZN(n585) );
  NOR2_X1 U649 ( .A1(n586), .A2(n585), .ZN(n757) );
  AND2_X1 U650 ( .A1(G40), .A2(n757), .ZN(n588) );
  NAND2_X1 U651 ( .A1(G137), .A2(n877), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n587), .B(KEYINPUT66), .ZN(n758) );
  NAND2_X1 U653 ( .A1(n588), .A2(n758), .ZN(n709) );
  INV_X1 U654 ( .A(n709), .ZN(n589) );
  NOR2_X1 U655 ( .A1(G164), .A2(G1384), .ZN(n710) );
  NAND2_X1 U656 ( .A1(n589), .A2(n710), .ZN(n668) );
  INV_X1 U657 ( .A(n703), .ZN(n590) );
  NOR2_X1 U658 ( .A1(G1976), .A2(G288), .ZN(n684) );
  NAND2_X1 U659 ( .A1(n590), .A2(n684), .ZN(n591) );
  AND2_X1 U660 ( .A1(KEYINPUT33), .A2(n591), .ZN(n691) );
  NAND2_X1 U661 ( .A1(n641), .A2(G1996), .ZN(n593) );
  XNOR2_X1 U662 ( .A(KEYINPUT26), .B(KEYINPUT100), .ZN(n592) );
  XNOR2_X1 U663 ( .A(n593), .B(n592), .ZN(n607) );
  AND2_X1 U664 ( .A1(n668), .A2(G1341), .ZN(n605) );
  NAND2_X1 U665 ( .A1(n785), .A2(G81), .ZN(n594) );
  XNOR2_X1 U666 ( .A(n594), .B(KEYINPUT12), .ZN(n596) );
  NAND2_X1 U667 ( .A1(G68), .A2(n786), .ZN(n595) );
  NAND2_X1 U668 ( .A1(n596), .A2(n595), .ZN(n598) );
  XOR2_X1 U669 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n597) );
  XNOR2_X1 U670 ( .A(n598), .B(n597), .ZN(n602) );
  NAND2_X1 U671 ( .A1(G56), .A2(n790), .ZN(n599) );
  XNOR2_X1 U672 ( .A(n599), .B(KEYINPUT69), .ZN(n600) );
  XNOR2_X1 U673 ( .A(KEYINPUT14), .B(n600), .ZN(n601) );
  NAND2_X1 U674 ( .A1(n789), .A2(G43), .ZN(n603) );
  NAND2_X1 U675 ( .A1(n604), .A2(n603), .ZN(n977) );
  NOR2_X1 U676 ( .A1(n605), .A2(n977), .ZN(n606) );
  AND2_X1 U677 ( .A1(n607), .A2(n606), .ZN(n618) );
  NAND2_X1 U678 ( .A1(G66), .A2(n790), .ZN(n614) );
  NAND2_X1 U679 ( .A1(G79), .A2(n786), .ZN(n609) );
  NAND2_X1 U680 ( .A1(G54), .A2(n789), .ZN(n608) );
  NAND2_X1 U681 ( .A1(n609), .A2(n608), .ZN(n612) );
  NAND2_X1 U682 ( .A1(G92), .A2(n785), .ZN(n610) );
  XNOR2_X1 U683 ( .A(KEYINPUT71), .B(n610), .ZN(n611) );
  NOR2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U685 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U686 ( .A(n615), .B(KEYINPUT15), .ZN(n616) );
  XNOR2_X1 U687 ( .A(KEYINPUT72), .B(n616), .ZN(n969) );
  XNOR2_X1 U688 ( .A(n617), .B(KEYINPUT101), .ZN(n624) );
  NAND2_X1 U689 ( .A1(n618), .A2(n969), .ZN(n622) );
  NOR2_X1 U690 ( .A1(G2067), .A2(n668), .ZN(n620) );
  NOR2_X1 U691 ( .A1(n641), .A2(G1348), .ZN(n619) );
  NOR2_X1 U692 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U693 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U694 ( .A1(n624), .A2(n623), .ZN(n635) );
  NAND2_X1 U695 ( .A1(G53), .A2(n789), .ZN(n626) );
  NAND2_X1 U696 ( .A1(G65), .A2(n790), .ZN(n625) );
  NAND2_X1 U697 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U698 ( .A1(G91), .A2(n785), .ZN(n628) );
  NAND2_X1 U699 ( .A1(G78), .A2(n786), .ZN(n627) );
  NAND2_X1 U700 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U701 ( .A1(n630), .A2(n629), .ZN(n978) );
  NAND2_X1 U702 ( .A1(n641), .A2(G2072), .ZN(n631) );
  XNOR2_X1 U703 ( .A(n631), .B(KEYINPUT27), .ZN(n633) );
  AND2_X1 U704 ( .A1(G1956), .A2(n668), .ZN(n632) );
  NOR2_X1 U705 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U706 ( .A1(n978), .A2(n636), .ZN(n634) );
  NAND2_X1 U707 ( .A1(n635), .A2(n634), .ZN(n639) );
  NOR2_X1 U708 ( .A1(n978), .A2(n636), .ZN(n637) );
  XOR2_X1 U709 ( .A(n637), .B(KEYINPUT28), .Z(n638) );
  NAND2_X1 U710 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U711 ( .A(n640), .B(KEYINPUT29), .ZN(n646) );
  XOR2_X1 U712 ( .A(G2078), .B(KEYINPUT25), .Z(n923) );
  NOR2_X1 U713 ( .A1(n923), .A2(n668), .ZN(n643) );
  NOR2_X1 U714 ( .A1(n641), .A2(G1961), .ZN(n642) );
  NOR2_X1 U715 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U716 ( .A(KEYINPUT99), .B(n644), .ZN(n655) );
  AND2_X1 U717 ( .A1(G171), .A2(n655), .ZN(n645) );
  NOR2_X1 U718 ( .A1(n646), .A2(n645), .ZN(n648) );
  XNOR2_X1 U719 ( .A(n648), .B(n647), .ZN(n675) );
  NOR2_X1 U720 ( .A1(G1966), .A2(n703), .ZN(n660) );
  NOR2_X1 U721 ( .A1(G2084), .A2(n668), .ZN(n659) );
  NOR2_X1 U722 ( .A1(n660), .A2(n659), .ZN(n649) );
  XOR2_X1 U723 ( .A(KEYINPUT103), .B(n649), .Z(n650) );
  NAND2_X1 U724 ( .A1(G8), .A2(n650), .ZN(n652) );
  XNOR2_X1 U725 ( .A(n652), .B(n651), .ZN(n654) );
  NOR2_X1 U726 ( .A1(G171), .A2(n655), .ZN(n656) );
  NOR2_X1 U727 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U728 ( .A(KEYINPUT31), .B(n658), .Z(n674) );
  AND2_X1 U729 ( .A1(n675), .A2(n674), .ZN(n663) );
  AND2_X1 U730 ( .A1(G8), .A2(n659), .ZN(n661) );
  OR2_X1 U731 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U732 ( .A1(G1976), .A2(G288), .ZN(n981) );
  INV_X1 U733 ( .A(n981), .ZN(n664) );
  OR2_X1 U734 ( .A1(n703), .A2(n664), .ZN(n686) );
  INV_X1 U735 ( .A(n686), .ZN(n665) );
  AND2_X1 U736 ( .A1(n698), .A2(n665), .ZN(n682) );
  INV_X1 U737 ( .A(G8), .ZN(n673) );
  NOR2_X1 U738 ( .A1(G1971), .A2(n703), .ZN(n666) );
  XNOR2_X1 U739 ( .A(n666), .B(KEYINPUT104), .ZN(n667) );
  NOR2_X1 U740 ( .A1(G166), .A2(n667), .ZN(n671) );
  NOR2_X1 U741 ( .A1(G2090), .A2(n668), .ZN(n669) );
  XNOR2_X1 U742 ( .A(n669), .B(KEYINPUT105), .ZN(n670) );
  NAND2_X1 U743 ( .A1(n671), .A2(n670), .ZN(n672) );
  OR2_X1 U744 ( .A1(n673), .A2(n672), .ZN(n677) );
  AND2_X1 U745 ( .A1(n674), .A2(n677), .ZN(n676) );
  NAND2_X1 U746 ( .A1(n676), .A2(n675), .ZN(n680) );
  INV_X1 U747 ( .A(n677), .ZN(n678) );
  OR2_X1 U748 ( .A1(n678), .A2(G286), .ZN(n679) );
  NAND2_X1 U749 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U750 ( .A(n681), .B(KEYINPUT32), .ZN(n697) );
  NAND2_X1 U751 ( .A1(n682), .A2(n697), .ZN(n688) );
  NOR2_X1 U752 ( .A1(G1971), .A2(G303), .ZN(n683) );
  NOR2_X1 U753 ( .A1(n684), .A2(n683), .ZN(n982) );
  XNOR2_X1 U754 ( .A(KEYINPUT106), .B(n982), .ZN(n685) );
  OR2_X1 U755 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U756 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U757 ( .A1(KEYINPUT33), .A2(n519), .ZN(n690) );
  NOR2_X1 U758 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U759 ( .A(n692), .B(KEYINPUT107), .ZN(n693) );
  XOR2_X1 U760 ( .A(G1981), .B(G305), .Z(n974) );
  NAND2_X1 U761 ( .A1(n693), .A2(n974), .ZN(n708) );
  NOR2_X1 U762 ( .A1(G1981), .A2(G305), .ZN(n694) );
  XOR2_X1 U763 ( .A(n694), .B(KEYINPUT24), .Z(n695) );
  XNOR2_X1 U764 ( .A(KEYINPUT98), .B(n695), .ZN(n696) );
  OR2_X1 U765 ( .A1(n703), .A2(n696), .ZN(n706) );
  NAND2_X1 U766 ( .A1(n698), .A2(n697), .ZN(n701) );
  NOR2_X1 U767 ( .A1(G2090), .A2(G303), .ZN(n699) );
  NAND2_X1 U768 ( .A1(G8), .A2(n699), .ZN(n700) );
  NAND2_X1 U769 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U770 ( .A(n702), .B(KEYINPUT108), .ZN(n704) );
  NAND2_X1 U771 ( .A1(n704), .A2(n703), .ZN(n705) );
  AND2_X1 U772 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U773 ( .A1(n710), .A2(n709), .ZN(n752) );
  XNOR2_X1 U774 ( .A(KEYINPUT96), .B(n752), .ZN(n728) );
  NAND2_X1 U775 ( .A1(G105), .A2(n878), .ZN(n711) );
  XNOR2_X1 U776 ( .A(n711), .B(KEYINPUT38), .ZN(n718) );
  NAND2_X1 U777 ( .A1(G117), .A2(n873), .ZN(n713) );
  NAND2_X1 U778 ( .A1(G129), .A2(n874), .ZN(n712) );
  NAND2_X1 U779 ( .A1(n713), .A2(n712), .ZN(n716) );
  NAND2_X1 U780 ( .A1(G141), .A2(n877), .ZN(n714) );
  XNOR2_X1 U781 ( .A(KEYINPUT95), .B(n714), .ZN(n715) );
  NOR2_X1 U782 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U783 ( .A1(n718), .A2(n717), .ZN(n888) );
  NAND2_X1 U784 ( .A1(G1996), .A2(n888), .ZN(n727) );
  NAND2_X1 U785 ( .A1(G95), .A2(n878), .ZN(n720) );
  NAND2_X1 U786 ( .A1(G107), .A2(n873), .ZN(n719) );
  NAND2_X1 U787 ( .A1(n720), .A2(n719), .ZN(n723) );
  NAND2_X1 U788 ( .A1(n874), .A2(G119), .ZN(n721) );
  XOR2_X1 U789 ( .A(KEYINPUT94), .B(n721), .Z(n722) );
  NOR2_X1 U790 ( .A1(n723), .A2(n722), .ZN(n725) );
  NAND2_X1 U791 ( .A1(n877), .A2(G131), .ZN(n724) );
  NAND2_X1 U792 ( .A1(n725), .A2(n724), .ZN(n891) );
  NAND2_X1 U793 ( .A1(G1991), .A2(n891), .ZN(n726) );
  NAND2_X1 U794 ( .A1(n727), .A2(n726), .ZN(n961) );
  NAND2_X1 U795 ( .A1(n728), .A2(n961), .ZN(n744) );
  XOR2_X1 U796 ( .A(G2067), .B(KEYINPUT37), .Z(n729) );
  XNOR2_X1 U797 ( .A(KEYINPUT93), .B(n729), .ZN(n750) );
  NAND2_X1 U798 ( .A1(G140), .A2(n877), .ZN(n731) );
  NAND2_X1 U799 ( .A1(G104), .A2(n878), .ZN(n730) );
  NAND2_X1 U800 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U801 ( .A(KEYINPUT34), .B(n732), .ZN(n737) );
  NAND2_X1 U802 ( .A1(G116), .A2(n873), .ZN(n734) );
  NAND2_X1 U803 ( .A1(G128), .A2(n874), .ZN(n733) );
  NAND2_X1 U804 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U805 ( .A(KEYINPUT35), .B(n735), .Z(n736) );
  NOR2_X1 U806 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U807 ( .A(KEYINPUT36), .B(n738), .ZN(n887) );
  NOR2_X1 U808 ( .A1(n750), .A2(n887), .ZN(n940) );
  NAND2_X1 U809 ( .A1(n752), .A2(n940), .ZN(n749) );
  NAND2_X1 U810 ( .A1(n744), .A2(n749), .ZN(n739) );
  XNOR2_X1 U811 ( .A(n739), .B(KEYINPUT97), .ZN(n741) );
  XNOR2_X1 U812 ( .A(G1986), .B(G290), .ZN(n973) );
  NAND2_X1 U813 ( .A1(n752), .A2(n973), .ZN(n740) );
  NAND2_X1 U814 ( .A1(n522), .A2(n521), .ZN(n755) );
  NOR2_X1 U815 ( .A1(G1986), .A2(G290), .ZN(n742) );
  NOR2_X1 U816 ( .A1(G1991), .A2(n891), .ZN(n956) );
  NOR2_X1 U817 ( .A1(n742), .A2(n956), .ZN(n743) );
  XNOR2_X1 U818 ( .A(n743), .B(KEYINPUT109), .ZN(n745) );
  NAND2_X1 U819 ( .A1(n745), .A2(n744), .ZN(n746) );
  OR2_X1 U820 ( .A1(n888), .A2(G1996), .ZN(n943) );
  NAND2_X1 U821 ( .A1(n746), .A2(n943), .ZN(n747) );
  XOR2_X1 U822 ( .A(KEYINPUT39), .B(n747), .Z(n748) );
  NAND2_X1 U823 ( .A1(n749), .A2(n748), .ZN(n751) );
  NAND2_X1 U824 ( .A1(n750), .A2(n887), .ZN(n941) );
  NAND2_X1 U825 ( .A1(n751), .A2(n941), .ZN(n753) );
  NAND2_X1 U826 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U827 ( .A1(n755), .A2(n520), .ZN(n756) );
  XNOR2_X1 U828 ( .A(n756), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U829 ( .A1(n758), .A2(n757), .ZN(G160) );
  INV_X1 U830 ( .A(G57), .ZN(G237) );
  NAND2_X1 U831 ( .A1(G94), .A2(G452), .ZN(n759) );
  XOR2_X1 U832 ( .A(KEYINPUT68), .B(n759), .Z(G173) );
  NAND2_X1 U833 ( .A1(G7), .A2(G661), .ZN(n760) );
  XNOR2_X1 U834 ( .A(n760), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U835 ( .A(G223), .ZN(n831) );
  NAND2_X1 U836 ( .A1(n831), .A2(G567), .ZN(n761) );
  XOR2_X1 U837 ( .A(KEYINPUT11), .B(n761), .Z(G234) );
  INV_X1 U838 ( .A(G860), .ZN(n797) );
  OR2_X1 U839 ( .A1(n977), .A2(n797), .ZN(G153) );
  NOR2_X1 U840 ( .A1(G868), .A2(n969), .ZN(n763) );
  INV_X1 U841 ( .A(G868), .ZN(n809) );
  NOR2_X1 U842 ( .A1(G171), .A2(n809), .ZN(n762) );
  NOR2_X1 U843 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U844 ( .A(KEYINPUT73), .B(n764), .ZN(G284) );
  INV_X1 U845 ( .A(n978), .ZN(G299) );
  NOR2_X1 U846 ( .A1(G286), .A2(n809), .ZN(n765) );
  XOR2_X1 U847 ( .A(KEYINPUT77), .B(n765), .Z(n768) );
  NOR2_X1 U848 ( .A1(G868), .A2(G299), .ZN(n766) );
  XNOR2_X1 U849 ( .A(KEYINPUT78), .B(n766), .ZN(n767) );
  NOR2_X1 U850 ( .A1(n768), .A2(n767), .ZN(G297) );
  NAND2_X1 U851 ( .A1(n797), .A2(G559), .ZN(n769) );
  NAND2_X1 U852 ( .A1(n769), .A2(n969), .ZN(n770) );
  XNOR2_X1 U853 ( .A(n770), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U854 ( .A1(G868), .A2(n977), .ZN(n773) );
  NAND2_X1 U855 ( .A1(n969), .A2(G868), .ZN(n771) );
  NOR2_X1 U856 ( .A1(G559), .A2(n771), .ZN(n772) );
  NOR2_X1 U857 ( .A1(n773), .A2(n772), .ZN(G282) );
  NAND2_X1 U858 ( .A1(G99), .A2(n878), .ZN(n775) );
  NAND2_X1 U859 ( .A1(G111), .A2(n873), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U861 ( .A(n776), .B(KEYINPUT79), .ZN(n778) );
  NAND2_X1 U862 ( .A1(G135), .A2(n877), .ZN(n777) );
  NAND2_X1 U863 ( .A1(n778), .A2(n777), .ZN(n781) );
  NAND2_X1 U864 ( .A1(n874), .A2(G123), .ZN(n779) );
  XOR2_X1 U865 ( .A(KEYINPUT18), .B(n779), .Z(n780) );
  NOR2_X1 U866 ( .A1(n781), .A2(n780), .ZN(n955) );
  XOR2_X1 U867 ( .A(n955), .B(G2096), .Z(n782) );
  XNOR2_X1 U868 ( .A(KEYINPUT80), .B(n782), .ZN(n783) );
  NOR2_X1 U869 ( .A1(G2100), .A2(n783), .ZN(n784) );
  XNOR2_X1 U870 ( .A(KEYINPUT81), .B(n784), .ZN(G156) );
  NAND2_X1 U871 ( .A1(G93), .A2(n785), .ZN(n788) );
  NAND2_X1 U872 ( .A1(G80), .A2(n786), .ZN(n787) );
  NAND2_X1 U873 ( .A1(n788), .A2(n787), .ZN(n795) );
  NAND2_X1 U874 ( .A1(G55), .A2(n789), .ZN(n792) );
  NAND2_X1 U875 ( .A1(G67), .A2(n790), .ZN(n791) );
  NAND2_X1 U876 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U877 ( .A(KEYINPUT83), .B(n793), .Z(n794) );
  NOR2_X1 U878 ( .A1(n795), .A2(n794), .ZN(n808) );
  XOR2_X1 U879 ( .A(n808), .B(KEYINPUT82), .Z(n799) );
  NAND2_X1 U880 ( .A1(n969), .A2(G559), .ZN(n796) );
  XOR2_X1 U881 ( .A(n977), .B(n796), .Z(n806) );
  NAND2_X1 U882 ( .A1(n806), .A2(n797), .ZN(n798) );
  XNOR2_X1 U883 ( .A(n799), .B(n798), .ZN(G145) );
  XNOR2_X1 U884 ( .A(n978), .B(G288), .ZN(n805) );
  XNOR2_X1 U885 ( .A(KEYINPUT19), .B(KEYINPUT86), .ZN(n801) );
  XNOR2_X1 U886 ( .A(G290), .B(n808), .ZN(n800) );
  XNOR2_X1 U887 ( .A(n801), .B(n800), .ZN(n802) );
  XNOR2_X1 U888 ( .A(G166), .B(n802), .ZN(n803) );
  XNOR2_X1 U889 ( .A(n803), .B(G305), .ZN(n804) );
  XNOR2_X1 U890 ( .A(n805), .B(n804), .ZN(n899) );
  XNOR2_X1 U891 ( .A(n806), .B(n899), .ZN(n807) );
  NAND2_X1 U892 ( .A1(n807), .A2(G868), .ZN(n811) );
  NAND2_X1 U893 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U894 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U895 ( .A(KEYINPUT87), .B(n812), .ZN(G295) );
  NAND2_X1 U896 ( .A1(G2084), .A2(G2078), .ZN(n813) );
  XOR2_X1 U897 ( .A(KEYINPUT20), .B(n813), .Z(n814) );
  NAND2_X1 U898 ( .A1(G2090), .A2(n814), .ZN(n815) );
  XNOR2_X1 U899 ( .A(n815), .B(KEYINPUT89), .ZN(n817) );
  XOR2_X1 U900 ( .A(KEYINPUT21), .B(KEYINPUT88), .Z(n816) );
  XNOR2_X1 U901 ( .A(n817), .B(n816), .ZN(n818) );
  NAND2_X1 U902 ( .A1(n818), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U903 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U904 ( .A1(G132), .A2(G82), .ZN(n819) );
  XNOR2_X1 U905 ( .A(n819), .B(KEYINPUT22), .ZN(n820) );
  XNOR2_X1 U906 ( .A(n820), .B(KEYINPUT90), .ZN(n821) );
  NOR2_X1 U907 ( .A1(G218), .A2(n821), .ZN(n822) );
  NAND2_X1 U908 ( .A1(G96), .A2(n822), .ZN(n839) );
  NAND2_X1 U909 ( .A1(G2106), .A2(n839), .ZN(n823) );
  XNOR2_X1 U910 ( .A(KEYINPUT91), .B(n823), .ZN(n828) );
  NAND2_X1 U911 ( .A1(G120), .A2(G108), .ZN(n824) );
  NOR2_X1 U912 ( .A1(G237), .A2(n824), .ZN(n825) );
  NAND2_X1 U913 ( .A1(G69), .A2(n825), .ZN(n838) );
  NAND2_X1 U914 ( .A1(G567), .A2(n838), .ZN(n826) );
  XOR2_X1 U915 ( .A(KEYINPUT92), .B(n826), .Z(n827) );
  NOR2_X1 U916 ( .A1(n828), .A2(n827), .ZN(G319) );
  INV_X1 U917 ( .A(G319), .ZN(n830) );
  NAND2_X1 U918 ( .A1(G661), .A2(G483), .ZN(n829) );
  NOR2_X1 U919 ( .A1(n830), .A2(n829), .ZN(n837) );
  NAND2_X1 U920 ( .A1(n837), .A2(G36), .ZN(G176) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n831), .ZN(G217) );
  INV_X1 U922 ( .A(G661), .ZN(n833) );
  NAND2_X1 U923 ( .A1(G2), .A2(G15), .ZN(n832) );
  NOR2_X1 U924 ( .A1(n833), .A2(n832), .ZN(n834) );
  XOR2_X1 U925 ( .A(KEYINPUT112), .B(n834), .Z(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n835) );
  XOR2_X1 U927 ( .A(KEYINPUT113), .B(n835), .Z(n836) );
  NAND2_X1 U928 ( .A1(n837), .A2(n836), .ZN(G188) );
  XNOR2_X1 U929 ( .A(G108), .B(KEYINPUT117), .ZN(G238) );
  INV_X1 U931 ( .A(G132), .ZN(G219) );
  INV_X1 U932 ( .A(G120), .ZN(G236) );
  INV_X1 U933 ( .A(G82), .ZN(G220) );
  NOR2_X1 U934 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U935 ( .A(G325), .ZN(G261) );
  XOR2_X1 U936 ( .A(KEYINPUT43), .B(KEYINPUT42), .Z(n841) );
  XNOR2_X1 U937 ( .A(G2678), .B(KEYINPUT115), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U939 ( .A(KEYINPUT114), .B(G2090), .Z(n843) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2072), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U942 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U943 ( .A(G2096), .B(G2100), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(n849) );
  XOR2_X1 U945 ( .A(G2084), .B(G2078), .Z(n848) );
  XNOR2_X1 U946 ( .A(n849), .B(n848), .ZN(G227) );
  XOR2_X1 U947 ( .A(G1986), .B(G1976), .Z(n851) );
  XNOR2_X1 U948 ( .A(G1961), .B(G1971), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U950 ( .A(n852), .B(G2474), .Z(n854) );
  XNOR2_X1 U951 ( .A(G1966), .B(G1981), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U953 ( .A(KEYINPUT41), .B(G1991), .Z(n856) );
  XNOR2_X1 U954 ( .A(G1996), .B(G1956), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n858), .B(n857), .ZN(G229) );
  NAND2_X1 U957 ( .A1(G124), .A2(n874), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n859), .B(KEYINPUT44), .ZN(n861) );
  NAND2_X1 U959 ( .A1(n878), .A2(G100), .ZN(n860) );
  NAND2_X1 U960 ( .A1(n861), .A2(n860), .ZN(n865) );
  NAND2_X1 U961 ( .A1(G136), .A2(n877), .ZN(n863) );
  NAND2_X1 U962 ( .A1(G112), .A2(n873), .ZN(n862) );
  NAND2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n864) );
  NOR2_X1 U964 ( .A1(n865), .A2(n864), .ZN(G162) );
  NAND2_X1 U965 ( .A1(G139), .A2(n877), .ZN(n867) );
  NAND2_X1 U966 ( .A1(G103), .A2(n878), .ZN(n866) );
  NAND2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n872) );
  NAND2_X1 U968 ( .A1(G115), .A2(n873), .ZN(n869) );
  NAND2_X1 U969 ( .A1(G127), .A2(n874), .ZN(n868) );
  NAND2_X1 U970 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U971 ( .A(KEYINPUT47), .B(n870), .Z(n871) );
  NOR2_X1 U972 ( .A1(n872), .A2(n871), .ZN(n947) );
  XNOR2_X1 U973 ( .A(n947), .B(n955), .ZN(n885) );
  NAND2_X1 U974 ( .A1(G118), .A2(n873), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G130), .A2(n874), .ZN(n875) );
  NAND2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n883) );
  NAND2_X1 U977 ( .A1(G142), .A2(n877), .ZN(n880) );
  NAND2_X1 U978 ( .A1(G106), .A2(n878), .ZN(n879) );
  NAND2_X1 U979 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U980 ( .A(KEYINPUT45), .B(n881), .Z(n882) );
  NOR2_X1 U981 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U982 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U983 ( .A(n887), .B(n886), .ZN(n890) );
  XOR2_X1 U984 ( .A(G160), .B(n888), .Z(n889) );
  XNOR2_X1 U985 ( .A(n890), .B(n889), .ZN(n896) );
  XNOR2_X1 U986 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n893) );
  XNOR2_X1 U987 ( .A(n891), .B(G162), .ZN(n892) );
  XNOR2_X1 U988 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U989 ( .A(G164), .B(n894), .Z(n895) );
  XNOR2_X1 U990 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U991 ( .A1(G37), .A2(n897), .ZN(G395) );
  XOR2_X1 U992 ( .A(n969), .B(n977), .Z(n898) );
  XNOR2_X1 U993 ( .A(G286), .B(n898), .ZN(n901) );
  XOR2_X1 U994 ( .A(G301), .B(n899), .Z(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U996 ( .A1(G37), .A2(n902), .ZN(n903) );
  XNOR2_X1 U997 ( .A(KEYINPUT116), .B(n903), .ZN(G397) );
  XOR2_X1 U998 ( .A(G2430), .B(G2451), .Z(n905) );
  XNOR2_X1 U999 ( .A(G2446), .B(G2427), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(n905), .B(n904), .ZN(n912) );
  XOR2_X1 U1001 ( .A(G2438), .B(KEYINPUT111), .Z(n907) );
  XNOR2_X1 U1002 ( .A(G2443), .B(G2454), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1004 ( .A(n908), .B(G2435), .Z(n910) );
  XNOR2_X1 U1005 ( .A(G1348), .B(G1341), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1007 ( .A(n912), .B(n911), .ZN(n913) );
  NAND2_X1 U1008 ( .A1(n913), .A2(G14), .ZN(n919) );
  NAND2_X1 U1009 ( .A1(G319), .A2(n919), .ZN(n916) );
  NOR2_X1 U1010 ( .A1(G227), .A2(G229), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(KEYINPUT49), .B(n914), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1014 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(G69), .ZN(G235) );
  INV_X1 U1017 ( .A(G96), .ZN(G221) );
  INV_X1 U1018 ( .A(n919), .ZN(G401) );
  XOR2_X1 U1019 ( .A(G1991), .B(G25), .Z(n920) );
  NAND2_X1 U1020 ( .A1(n920), .A2(G28), .ZN(n929) );
  XNOR2_X1 U1021 ( .A(G1996), .B(G32), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(G33), .B(G2072), .ZN(n921) );
  NOR2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(n923), .B(G27), .ZN(n925) );
  XNOR2_X1 U1025 ( .A(G2067), .B(G26), .ZN(n924) );
  NOR2_X1 U1026 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1029 ( .A(KEYINPUT53), .B(n930), .Z(n933) );
  XOR2_X1 U1030 ( .A(KEYINPUT54), .B(G34), .Z(n931) );
  XNOR2_X1 U1031 ( .A(G2084), .B(n931), .ZN(n932) );
  NAND2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n935) );
  XNOR2_X1 U1033 ( .A(G35), .B(G2090), .ZN(n934) );
  NOR2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1035 ( .A1(n936), .A2(KEYINPUT55), .ZN(n1028) );
  INV_X1 U1036 ( .A(n936), .ZN(n938) );
  NOR2_X1 U1037 ( .A1(G29), .A2(KEYINPUT55), .ZN(n937) );
  NAND2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1039 ( .A1(G11), .A2(n939), .ZN(n1026) );
  INV_X1 U1040 ( .A(KEYINPUT55), .ZN(n967) );
  INV_X1 U1041 ( .A(n940), .ZN(n942) );
  NAND2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n954) );
  XNOR2_X1 U1043 ( .A(G2090), .B(G162), .ZN(n944) );
  NAND2_X1 U1044 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1045 ( .A(n945), .B(KEYINPUT119), .ZN(n946) );
  XOR2_X1 U1046 ( .A(KEYINPUT51), .B(n946), .Z(n952) );
  XOR2_X1 U1047 ( .A(G2072), .B(n947), .Z(n949) );
  XOR2_X1 U1048 ( .A(G164), .B(G2078), .Z(n948) );
  NOR2_X1 U1049 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1050 ( .A(KEYINPUT50), .B(n950), .ZN(n951) );
  NAND2_X1 U1051 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n963) );
  NOR2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1054 ( .A(KEYINPUT118), .B(n957), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(G160), .B(G2084), .ZN(n958) );
  NAND2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(KEYINPUT120), .B(n964), .ZN(n965) );
  XOR2_X1 U1060 ( .A(KEYINPUT52), .B(n965), .Z(n966) );
  NAND2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n968), .A2(G29), .ZN(n1024) );
  XNOR2_X1 U1063 ( .A(G16), .B(KEYINPUT56), .ZN(n993) );
  XNOR2_X1 U1064 ( .A(n969), .B(G1348), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(G303), .A2(G1971), .ZN(n970) );
  NAND2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n991) );
  XNOR2_X1 U1068 ( .A(G1966), .B(G168), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(KEYINPUT57), .B(n976), .ZN(n986) );
  XOR2_X1 U1071 ( .A(n977), .B(G1341), .Z(n980) );
  XNOR2_X1 U1072 ( .A(n978), .B(G1956), .ZN(n979) );
  NAND2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n984) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n989) );
  XOR2_X1 U1077 ( .A(G1961), .B(G301), .Z(n987) );
  XNOR2_X1 U1078 ( .A(KEYINPUT121), .B(n987), .ZN(n988) );
  NOR2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n1021) );
  INV_X1 U1082 ( .A(G16), .ZN(n1019) );
  XNOR2_X1 U1083 ( .A(KEYINPUT123), .B(G1341), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(n994), .B(G19), .ZN(n999) );
  XOR2_X1 U1085 ( .A(G1348), .B(KEYINPUT59), .Z(n995) );
  XNOR2_X1 U1086 ( .A(G4), .B(n995), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(G20), .B(G1956), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(KEYINPUT124), .B(G1981), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(G6), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(KEYINPUT60), .B(n1003), .ZN(n1014) );
  XNOR2_X1 U1094 ( .A(G1961), .B(KEYINPUT122), .ZN(n1004) );
  XNOR2_X1 U1095 ( .A(n1004), .B(G5), .ZN(n1012) );
  XNOR2_X1 U1096 ( .A(G1971), .B(G22), .ZN(n1006) );
  XNOR2_X1 U1097 ( .A(G23), .B(G1976), .ZN(n1005) );
  NOR2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(G1986), .B(KEYINPUT125), .ZN(n1007) );
  XNOR2_X1 U1100 ( .A(n1007), .B(G24), .ZN(n1008) );
  NAND2_X1 U1101 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1102 ( .A(KEYINPUT58), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  XNOR2_X1 U1105 ( .A(G21), .B(G1966), .ZN(n1015) );
  NOR2_X1 U1106 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1107 ( .A(KEYINPUT61), .B(n1017), .ZN(n1018) );
  NAND2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1110 ( .A(KEYINPUT126), .B(n1022), .Z(n1023) );
  NAND2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1114 ( .A(n1029), .B(KEYINPUT62), .ZN(n1030) );
  XNOR2_X1 U1115 ( .A(KEYINPUT127), .B(n1030), .ZN(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

