//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n796, new_n797, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934;
  XNOR2_X1  g000(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(G127gat), .B(G155gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G231gat), .ZN(new_n207));
  INV_X1    g006(.A(G233gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G15gat), .B(G22gat), .ZN(new_n210));
  INV_X1    g009(.A(G1gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT16), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(G1gat), .B2(new_n210), .ZN(new_n214));
  INV_X1    g013(.A(G8gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n214), .B(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT21), .ZN(new_n217));
  INV_X1    g016(.A(G57gat), .ZN(new_n218));
  OR3_X1    g017(.A1(new_n218), .A2(KEYINPUT92), .A3(G64gat), .ZN(new_n219));
  INV_X1    g018(.A(G64gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G57gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT92), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n218), .A2(G64gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n219), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G71gat), .A2(G78gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(G71gat), .A2(G78gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT9), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n225), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n224), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT91), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n223), .A2(new_n221), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n231), .B1(new_n223), .B2(new_n221), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n225), .A2(new_n228), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NOR3_X1   g034(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT90), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n227), .A2(new_n237), .A3(new_n225), .ZN(new_n238));
  INV_X1    g037(.A(new_n225), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT90), .B1(new_n239), .B2(new_n226), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n230), .B1(new_n236), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n216), .B1(new_n217), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G183gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n242), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n246), .A2(KEYINPUT21), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n243), .B(G183gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n247), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n209), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n249), .A2(new_n251), .A3(new_n209), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n206), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n249), .A2(new_n251), .A3(new_n209), .ZN(new_n256));
  NOR3_X1   g055(.A1(new_n256), .A2(new_n252), .A3(new_n205), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n203), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n253), .A2(new_n206), .A3(new_n254), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n205), .B1(new_n256), .B2(new_n252), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(new_n202), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT87), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT87), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n265), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT14), .ZN(new_n267));
  INV_X1    g066(.A(G29gat), .ZN(new_n268));
  INV_X1    g067(.A(G36gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n264), .A2(new_n266), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G29gat), .A2(G36gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G50gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n274), .A2(G43gat), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(G43gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(KEYINPUT15), .A3(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT17), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT88), .B(G43gat), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n275), .B1(new_n282), .B2(new_n274), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n272), .B1(new_n283), .B2(KEYINPUT15), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT89), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n267), .A2(new_n268), .A3(new_n269), .A4(KEYINPUT89), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(new_n287), .A3(new_n263), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(new_n278), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n280), .B(new_n281), .C1(new_n284), .C2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G43gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT88), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT88), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G43gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n295), .A3(new_n274), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(new_n276), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT15), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n299), .A2(new_n278), .A3(new_n272), .A4(new_n288), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n281), .B1(new_n300), .B2(new_n280), .ZN(new_n301));
  NAND2_X1  g100(.A1(G99gat), .A2(G106gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT8), .ZN(new_n303));
  NAND2_X1  g102(.A1(G85gat), .A2(G92gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT7), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G85gat), .ZN(new_n307));
  INV_X1    g106(.A(G92gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n303), .A2(new_n306), .A3(new_n309), .A4(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G99gat), .B(G106gat), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT93), .ZN(new_n315));
  AOI22_X1  g114(.A1(KEYINPUT8), .A2(new_n302), .B1(new_n307), .B2(new_n308), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n316), .A2(new_n312), .A3(new_n306), .A4(new_n310), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n314), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n311), .A2(KEYINPUT93), .A3(new_n313), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(KEYINPUT94), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT94), .B1(new_n318), .B2(new_n319), .ZN(new_n322));
  OAI22_X1  g121(.A1(new_n291), .A2(new_n301), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n318), .A2(new_n319), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT94), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n300), .A2(new_n280), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(new_n328), .A3(new_n320), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n323), .A2(new_n324), .A3(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G190gat), .B(G218gat), .ZN(new_n331));
  OR2_X1    g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n331), .ZN(new_n333));
  XOR2_X1   g132(.A(G134gat), .B(G162gat), .Z(new_n334));
  AOI21_X1  g133(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n332), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n336), .B1(new_n332), .B2(new_n333), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT84), .ZN(new_n340));
  XNOR2_X1  g139(.A(G155gat), .B(G162gat), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT2), .ZN(new_n342));
  INV_X1    g141(.A(G148gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G141gat), .ZN(new_n344));
  INV_X1    g143(.A(G141gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G148gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n341), .B1(new_n342), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT74), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n342), .B1(G155gat), .B2(G162gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(KEYINPUT77), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n344), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n343), .A2(KEYINPUT76), .A3(G141gat), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n346), .A2(KEYINPUT75), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n346), .A2(KEYINPUT75), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n354), .B(new_n355), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n352), .A2(new_n358), .A3(new_n341), .ZN(new_n359));
  XOR2_X1   g158(.A(G127gat), .B(G134gat), .Z(new_n360));
  INV_X1    g159(.A(G113gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(G120gat), .ZN(new_n362));
  INV_X1    g161(.A(G120gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(G113gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n360), .B1(new_n365), .B2(KEYINPUT1), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n360), .A2(KEYINPUT1), .ZN(new_n367));
  OR3_X1    g166(.A1(new_n361), .A2(KEYINPUT69), .A3(G120gat), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT69), .B1(new_n361), .B2(G120gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n367), .B1(new_n364), .B2(new_n370), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n350), .A2(new_n359), .A3(new_n366), .A4(new_n371), .ZN(new_n372));
  XOR2_X1   g171(.A(new_n372), .B(KEYINPUT4), .Z(new_n373));
  NAND2_X1  g172(.A1(new_n350), .A2(new_n359), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT3), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT78), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n374), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT79), .B1(new_n374), .B2(KEYINPUT3), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT79), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n350), .A2(new_n380), .A3(new_n381), .A4(new_n359), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n377), .A2(new_n378), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n371), .A2(new_n366), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n373), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G225gat), .A2(G233gat), .ZN(new_n386));
  XOR2_X1   g185(.A(new_n386), .B(KEYINPUT80), .Z(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n340), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n383), .A2(new_n384), .ZN(new_n390));
  INV_X1    g189(.A(new_n373), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n392), .A2(KEYINPUT84), .A3(new_n387), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT39), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G1gat), .B(G29gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(G85gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT0), .B(G57gat), .ZN(new_n399));
  XOR2_X1   g198(.A(new_n398), .B(new_n399), .Z(new_n400));
  AOI21_X1  g199(.A(new_n387), .B1(new_n374), .B2(new_n384), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n395), .B1(new_n401), .B2(new_n372), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n389), .A2(new_n393), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n396), .A2(new_n400), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT40), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n385), .A2(KEYINPUT5), .A3(new_n388), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT5), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n400), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n374), .A2(new_n384), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n411), .A2(KEYINPUT5), .A3(new_n372), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n387), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n407), .A2(new_n409), .A3(new_n410), .A4(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G197gat), .B(G204gat), .ZN(new_n415));
  INV_X1    g214(.A(G211gat), .ZN(new_n416));
  INV_X1    g215(.A(G218gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n415), .B1(KEYINPUT22), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G211gat), .B(G218gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(KEYINPUT27), .B(G183gat), .ZN(new_n423));
  INV_X1    g222(.A(G190gat), .ZN(new_n424));
  AND2_X1   g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n426));
  AOI22_X1  g225(.A1(new_n425), .A2(new_n426), .B1(G183gat), .B2(G190gat), .ZN(new_n427));
  NOR2_X1   g226(.A1(G169gat), .A2(G176gat), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT68), .ZN(new_n430));
  OR3_X1    g229(.A1(new_n429), .A2(new_n430), .A3(KEYINPUT26), .ZN(new_n431));
  INV_X1    g230(.A(G169gat), .ZN(new_n432));
  INV_X1    g231(.A(G176gat), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n429), .A2(KEYINPUT26), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n430), .B1(new_n429), .B2(KEYINPUT26), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n431), .A2(new_n435), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n427), .B(new_n438), .C1(new_n425), .C2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT23), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n441), .A2(G169gat), .A3(G176gat), .ZN(new_n442));
  OR3_X1    g241(.A1(new_n428), .A2(KEYINPUT66), .A3(KEYINPUT23), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT66), .B1(new_n428), .B2(KEYINPUT23), .ZN(new_n444));
  AOI211_X1 g243(.A(new_n442), .B(new_n434), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n244), .A2(new_n424), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n446), .B(KEYINPUT65), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT24), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n448), .B1(new_n244), .B2(new_n424), .ZN(new_n449));
  OR2_X1    g248(.A1(new_n449), .A2(KEYINPUT64), .ZN(new_n450));
  NAND3_X1  g249(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(KEYINPUT64), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n447), .A2(new_n450), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT25), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n445), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n449), .A2(new_n446), .A3(new_n451), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n445), .A2(new_n456), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n440), .B(new_n455), .C1(new_n457), .C2(new_n454), .ZN(new_n458));
  AND2_X1   g257(.A1(G226gat), .A2(G233gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT29), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n422), .B(new_n460), .C1(new_n462), .C2(new_n459), .ZN(new_n463));
  OR2_X1    g262(.A1(new_n463), .A2(KEYINPUT73), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n462), .A2(new_n459), .ZN(new_n465));
  INV_X1    g264(.A(new_n460), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n421), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n463), .A2(KEYINPUT73), .ZN(new_n468));
  XNOR2_X1  g267(.A(G8gat), .B(G36gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(G64gat), .B(G92gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n464), .A2(new_n467), .A3(new_n468), .A4(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT30), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n464), .A2(new_n467), .A3(new_n468), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n471), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n473), .A2(new_n474), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n475), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n396), .A2(KEYINPUT40), .A3(new_n400), .A4(new_n403), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n406), .A2(new_n414), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n381), .B1(new_n421), .B2(KEYINPUT29), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n374), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT29), .B1(new_n379), .B2(new_n382), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n483), .B1(new_n484), .B2(new_n422), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT81), .ZN(new_n486));
  NAND2_X1  g285(.A1(G228gat), .A2(G233gat), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT81), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n488), .B(new_n483), .C1(new_n484), .C2(new_n422), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n486), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n485), .A2(KEYINPUT81), .A3(G228gat), .A4(G233gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(G22gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n490), .A2(G22gat), .A3(new_n491), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT82), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n497), .B1(new_n492), .B2(new_n493), .ZN(new_n498));
  XOR2_X1   g297(.A(G78gat), .B(G106gat), .Z(new_n499));
  XNOR2_X1  g298(.A(new_n499), .B(KEYINPUT31), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(new_n274), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n496), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n494), .A2(new_n497), .A3(new_n495), .A4(new_n501), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT38), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT37), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n464), .A2(new_n507), .A3(new_n467), .A4(new_n468), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT86), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n508), .A2(new_n509), .ZN(new_n511));
  OR2_X1    g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n476), .A2(KEYINPUT37), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n506), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT85), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n463), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n516), .A2(new_n507), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n467), .A2(new_n515), .A3(new_n463), .ZN(new_n518));
  AOI211_X1 g317(.A(KEYINPUT38), .B(new_n472), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n519), .B1(new_n510), .B2(new_n511), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n407), .A2(new_n409), .A3(new_n413), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT6), .ZN(new_n522));
  OR3_X1    g321(.A1(new_n521), .A2(new_n522), .A3(new_n400), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n400), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n524), .A2(new_n522), .A3(new_n414), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n476), .A2(new_n506), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(new_n472), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n520), .A2(new_n523), .A3(new_n525), .A4(new_n527), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n481), .B(new_n505), .C1(new_n514), .C2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT83), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n505), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n479), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n525), .A2(new_n523), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n503), .A2(KEYINPUT83), .A3(new_n504), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G15gat), .B(G43gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(G71gat), .B(G99gat), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n537), .B(new_n538), .Z(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n458), .B(new_n384), .ZN(new_n541));
  NAND2_X1  g340(.A1(G227gat), .A2(G233gat), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT33), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n540), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(KEYINPUT32), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n547), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT70), .B1(new_n541), .B2(new_n543), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n551), .A2(KEYINPUT34), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n551), .A2(KEYINPUT34), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n548), .B(new_n549), .C1(new_n552), .C2(new_n553), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(KEYINPUT36), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n555), .A2(KEYINPUT72), .A3(new_n556), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n558), .B1(KEYINPUT72), .B2(new_n556), .ZN(new_n559));
  XNOR2_X1  g358(.A(KEYINPUT71), .B(KEYINPUT36), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n557), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n529), .A2(new_n536), .A3(new_n562), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n559), .A2(new_n505), .A3(new_n533), .A4(new_n532), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT35), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n555), .A2(new_n556), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n566), .B1(new_n503), .B2(new_n504), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n532), .A2(new_n533), .A3(KEYINPUT35), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n564), .A2(new_n565), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AOI211_X1 g368(.A(new_n262), .B(new_n339), .C1(new_n563), .C2(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n216), .B1(new_n291), .B2(new_n301), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n214), .B(G8gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(new_n328), .ZN(new_n573));
  NAND2_X1  g372(.A1(G229gat), .A2(G233gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT18), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n572), .B(new_n328), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n574), .B(KEYINPUT13), .Z(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n571), .A2(KEYINPUT18), .A3(new_n573), .A4(new_n574), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n577), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G113gat), .B(G141gat), .ZN(new_n583));
  INV_X1    g382(.A(G197gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT11), .B(G169gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT12), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n582), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n577), .A2(new_n580), .A3(new_n588), .A4(new_n581), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(G230gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n594), .A2(new_n208), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n223), .A2(new_n221), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT91), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n223), .A2(new_n221), .A3(new_n231), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(new_n234), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n238), .A2(new_n240), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(KEYINPUT10), .A3(new_n230), .ZN(new_n603));
  NOR3_X1   g402(.A1(new_n321), .A2(new_n322), .A3(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(KEYINPUT95), .B(KEYINPUT10), .Z(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n325), .A2(new_n242), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n314), .A2(new_n317), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n602), .A2(new_n608), .A3(new_n230), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n606), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n596), .B1(new_n604), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n607), .A2(new_n609), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n611), .B1(new_n596), .B2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G176gat), .B(G204gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(new_n343), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT96), .B(G120gat), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n615), .B(new_n616), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n613), .B(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n593), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n570), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n620), .A2(new_n533), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(new_n211), .ZN(G1324gat));
  NOR2_X1   g421(.A1(new_n620), .A2(new_n532), .ZN(new_n623));
  NAND2_X1  g422(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n624));
  OR2_X1    g423(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n626), .A2(KEYINPUT42), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(KEYINPUT42), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n627), .B(new_n628), .C1(new_n215), .C2(new_n623), .ZN(G1325gat));
  INV_X1    g428(.A(G15gat), .ZN(new_n630));
  INV_X1    g429(.A(new_n559), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n630), .B1(new_n620), .B2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT97), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n620), .A2(new_n630), .A3(new_n562), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(G1326gat));
  NAND2_X1  g434(.A1(new_n531), .A2(new_n535), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n620), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(KEYINPUT43), .B(G22gat), .Z(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(G1327gat));
  NAND2_X1  g438(.A1(new_n262), .A2(new_n619), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n563), .A2(new_n569), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n339), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n339), .B(KEYINPUT100), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT99), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n644), .B1(new_n645), .B2(KEYINPUT44), .ZN(new_n646));
  OAI21_X1  g445(.A(KEYINPUT44), .B1(new_n642), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n641), .A2(new_n645), .A3(new_n646), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n640), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(G29gat), .B1(new_n650), .B2(new_n533), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n642), .A2(new_n640), .ZN(new_n652));
  INV_X1    g451(.A(new_n533), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n652), .A2(new_n268), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g453(.A(KEYINPUT98), .B(KEYINPUT45), .Z(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n651), .A2(new_n656), .ZN(G1328gat));
  NAND3_X1  g456(.A1(new_n652), .A2(new_n269), .A3(new_n479), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n658), .B(KEYINPUT46), .Z(new_n659));
  OAI21_X1  g458(.A(G36gat), .B1(new_n650), .B2(new_n532), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(G1329gat));
  INV_X1    g460(.A(new_n562), .ZN(new_n662));
  INV_X1    g461(.A(new_n640), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664));
  INV_X1    g463(.A(new_n339), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n665), .B1(new_n563), .B2(new_n569), .ZN(new_n666));
  INV_X1    g465(.A(new_n646), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n664), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n648), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n662), .B(new_n663), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n631), .A2(new_n282), .ZN(new_n671));
  AOI22_X1  g470(.A1(new_n670), .A2(new_n282), .B1(new_n652), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT47), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(KEYINPUT101), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n673), .A2(KEYINPUT101), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1330gat));
  OAI21_X1  g476(.A(G50gat), .B1(new_n650), .B2(new_n505), .ZN(new_n678));
  NOR4_X1   g477(.A1(new_n642), .A2(G50gat), .A3(new_n636), .A4(new_n640), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n678), .A2(KEYINPUT48), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n636), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n649), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n679), .B1(new_n683), .B2(G50gat), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n681), .B1(KEYINPUT48), .B2(new_n684), .ZN(G1331gat));
  AND3_X1   g484(.A1(new_n570), .A2(new_n593), .A3(new_n618), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n653), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G57gat), .ZN(G1332gat));
  INV_X1    g487(.A(KEYINPUT49), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n686), .B(new_n479), .C1(new_n689), .C2(new_n220), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n220), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1333gat));
  AOI21_X1  g491(.A(G71gat), .B1(new_n686), .B2(new_n559), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n662), .A2(G71gat), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n693), .B1(new_n686), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT50), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1334gat));
  NAND2_X1  g496(.A1(new_n686), .A2(new_n682), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT102), .B(G78gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1335gat));
  AOI21_X1  g499(.A(KEYINPUT103), .B1(new_n641), .B2(new_n339), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n262), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n703), .A2(new_n592), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n666), .A2(KEYINPUT103), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n702), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT51), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT103), .ZN(new_n709));
  AOI211_X1 g508(.A(new_n709), .B(new_n665), .C1(new_n563), .C2(new_n569), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n701), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n711), .A2(KEYINPUT51), .A3(new_n704), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n713), .A2(new_n307), .A3(new_n653), .A4(new_n618), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n618), .B(new_n704), .C1(new_n668), .C2(new_n669), .ZN(new_n715));
  OAI21_X1  g514(.A(G85gat), .B1(new_n715), .B2(new_n533), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(G1336gat));
  NAND3_X1  g516(.A1(new_n479), .A2(new_n308), .A3(new_n618), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT105), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT51), .B1(new_n711), .B2(new_n704), .ZN(new_n720));
  INV_X1    g519(.A(new_n704), .ZN(new_n721));
  NOR4_X1   g520(.A1(new_n701), .A2(new_n710), .A3(new_n707), .A4(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n719), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G92gat), .B1(new_n715), .B2(new_n532), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n725), .A2(new_n727), .A3(KEYINPUT52), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT52), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n723), .B(new_n726), .C1(new_n724), .C2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(G1337gat));
  NOR2_X1   g530(.A1(new_n631), .A2(G99gat), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n713), .A2(new_n618), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G99gat), .B1(new_n715), .B2(new_n562), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(G1338gat));
  NOR2_X1   g534(.A1(new_n715), .A2(new_n636), .ZN(new_n736));
  INV_X1    g535(.A(G106gat), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n618), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n505), .A2(G106gat), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT106), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n741), .B1(new_n708), .B2(new_n712), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT53), .B1(new_n738), .B2(new_n742), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n742), .A2(KEYINPUT53), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT107), .B1(new_n715), .B2(new_n505), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n739), .B1(new_n647), .B2(new_n648), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT107), .ZN(new_n747));
  INV_X1    g546(.A(new_n505), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n746), .A2(new_n747), .A3(new_n748), .A4(new_n704), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n745), .A2(new_n749), .A3(G106gat), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n743), .B1(new_n744), .B2(new_n750), .ZN(G1339gat));
  AOI22_X1  g550(.A1(new_n602), .A2(new_n230), .B1(new_n318), .B2(new_n319), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n602), .A2(new_n608), .A3(new_n230), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n605), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n327), .A2(KEYINPUT10), .A3(new_n246), .A4(new_n320), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n754), .A2(new_n755), .A3(new_n595), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n611), .A2(KEYINPUT54), .A3(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n611), .A2(KEYINPUT108), .A3(new_n756), .A4(KEYINPUT54), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n617), .B1(new_n611), .B2(KEYINPUT54), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n613), .A2(new_n617), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n762), .B1(new_n759), .B2(new_n760), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n767), .B1(new_n768), .B2(KEYINPUT55), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n592), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n578), .A2(new_n579), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n574), .B1(new_n571), .B2(new_n573), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n587), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n591), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n618), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n643), .B1(new_n771), .B2(new_n776), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n643), .A2(new_n775), .A3(new_n770), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n262), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n258), .A2(new_n665), .A3(new_n739), .A4(new_n261), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n780), .A2(new_n592), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n783), .A2(new_n682), .A3(new_n631), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n533), .A2(new_n479), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(G113gat), .B1(new_n786), .B2(new_n593), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n782), .A2(new_n653), .A3(new_n567), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n532), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n592), .A2(new_n361), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n787), .B1(new_n789), .B2(new_n790), .ZN(G1340gat));
  OAI21_X1  g590(.A(G120gat), .B1(new_n786), .B2(new_n739), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n479), .A2(new_n739), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n788), .A2(new_n363), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(G1341gat));
  OAI21_X1  g594(.A(G127gat), .B1(new_n786), .B2(new_n262), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n262), .A2(G127gat), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n789), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT109), .ZN(G1342gat));
  OR2_X1    g598(.A1(new_n789), .A2(G134gat), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n800), .A2(KEYINPUT56), .A3(new_n665), .ZN(new_n801));
  XOR2_X1   g600(.A(new_n801), .B(KEYINPUT110), .Z(new_n802));
  OAI21_X1  g601(.A(G134gat), .B1(new_n786), .B2(new_n665), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT56), .B1(new_n800), .B2(new_n665), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(KEYINPUT111), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n802), .A2(new_n803), .A3(new_n805), .ZN(G1343gat));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n807), .B1(new_n761), .B2(new_n763), .ZN(new_n808));
  AOI211_X1 g607(.A(KEYINPUT112), .B(new_n762), .C1(new_n759), .C2(new_n760), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n808), .A2(new_n809), .A3(KEYINPUT55), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n761), .A2(KEYINPUT55), .A3(new_n763), .ZN(new_n811));
  INV_X1    g610(.A(new_n767), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n811), .A2(new_n592), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n776), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n778), .B1(new_n665), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n781), .B1(new_n815), .B2(new_n703), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n816), .A2(KEYINPUT57), .A3(new_n682), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT113), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n816), .A2(new_n819), .A3(KEYINPUT57), .A4(new_n682), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n783), .A2(new_n505), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n818), .B(new_n820), .C1(KEYINPUT57), .C2(new_n821), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n562), .A2(new_n785), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(new_n592), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n824), .A2(new_n825), .A3(G141gat), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n825), .B1(new_n824), .B2(G141gat), .ZN(new_n827));
  NOR4_X1   g626(.A1(new_n783), .A2(new_n533), .A3(new_n662), .A4(new_n505), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n532), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n829), .A2(G141gat), .A3(new_n593), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n826), .A2(new_n827), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT58), .B1(new_n824), .B2(G141gat), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n834));
  INV_X1    g633(.A(new_n830), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n834), .B1(new_n833), .B2(new_n835), .ZN(new_n837));
  OAI22_X1  g636(.A1(new_n831), .A2(new_n832), .B1(new_n836), .B2(new_n837), .ZN(G1344gat));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n808), .A2(new_n809), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n813), .B1(new_n840), .B2(new_n765), .ZN(new_n841));
  INV_X1    g640(.A(new_n776), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n665), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AND4_X1   g642(.A1(new_n339), .A2(new_n766), .A3(new_n769), .A4(new_n775), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n703), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n780), .A2(new_n592), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT118), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n844), .B1(new_n814), .B2(new_n665), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n781), .B(new_n849), .C1(new_n703), .C2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n848), .A2(new_n682), .A3(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT57), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n852), .A2(KEYINPUT119), .A3(new_n853), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n782), .A2(KEYINPUT57), .A3(new_n748), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n782), .A2(KEYINPUT117), .A3(KEYINPUT57), .A4(new_n748), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n739), .B1(new_n858), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n343), .B1(new_n864), .B2(new_n823), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n839), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n822), .A2(new_n823), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n866), .B(G148gat), .C1(new_n868), .C2(new_n739), .ZN(new_n869));
  INV_X1    g668(.A(new_n857), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT119), .B1(new_n852), .B2(new_n853), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n863), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n618), .A3(new_n823), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(G148gat), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(KEYINPUT120), .A3(KEYINPUT59), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n867), .A2(new_n869), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n828), .A2(new_n343), .A3(new_n793), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT116), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(G1345gat));
  OAI21_X1  g678(.A(G155gat), .B1(new_n868), .B2(new_n262), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n262), .A2(G155gat), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n880), .B1(new_n829), .B2(new_n881), .ZN(G1346gat));
  OAI21_X1  g681(.A(G162gat), .B1(new_n868), .B2(new_n644), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n665), .A2(G162gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n883), .B1(new_n829), .B2(new_n884), .ZN(G1347gat));
  NOR2_X1   g684(.A1(new_n653), .A2(new_n532), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n784), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(G169gat), .B1(new_n887), .B2(new_n593), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n782), .A2(new_n567), .A3(new_n886), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n432), .A3(new_n592), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(G1348gat));
  AOI21_X1  g690(.A(G176gat), .B1(new_n889), .B2(new_n618), .ZN(new_n892));
  INV_X1    g691(.A(new_n887), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n739), .A2(new_n433), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(G1349gat));
  NAND3_X1  g694(.A1(new_n889), .A2(new_n423), .A3(new_n703), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT121), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n893), .A2(new_n703), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n897), .B1(new_n898), .B2(G183gat), .ZN(new_n899));
  XNOR2_X1  g698(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n899), .B(new_n900), .ZN(G1350gat));
  OAI21_X1  g700(.A(G190gat), .B1(new_n887), .B2(new_n665), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT61), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n889), .A2(new_n424), .A3(new_n643), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1351gat));
  AND2_X1   g704(.A1(new_n562), .A2(new_n886), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n821), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT123), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n584), .A3(new_n592), .ZN(new_n909));
  XOR2_X1   g708(.A(new_n906), .B(KEYINPUT124), .Z(new_n910));
  AND2_X1   g709(.A1(new_n872), .A2(new_n910), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n911), .A2(new_n592), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n909), .B1(new_n912), .B2(new_n584), .ZN(G1352gat));
  INV_X1    g712(.A(G204gat), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n907), .A2(new_n914), .A3(new_n618), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT62), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n914), .B1(new_n864), .B2(new_n910), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT125), .ZN(new_n918));
  OR3_X1    g717(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n916), .B2(new_n917), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(G1353gat));
  NAND3_X1  g720(.A1(new_n908), .A2(new_n416), .A3(new_n703), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n911), .A2(new_n703), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n923), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT63), .B1(new_n923), .B2(G211gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(G1354gat));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n644), .A2(G218gat), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n908), .A2(new_n928), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n911), .A2(new_n339), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n927), .B(new_n929), .C1(new_n930), .C2(new_n417), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n417), .B1(new_n911), .B2(new_n339), .ZN(new_n932));
  INV_X1    g731(.A(new_n929), .ZN(new_n933));
  OAI21_X1  g732(.A(KEYINPUT126), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n931), .A2(new_n934), .ZN(G1355gat));
endmodule


