//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 0 1 1 0 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n566, new_n568, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n592, new_n593, new_n594, new_n595, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n630,
    new_n631, new_n634, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1180, new_n1181, new_n1182, new_n1183;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT64), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT65), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n460), .B1(G567), .B2(new_n456), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT66), .B(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n462), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n465), .A2(G2104), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n466), .B1(new_n476), .B2(KEYINPUT67), .ZN(new_n477));
  OR3_X1    g052(.A1(new_n463), .A2(KEYINPUT67), .A3(KEYINPUT3), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n462), .A2(G137), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n475), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n482));
  OR2_X1    g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n481), .A2(new_n482), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n471), .B1(new_n483), .B2(new_n484), .ZN(G160));
  OAI221_X1 g060(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n462), .C2(G112), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT69), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n479), .A2(new_n462), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n477), .A2(new_n472), .A3(new_n478), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI22_X1  g065(.A1(G124), .A2(new_n488), .B1(new_n490), .B2(G136), .ZN(new_n491));
  AND2_X1   g066(.A1(new_n487), .A2(new_n491), .ZN(G162));
  NAND3_X1  g067(.A1(new_n477), .A2(G126), .A3(new_n478), .ZN(new_n493));
  NAND2_X1  g068(.A1(G114), .A2(G2104), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n495), .A2(G2105), .B1(G102), .B2(new_n474), .ZN(new_n496));
  OR2_X1    g071(.A1(new_n496), .A2(KEYINPUT70), .ZN(new_n497));
  INV_X1    g072(.A(new_n479), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n462), .A2(KEYINPUT4), .A3(G138), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n468), .A2(new_n462), .A3(G138), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n498), .A2(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n496), .A2(KEYINPUT70), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n497), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  XNOR2_X1  g081(.A(KEYINPUT5), .B(G543), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  AND2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n515), .B(new_n517), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n512), .A2(new_n513), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n510), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  AND2_X1   g099(.A1(G63), .A2(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n507), .A2(new_n525), .ZN(new_n526));
  AND3_X1   g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  AND2_X1   g102(.A1(KEYINPUT71), .A2(KEYINPUT7), .ZN(new_n528));
  NOR2_X1   g103(.A1(KEYINPUT71), .A2(KEYINPUT7), .ZN(new_n529));
  NOR3_X1   g104(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  OR2_X1    g106(.A1(KEYINPUT71), .A2(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g107(.A1(KEYINPUT71), .A2(KEYINPUT7), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n526), .B1(new_n530), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g110(.A(G51), .B(G543), .C1(new_n518), .C2(new_n519), .ZN(new_n536));
  INV_X1    g111(.A(G89), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n520), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g113(.A(KEYINPUT72), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n532), .A2(new_n531), .A3(new_n533), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n540), .A2(new_n541), .B1(new_n507), .B2(new_n525), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT72), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n507), .A2(new_n511), .A3(G89), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n542), .A2(new_n543), .A3(new_n544), .A4(new_n536), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n539), .A2(new_n545), .ZN(G168));
  OAI211_X1 g121(.A(G52), .B(G543), .C1(new_n518), .C2(new_n519), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n520), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n515), .A2(new_n517), .A3(G64), .ZN(new_n550));
  NAND2_X1  g125(.A1(G77), .A2(G543), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n509), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n549), .A2(new_n552), .ZN(G171));
  INV_X1    g128(.A(new_n520), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G81), .ZN(new_n555));
  INV_X1    g130(.A(new_n512), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G43), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n515), .A2(new_n517), .A3(G56), .ZN(new_n558));
  NAND2_X1  g133(.A1(G68), .A2(G543), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n560), .A2(KEYINPUT73), .A3(G651), .ZN(new_n561));
  AOI21_X1  g136(.A(KEYINPUT73), .B1(new_n560), .B2(G651), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n555), .B(new_n557), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  AND3_X1   g140(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G36), .ZN(G176));
  XOR2_X1   g142(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n568));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n568), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(G188));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT76), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G65), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n515), .A2(new_n517), .A3(new_n573), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n576), .A2(KEYINPUT77), .A3(new_n577), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n580), .A2(G651), .A3(new_n581), .ZN(new_n582));
  OAI211_X1 g157(.A(G53), .B(G543), .C1(new_n518), .C2(new_n519), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT9), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n554), .A2(KEYINPUT75), .A3(G91), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT75), .ZN(new_n586));
  INV_X1    g161(.A(G91), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n520), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n582), .A2(new_n584), .A3(new_n589), .ZN(G299));
  INV_X1    g165(.A(G171), .ZN(G301));
  NAND3_X1  g166(.A1(new_n539), .A2(KEYINPUT78), .A3(new_n545), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(KEYINPUT78), .B1(new_n539), .B2(new_n545), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G286));
  NAND2_X1  g171(.A1(new_n556), .A2(G49), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n554), .A2(G87), .ZN(new_n598));
  OAI21_X1  g173(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(G288));
  AOI22_X1  g175(.A1(new_n507), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(new_n509), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n602), .B1(G86), .B2(new_n554), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n556), .A2(G48), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(G305));
  INV_X1    g180(.A(G47), .ZN(new_n606));
  INV_X1    g181(.A(G85), .ZN(new_n607));
  OAI22_X1  g182(.A1(new_n512), .A2(new_n606), .B1(new_n520), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT79), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n608), .B(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n611), .A2(new_n509), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n610), .A2(new_n612), .ZN(G290));
  NAND2_X1  g188(.A1(G301), .A2(G868), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n615));
  INV_X1    g190(.A(G92), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n520), .B2(new_n616), .ZN(new_n617));
  NAND4_X1  g192(.A1(new_n507), .A2(new_n511), .A3(KEYINPUT10), .A4(G92), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AND2_X1   g194(.A1(new_n507), .A2(G66), .ZN(new_n620));
  NAND2_X1  g195(.A1(G79), .A2(G543), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT80), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(G651), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n556), .A2(G54), .ZN(new_n625));
  AND3_X1   g200(.A1(new_n619), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n614), .B1(new_n626), .B2(G868), .ZN(G284));
  OAI21_X1  g202(.A(new_n614), .B1(new_n626), .B2(G868), .ZN(G321));
  NAND2_X1  g203(.A1(G286), .A2(G868), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT81), .Z(new_n630));
  AND3_X1   g205(.A1(new_n582), .A2(new_n584), .A3(new_n589), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(G868), .B2(new_n631), .ZN(G297));
  OAI21_X1  g207(.A(new_n630), .B1(G868), .B2(new_n631), .ZN(G280));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n626), .B1(new_n634), .B2(G860), .ZN(G148));
  NAND3_X1  g210(.A1(new_n619), .A2(new_n624), .A3(new_n625), .ZN(new_n636));
  OAI21_X1  g211(.A(G868), .B1(new_n636), .B2(G559), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n564), .B2(G868), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g214(.A1(new_n490), .A2(G135), .ZN(new_n640));
  INV_X1    g215(.A(KEYINPUT83), .ZN(new_n641));
  AOI22_X1  g216(.A1(new_n640), .A2(new_n641), .B1(G123), .B2(new_n488), .ZN(new_n642));
  OAI221_X1 g217(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n462), .C2(G111), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n642), .B(new_n643), .C1(new_n641), .C2(new_n640), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2096), .Z(new_n645));
  NOR2_X1   g220(.A1(new_n467), .A2(new_n473), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(KEYINPUT13), .B(G2100), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n645), .A2(new_n650), .ZN(G156));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XOR2_X1   g228(.A(G2443), .B(G2446), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(KEYINPUT84), .B(G2438), .Z(new_n658));
  XNOR2_X1  g233(.A(G2427), .B(G2430), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(KEYINPUT15), .B(G2435), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(KEYINPUT14), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n657), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(G14), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(G401));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2067), .B(G2678), .Z(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n669), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n671), .A2(new_n672), .A3(KEYINPUT17), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT18), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2072), .B(G2078), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n675), .B(new_n676), .C1(new_n674), .C2(new_n670), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(new_n676), .B2(new_n675), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2096), .B(G2100), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G227));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n682), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n683), .A2(new_n684), .ZN(new_n688));
  AOI22_X1  g263(.A1(new_n686), .A2(KEYINPUT20), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n688), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n690), .A2(new_n682), .A3(new_n685), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n689), .B(new_n691), .C1(KEYINPUT20), .C2(new_n686), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1986), .B(G1996), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n692), .B(new_n693), .Z(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G1981), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1991), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n694), .A2(new_n697), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(G229));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G25), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n488), .A2(G119), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n490), .A2(G131), .ZN(new_n704));
  OAI221_X1 g279(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n462), .C2(G107), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n702), .B1(new_n707), .B2(new_n701), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT35), .B(G1991), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT85), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n708), .B(new_n710), .Z(new_n711));
  INV_X1    g286(.A(G1986), .ZN(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n610), .B2(new_n612), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n713), .B2(G24), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n711), .B1(new_n712), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n713), .A2(G6), .ZN(new_n717));
  INV_X1    g292(.A(G305), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n717), .B1(new_n718), .B2(new_n713), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT32), .B(G1981), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n713), .A2(G22), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G166), .B2(new_n713), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT87), .B(G1971), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n713), .A2(G23), .ZN(new_n726));
  INV_X1    g301(.A(G288), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n726), .B1(new_n727), .B2(new_n713), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT86), .B(KEYINPUT33), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1976), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n728), .B(new_n730), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n721), .A2(new_n725), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n716), .B1(KEYINPUT34), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(KEYINPUT34), .B2(new_n732), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n712), .B2(new_n715), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT36), .Z(new_n736));
  NAND2_X1  g311(.A1(new_n701), .A2(G35), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G162), .B2(new_n701), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT29), .B(G2090), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n462), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n741), .A2(new_n477), .A3(G129), .A4(new_n478), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n477), .A2(G141), .A3(new_n472), .A4(new_n478), .ZN(new_n743));
  NAND3_X1  g318(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT26), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n474), .A2(G105), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n742), .A2(new_n743), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G29), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G29), .B2(G32), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT27), .B(G1996), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n740), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n626), .A2(new_n713), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G4), .B2(new_n713), .ZN(new_n754));
  INV_X1    g329(.A(G1348), .ZN(new_n755));
  OAI22_X1  g330(.A1(new_n754), .A2(new_n755), .B1(new_n701), .B2(new_n644), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n755), .B2(new_n754), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n750), .A2(new_n751), .ZN(new_n758));
  NOR2_X1   g333(.A1(G5), .A2(G16), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G171), .B2(G16), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(G1961), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n760), .A2(G1961), .ZN(new_n762));
  INV_X1    g337(.A(G28), .ZN(new_n763));
  AOI21_X1  g338(.A(G29), .B1(new_n763), .B2(KEYINPUT30), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(KEYINPUT30), .B2(new_n763), .ZN(new_n765));
  AND4_X1   g340(.A1(new_n758), .A2(new_n761), .A3(new_n762), .A4(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n752), .A2(new_n757), .A3(new_n766), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT31), .B(G11), .Z(new_n768));
  NOR2_X1   g343(.A1(G16), .A2(G21), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G168), .B2(G16), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G1966), .ZN(new_n771));
  NAND2_X1  g346(.A1(KEYINPUT24), .A2(G34), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(KEYINPUT24), .A2(G34), .ZN(new_n774));
  NOR3_X1   g349(.A1(new_n773), .A2(new_n774), .A3(G29), .ZN(new_n775));
  INV_X1    g350(.A(G160), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(G29), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n771), .B1(new_n778), .B2(G2084), .ZN(new_n779));
  INV_X1    g354(.A(G2084), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n713), .A2(G19), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n564), .B2(new_n713), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n777), .A2(new_n780), .B1(G1341), .B2(new_n782), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n779), .B(new_n783), .C1(G1341), .C2(new_n782), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n701), .A2(G27), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G164), .B2(new_n701), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G2078), .ZN(new_n787));
  NOR4_X1   g362(.A1(new_n767), .A2(new_n768), .A3(new_n784), .A4(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(KEYINPUT23), .B1(new_n631), .B2(new_n713), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n713), .A2(G20), .ZN(new_n790));
  MUX2_X1   g365(.A(KEYINPUT23), .B(new_n789), .S(new_n790), .Z(new_n791));
  XOR2_X1   g366(.A(KEYINPUT93), .B(G1956), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(G29), .A2(G33), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT25), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n490), .A2(G139), .ZN(new_n797));
  NAND2_X1  g372(.A1(G115), .A2(G2104), .ZN(new_n798));
  INV_X1    g373(.A(G127), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n467), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(new_n741), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n796), .A2(new_n797), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(KEYINPUT91), .ZN(new_n803));
  INV_X1    g378(.A(G139), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n801), .B1(new_n804), .B2(new_n489), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n795), .B(KEYINPUT25), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT91), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n803), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n794), .B1(new_n810), .B2(G29), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT92), .B(G2072), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n701), .A2(G26), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n490), .A2(KEYINPUT88), .A3(G140), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT88), .ZN(new_n818));
  INV_X1    g393(.A(G140), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n489), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  OAI221_X1 g396(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n462), .C2(G116), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT89), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n488), .A2(G128), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n821), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n816), .B1(new_n826), .B2(G29), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G2067), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n813), .A2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n736), .A2(new_n788), .A3(new_n793), .A4(new_n830), .ZN(G150));
  INV_X1    g406(.A(G150), .ZN(G311));
  NAND2_X1  g407(.A1(new_n626), .A2(G559), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT38), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n835), .A2(new_n509), .ZN(new_n836));
  INV_X1    g411(.A(G55), .ZN(new_n837));
  INV_X1    g412(.A(G93), .ZN(new_n838));
  OAI22_X1  g413(.A1(new_n512), .A2(new_n837), .B1(new_n520), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n563), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n834), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT39), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT94), .ZN(new_n846));
  INV_X1    g421(.A(G860), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n846), .B(new_n847), .C1(new_n844), .C2(new_n843), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n840), .A2(new_n847), .ZN(new_n849));
  XNOR2_X1  g424(.A(KEYINPUT95), .B(KEYINPUT37), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n848), .A2(new_n851), .ZN(G145));
  XOR2_X1   g427(.A(G160), .B(new_n648), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(G162), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n821), .A2(new_n824), .A3(new_n825), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n747), .B1(new_n496), .B2(new_n503), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n496), .A2(new_n503), .A3(new_n747), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n856), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n859), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n826), .B1(new_n861), .B2(new_n857), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n810), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n807), .A2(KEYINPUT98), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n488), .A2(G130), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT99), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n488), .A2(KEYINPUT99), .A3(G130), .ZN(new_n871));
  AOI22_X1  g446(.A1(new_n870), .A2(new_n871), .B1(G142), .B2(new_n490), .ZN(new_n872));
  OAI221_X1 g447(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n462), .C2(G118), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n872), .A2(new_n706), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n706), .B1(new_n872), .B2(new_n873), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n802), .A2(KEYINPUT98), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n860), .A2(new_n862), .A3(new_n877), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n867), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n876), .B1(new_n867), .B2(new_n878), .ZN(new_n880));
  XOR2_X1   g455(.A(KEYINPUT96), .B(KEYINPUT97), .Z(new_n881));
  XNOR2_X1  g456(.A(new_n644), .B(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NOR3_X1   g458(.A1(new_n879), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  AOI211_X1 g459(.A(new_n865), .B(new_n810), .C1(new_n860), .C2(new_n862), .ZN(new_n885));
  INV_X1    g460(.A(new_n878), .ZN(new_n886));
  OAI22_X1  g461(.A1(new_n885), .A2(new_n886), .B1(new_n875), .B2(new_n874), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n867), .A2(new_n876), .A3(new_n878), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n882), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n855), .B1(new_n884), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(G37), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n883), .B1(new_n879), .B2(new_n880), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n887), .A2(new_n888), .A3(new_n882), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(new_n893), .A3(new_n854), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n890), .A2(new_n891), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n890), .A2(KEYINPUT100), .A3(new_n891), .A4(new_n894), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XOR2_X1   g474(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n900));
  XNOR2_X1  g475(.A(new_n899), .B(new_n900), .ZN(G395));
  XNOR2_X1  g476(.A(G303), .B(G288), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(G290), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(G305), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n904), .A2(KEYINPUT102), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT42), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT41), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT9), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n583), .B(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n577), .ZN(new_n910));
  XNOR2_X1  g485(.A(KEYINPUT76), .B(G65), .ZN(new_n911));
  AOI211_X1 g486(.A(new_n579), .B(new_n910), .C1(new_n507), .C2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT77), .B1(new_n576), .B2(new_n577), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n909), .B1(new_n914), .B2(G651), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n626), .B1(new_n915), .B2(new_n589), .ZN(new_n916));
  NOR2_X1   g491(.A1(G299), .A2(new_n636), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n907), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n631), .A2(new_n626), .ZN(new_n919));
  NAND2_X1  g494(.A1(G299), .A2(new_n636), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(KEYINPUT41), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n916), .A2(new_n917), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n563), .B(new_n840), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n636), .A2(G559), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n925), .B(new_n926), .ZN(new_n927));
  MUX2_X1   g502(.A(new_n923), .B(new_n924), .S(new_n927), .Z(new_n928));
  XNOR2_X1  g503(.A(new_n906), .B(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(G868), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n930), .B1(G868), .B2(new_n840), .ZN(G295));
  OAI21_X1  g506(.A(new_n930), .B1(G868), .B2(new_n840), .ZN(G331));
  AOI21_X1  g507(.A(KEYINPUT103), .B1(G168), .B2(G301), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT103), .ZN(new_n934));
  AOI211_X1 g509(.A(new_n934), .B(G171), .C1(new_n539), .C2(new_n545), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT78), .ZN(new_n937));
  NAND2_X1  g512(.A1(G168), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(G301), .B1(new_n938), .B2(new_n592), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n925), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(G168), .A2(G301), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n934), .ZN(new_n942));
  NAND3_X1  g517(.A1(G168), .A2(KEYINPUT103), .A3(G301), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(G171), .B1(new_n593), .B2(new_n594), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(new_n842), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n940), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n923), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n940), .A2(new_n946), .A3(new_n924), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT106), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n948), .B(new_n949), .C1(new_n904), .C2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n903), .B(new_n718), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n948), .A2(new_n949), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n940), .A2(new_n946), .A3(new_n924), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n952), .B(new_n953), .C1(KEYINPUT106), .C2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n951), .A2(new_n955), .A3(new_n891), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT104), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n922), .B1(new_n946), .B2(new_n940), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n958), .B1(new_n954), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n948), .A2(KEYINPUT104), .A3(new_n949), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(new_n952), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n891), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT105), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n952), .A2(new_n953), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n962), .A2(KEYINPUT105), .A3(new_n891), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n965), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n957), .B(KEYINPUT44), .C1(new_n969), .C2(KEYINPUT43), .ZN(new_n970));
  OR2_X1    g545(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n962), .A2(KEYINPUT105), .A3(new_n891), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT105), .B1(new_n962), .B2(new_n891), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n972), .A2(new_n973), .A3(new_n966), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT43), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n971), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n976), .A2(KEYINPUT107), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT107), .B1(new_n976), .B2(new_n977), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n970), .B1(new_n978), .B2(new_n979), .ZN(G397));
  AOI21_X1  g555(.A(G1384), .B1(new_n496), .B2(new_n503), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(G160), .A2(G40), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n706), .B(new_n710), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n826), .B(G2067), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n747), .B(G1996), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n987), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n992), .B(KEYINPUT109), .ZN(new_n993));
  XNOR2_X1  g568(.A(G290), .B(G1986), .ZN(new_n994));
  AOI211_X1 g569(.A(new_n989), .B(new_n993), .C1(new_n987), .C2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n996));
  AND2_X1   g571(.A1(G160), .A2(G40), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n981), .ZN(new_n998));
  INV_X1    g573(.A(G1976), .ZN(new_n999));
  NOR2_X1   g574(.A1(G288), .A2(new_n999), .ZN(new_n1000));
  OR2_X1    g575(.A1(new_n1000), .A2(KEYINPUT111), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(KEYINPUT111), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n998), .A2(G8), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(G288), .A2(new_n999), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n996), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1003), .A2(KEYINPUT112), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n986), .A2(new_n982), .ZN(new_n1008));
  INV_X1    g583(.A(G8), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1010), .A2(new_n1011), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1010), .A2(KEYINPUT111), .A3(new_n999), .A4(G288), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1012), .A2(new_n1013), .A3(new_n996), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1007), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(G1981), .B1(new_n602), .B2(KEYINPUT113), .ZN(new_n1016));
  XNOR2_X1  g591(.A(G305), .B(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT49), .ZN(new_n1018));
  XOR2_X1   g593(.A(G305), .B(new_n1016), .Z(new_n1019));
  INV_X1    g594(.A(KEYINPUT49), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT114), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n1017), .A2(new_n1022), .A3(KEYINPUT49), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1018), .B(new_n1010), .C1(new_n1021), .C2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1015), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT115), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n997), .B1(KEYINPUT50), .B2(new_n982), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT50), .ZN(new_n1028));
  INV_X1    g603(.A(G1384), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1028), .B1(new_n505), .B2(new_n1029), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n1027), .A2(new_n1030), .A3(G2084), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT45), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n986), .B1(new_n1032), .B2(new_n982), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n505), .A2(new_n1029), .A3(new_n983), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1966), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(G8), .B(new_n595), .C1(new_n1031), .C2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n505), .A2(new_n1029), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT50), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n986), .B1(new_n1028), .B2(new_n981), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1040), .A2(G2090), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1037), .A2(new_n984), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n986), .B1(KEYINPUT45), .B2(new_n981), .ZN(new_n1043));
  AOI21_X1  g618(.A(G1971), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(G8), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G303), .A2(G8), .ZN(new_n1046));
  XNOR2_X1  g621(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1046), .B(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1036), .B1(new_n1045), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1024), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1051), .B1(new_n1007), .B2(new_n1014), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI211_X1 g629(.A(G8), .B(new_n1048), .C1(new_n1041), .C2(new_n1044), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1055), .A2(KEYINPUT63), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1026), .A2(new_n1050), .A3(new_n1054), .A4(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1044), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n981), .A2(new_n1028), .ZN(new_n1059));
  OR3_X1    g634(.A1(new_n986), .A2(new_n1059), .A3(KEYINPUT116), .ZN(new_n1060));
  INV_X1    g635(.A(G2090), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n505), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT116), .B1(new_n986), .B2(new_n1059), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1009), .B1(new_n1058), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1055), .B1(new_n1065), .B2(new_n1048), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1025), .A2(new_n1066), .A3(new_n1036), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1057), .B1(KEYINPUT63), .B2(new_n1067), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n545), .B(new_n539), .C1(new_n1031), .C2(new_n1035), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1070));
  INV_X1    g645(.A(G1966), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1038), .A2(new_n780), .A3(new_n1039), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1072), .A2(G168), .A3(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1069), .A2(new_n1074), .A3(G8), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n1076));
  OAI21_X1  g651(.A(G8), .B1(new_n1031), .B2(new_n1035), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1076), .B1(new_n1077), .B2(KEYINPUT121), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1074), .A2(G8), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT62), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1025), .A2(new_n1066), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1080), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1077), .A2(KEYINPUT121), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1084), .B1(new_n1085), .B2(new_n1076), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT62), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT123), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n1070), .B2(G2078), .ZN(new_n1091));
  INV_X1    g666(.A(G2078), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1033), .A2(KEYINPUT123), .A3(new_n1034), .A4(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1091), .A2(KEYINPUT53), .A3(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1042), .A2(new_n1092), .A3(new_n1043), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n1096));
  INV_X1    g671(.A(G1961), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1095), .A2(new_n1096), .B1(new_n1040), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(G301), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1082), .A2(new_n1083), .A3(new_n1089), .A4(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1024), .A2(new_n999), .A3(new_n727), .ZN(new_n1101));
  OR2_X1    g676(.A1(G305), .A2(G1981), .ZN(new_n1102));
  AOI211_X1 g677(.A(new_n1009), .B(new_n1008), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1052), .B(KEYINPUT115), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1055), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1103), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1068), .A2(new_n1100), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT124), .B(G2078), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1043), .A2(KEYINPUT53), .A3(new_n985), .A4(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1098), .A2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1112), .A2(G171), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1109), .B1(new_n1113), .B2(new_n1099), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(G171), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1094), .A2(G301), .A3(new_n1098), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1115), .A2(KEYINPUT54), .A3(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1108), .A2(new_n1114), .A3(new_n1083), .A4(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1119));
  XOR2_X1   g694(.A(KEYINPUT119), .B(G1996), .Z(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT58), .B(G1341), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1008), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n564), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n998), .A2(G2067), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1128), .B1(new_n1040), .B2(new_n755), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT60), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1129), .A2(new_n1130), .A3(new_n626), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1126), .A2(new_n1127), .A3(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1060), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1133));
  INV_X1    g708(.A(G1956), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT56), .B(G2072), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1042), .A2(new_n1043), .A3(new_n1136), .ZN(new_n1137));
  XOR2_X1   g712(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n1138));
  NAND2_X1  g713(.A1(G299), .A2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT118), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT57), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1140), .B1(new_n1141), .B2(G299), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1135), .A2(new_n1137), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1144));
  OAI21_X1  g719(.A(KEYINPUT120), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT61), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1129), .A2(new_n636), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1129), .A2(new_n636), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT60), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n1150));
  OAI211_X1 g725(.A(KEYINPUT120), .B(new_n1150), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1132), .A2(new_n1146), .A3(new_n1149), .A4(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1143), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1153), .B1(new_n1144), .B2(new_n1148), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1118), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n995), .B1(new_n1107), .B2(new_n1155), .ZN(new_n1156));
  NOR4_X1   g731(.A1(new_n985), .A2(new_n986), .A3(G1986), .A4(G290), .ZN(new_n1157));
  XOR2_X1   g732(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1158));
  XNOR2_X1  g733(.A(new_n1157), .B(new_n1158), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n993), .A2(new_n1159), .A3(new_n989), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n987), .B1(new_n990), .B2(new_n747), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT125), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n985), .A2(new_n986), .A3(G1996), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1163), .B(KEYINPUT46), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1165), .B(KEYINPUT47), .ZN(new_n1166));
  OR2_X1    g741(.A1(new_n706), .A2(new_n710), .ZN(new_n1167));
  OAI22_X1  g742(.A1(new_n993), .A2(new_n1167), .B1(G2067), .B2(new_n826), .ZN(new_n1168));
  AOI211_X1 g743(.A(new_n1160), .B(new_n1166), .C1(new_n987), .C2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1156), .A2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g745(.A(G227), .B1(new_n897), .B2(new_n898), .ZN(new_n1172));
  OAI211_X1 g746(.A(new_n665), .B(G319), .C1(new_n698), .C2(new_n699), .ZN(new_n1173));
  INV_X1    g747(.A(new_n1173), .ZN(new_n1174));
  AND4_X1   g748(.A1(KEYINPUT127), .A2(new_n1172), .A3(new_n976), .A4(new_n1174), .ZN(new_n1175));
  NAND2_X1  g749(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n1176));
  AOI21_X1  g750(.A(new_n1173), .B1(new_n1176), .B2(new_n971), .ZN(new_n1177));
  AOI21_X1  g751(.A(KEYINPUT127), .B1(new_n1177), .B2(new_n1172), .ZN(new_n1178));
  NOR2_X1   g752(.A1(new_n1175), .A2(new_n1178), .ZN(G308));
  NAND3_X1  g753(.A1(new_n1172), .A2(new_n976), .A3(new_n1174), .ZN(new_n1180));
  INV_X1    g754(.A(KEYINPUT127), .ZN(new_n1181));
  NAND2_X1  g755(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g756(.A1(new_n1177), .A2(KEYINPUT127), .A3(new_n1172), .ZN(new_n1183));
  NAND2_X1  g757(.A1(new_n1182), .A2(new_n1183), .ZN(G225));
endmodule


