//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 1 1 0 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1276, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT0), .Z(new_n217));
  AND2_X1   g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G20), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT65), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n206), .A2(new_n207), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n217), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT66), .Z(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  INV_X1    g0025(.A(G87), .ZN(new_n226));
  INV_X1    g0026(.A(G250), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n224), .B1(new_n202), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  INV_X1    g0030(.A(G97), .ZN(new_n231));
  INV_X1    g0031(.A(G257), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n229), .B1(new_n201), .B2(new_n230), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n214), .B1(new_n228), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT1), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n223), .A2(new_n235), .ZN(G361));
  XOR2_X1   g0036(.A(G226), .B(G232), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G238), .B(G244), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n207), .A2(G68), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n202), .A2(G50), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n249), .B(new_n254), .ZN(G351));
  NAND2_X1  g0055(.A1(G1), .A2(G13), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n256), .B1(G33), .B2(G41), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT3), .B(G33), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(G226), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G97), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NOR3_X1   g0067(.A1(new_n267), .A2(new_n230), .A3(new_n259), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n257), .B1(new_n262), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n218), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  AOI21_X1  g0073(.A(G1), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n271), .A2(G274), .A3(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n257), .A2(new_n274), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n276), .B1(G238), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n269), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT13), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT13), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n269), .A2(new_n278), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT14), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(new_n284), .A3(G169), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT75), .ZN(new_n286));
  INV_X1    g0086(.A(G169), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n287), .B1(new_n280), .B2(new_n282), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT75), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(new_n289), .A3(new_n284), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G179), .ZN(new_n292));
  OAI22_X1  g0092(.A1(new_n288), .A2(new_n284), .B1(new_n283), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  AND3_X1   g0095(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n202), .ZN(new_n297));
  XOR2_X1   g0097(.A(new_n297), .B(KEYINPUT12), .Z(new_n298));
  NAND3_X1  g0098(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n256), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n212), .A2(G33), .A3(G77), .ZN(new_n302));
  NOR2_X1   g0102(.A1(G20), .A2(G33), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n303), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n301), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n298), .B1(KEYINPUT11), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT72), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n307), .B1(new_n296), .B2(new_n300), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n309), .A2(KEYINPUT72), .A3(new_n256), .A4(new_n299), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n211), .A2(G20), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n308), .A2(G68), .A3(new_n310), .A4(new_n311), .ZN(new_n312));
  OR2_X1    g0112(.A1(new_n305), .A2(KEYINPUT11), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n306), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT74), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n306), .A2(KEYINPUT74), .A3(new_n312), .A4(new_n313), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n295), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n283), .A2(G200), .ZN(new_n321));
  INV_X1    g0121(.A(G190), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n318), .B(new_n321), .C1(new_n322), .C2(new_n283), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n208), .A2(G20), .ZN(new_n325));
  INV_X1    g0125(.A(G150), .ZN(new_n326));
  INV_X1    g0126(.A(new_n303), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT8), .B(G58), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n328), .B(KEYINPUT69), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n212), .A2(G33), .ZN(new_n330));
  OAI221_X1 g0130(.A(new_n325), .B1(new_n326), .B2(new_n327), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n300), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n301), .A2(new_n311), .ZN(new_n333));
  MUX2_X1   g0133(.A(new_n309), .B(new_n333), .S(G50), .Z(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n258), .A2(G222), .A3(new_n259), .ZN(new_n336));
  INV_X1    g0136(.A(G77), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n258), .A2(G1698), .ZN(new_n338));
  INV_X1    g0138(.A(G223), .ZN(new_n339));
  OAI221_X1 g0139(.A(new_n336), .B1(new_n337), .B2(new_n258), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n257), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n276), .B1(G226), .B2(new_n277), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n287), .ZN(new_n344));
  XNOR2_X1  g0144(.A(KEYINPUT70), .B(G179), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n335), .B(new_n344), .C1(new_n343), .C2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n277), .A2(G244), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n275), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT71), .ZN(new_n350));
  INV_X1    g0150(.A(G107), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n338), .A2(new_n225), .B1(new_n351), .B2(new_n258), .ZN(new_n352));
  NOR3_X1   g0152(.A1(new_n267), .A2(new_n230), .A3(G1698), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n257), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT71), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n348), .A2(new_n355), .A3(new_n275), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n350), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  OR2_X1    g0157(.A1(new_n357), .A2(new_n346), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G20), .A2(G77), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT15), .B(G87), .ZN(new_n360));
  OAI221_X1 g0160(.A(new_n359), .B1(new_n328), .B2(new_n327), .C1(new_n330), .C2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n300), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n308), .A2(G77), .A3(new_n310), .A4(new_n311), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n296), .A2(new_n337), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT73), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n362), .A2(KEYINPUT73), .A3(new_n363), .A4(new_n364), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n357), .A2(new_n287), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n358), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n357), .A2(G200), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n350), .A2(new_n354), .A3(G190), .A4(new_n356), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n372), .A2(new_n368), .A3(new_n367), .A4(new_n373), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT10), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT9), .ZN(new_n377));
  AND3_X1   g0177(.A1(new_n332), .A2(new_n377), .A3(new_n334), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n377), .B1(new_n332), .B2(new_n334), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n343), .A2(new_n322), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n381), .B1(G200), .B2(new_n343), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n376), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n382), .B(new_n376), .C1(new_n378), .C2(new_n379), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n347), .B(new_n375), .C1(new_n383), .C2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n324), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n258), .A2(G226), .A3(G1698), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n264), .A2(new_n266), .A3(G223), .A4(new_n259), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G87), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n257), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n271), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n275), .B1(new_n394), .B2(new_n230), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n287), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n395), .B1(new_n257), .B2(new_n391), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n345), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(KEYINPUT7), .B1(new_n267), .B2(new_n212), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT7), .ZN(new_n404));
  AOI211_X1 g0204(.A(new_n404), .B(G20), .C1(new_n264), .C2(new_n266), .ZN(new_n405));
  OAI21_X1  g0205(.A(G68), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(G159), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n327), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G58), .A2(G68), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n203), .A2(new_n205), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT76), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n412), .A3(G20), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(G20), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT76), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n406), .A2(new_n409), .A3(new_n413), .A4(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT16), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n404), .B1(new_n258), .B2(G20), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n267), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n408), .B1(new_n420), .B2(G68), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT16), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n411), .A2(new_n412), .A3(G20), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n412), .B1(new_n411), .B2(G20), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n421), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n301), .B1(new_n417), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n329), .A2(new_n333), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n428), .B1(new_n296), .B2(new_n329), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n402), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT18), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n421), .A2(new_n422), .A3(new_n425), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n422), .B1(new_n421), .B2(new_n425), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n300), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n429), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT18), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n437), .A3(new_n402), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n392), .A2(new_n322), .A3(new_n396), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT77), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT77), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n399), .A2(new_n441), .A3(new_n322), .ZN(new_n442));
  INV_X1    g0242(.A(G200), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n397), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n440), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n435), .A2(new_n429), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT17), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n417), .A2(new_n426), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n430), .B1(new_n449), .B2(new_n300), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(KEYINPUT17), .A3(new_n445), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n432), .A2(new_n438), .A3(new_n448), .A4(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  OR2_X1    g0253(.A1(new_n453), .A2(KEYINPUT78), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(KEYINPUT78), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n387), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  OR3_X1    g0257(.A1(new_n309), .A2(KEYINPUT80), .A3(G97), .ZN(new_n458));
  OAI21_X1  g0258(.A(KEYINPUT80), .B1(new_n309), .B2(G97), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n211), .A2(G33), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n301), .A2(new_n309), .A3(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n460), .B1(new_n231), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n420), .A2(G107), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT79), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n327), .A2(new_n337), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n351), .A2(KEYINPUT6), .A3(G97), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT6), .ZN(new_n470));
  XNOR2_X1  g0270(.A(G97), .B(G107), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n465), .B(new_n467), .C1(new_n472), .C2(new_n212), .ZN(new_n473));
  AND2_X1   g0273(.A1(G97), .A2(G107), .ZN(new_n474));
  NOR2_X1   g0274(.A1(G97), .A2(G107), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n470), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n212), .B1(new_n476), .B2(new_n468), .ZN(new_n477));
  OAI21_X1  g0277(.A(KEYINPUT79), .B1(new_n477), .B2(new_n466), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n464), .A2(new_n473), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n463), .B1(new_n479), .B2(new_n300), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n264), .A2(new_n266), .A3(G244), .A4(new_n259), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT4), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G283), .ZN(new_n484));
  INV_X1    g0284(.A(G244), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n258), .A2(new_n259), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n483), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n264), .A2(new_n266), .A3(G250), .A4(G1698), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT81), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT81), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n258), .A2(new_n491), .A3(G250), .A4(G1698), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n257), .B1(new_n488), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(G274), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n495), .B1(new_n218), .B2(new_n270), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n273), .A2(G1), .ZN(new_n497));
  XNOR2_X1  g0297(.A(KEYINPUT5), .B(G41), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  AND2_X1   g0299(.A1(KEYINPUT5), .A2(G41), .ZN(new_n500));
  NOR2_X1   g0300(.A1(KEYINPUT5), .A2(G41), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n497), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n502), .A2(G257), .A3(new_n271), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT82), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n502), .A2(KEYINPUT82), .A3(G257), .A4(new_n271), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n499), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n494), .A2(new_n507), .A3(G190), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n480), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT83), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n494), .A2(new_n507), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n510), .B1(new_n511), .B2(G200), .ZN(new_n512));
  AOI211_X1 g0312(.A(KEYINPUT83), .B(new_n443), .C1(new_n494), .C2(new_n507), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n509), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n479), .A2(new_n300), .ZN(new_n515));
  INV_X1    g0315(.A(new_n463), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n511), .A2(new_n287), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n494), .A2(new_n507), .A3(new_n345), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT84), .B1(new_n514), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n511), .A2(G200), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT83), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n511), .A2(new_n510), .A3(G200), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n523), .A2(new_n480), .A3(new_n508), .A4(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT84), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n521), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(G238), .A2(G1698), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n485), .A2(G1698), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n258), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G116), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n271), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n496), .A2(new_n497), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n227), .B1(new_n211), .B2(G45), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n271), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n540), .A2(KEYINPUT85), .A3(new_n345), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n264), .A2(new_n266), .A3(new_n212), .A4(G68), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT19), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n212), .B1(new_n261), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n475), .A2(new_n226), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n212), .A2(G33), .A3(G97), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT86), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n547), .A2(new_n548), .A3(new_n543), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n548), .B1(new_n547), .B2(new_n543), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n542), .B(new_n546), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n300), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n360), .A2(new_n296), .ZN(new_n553));
  INV_X1    g0353(.A(new_n462), .ZN(new_n554));
  INV_X1    g0354(.A(new_n360), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n552), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n496), .A2(new_n497), .B1(new_n271), .B2(new_n537), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n530), .B1(new_n485), .B2(G1698), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n559), .A2(new_n258), .B1(G33), .B2(G116), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n345), .B(new_n558), .C1(new_n560), .C2(new_n271), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT85), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n558), .B1(new_n560), .B2(new_n271), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n287), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n541), .A2(new_n557), .A3(new_n563), .A4(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n551), .A2(new_n300), .B1(new_n296), .B2(new_n360), .ZN(new_n567));
  OAI21_X1  g0367(.A(G200), .B1(new_n535), .B2(new_n539), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n554), .A2(G87), .ZN(new_n569));
  OAI211_X1 g0369(.A(G190), .B(new_n558), .C1(new_n560), .C2(new_n271), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n567), .A2(new_n568), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n529), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n264), .A2(new_n266), .A3(new_n212), .A4(G87), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT22), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT22), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n258), .A2(new_n577), .A3(new_n212), .A4(G87), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT23), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(G20), .B2(new_n351), .ZN(new_n581));
  NOR3_X1   g0381(.A1(new_n212), .A2(KEYINPUT23), .A3(G107), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n534), .A2(G20), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT24), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n584), .A2(KEYINPUT89), .ZN(new_n585));
  NOR4_X1   g0385(.A1(new_n581), .A2(new_n582), .A3(new_n583), .A4(new_n585), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n584), .A2(KEYINPUT89), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n579), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n587), .B1(new_n579), .B2(new_n586), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n300), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n554), .A2(G107), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT25), .B1(new_n296), .B2(new_n351), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n296), .A2(KEYINPUT25), .A3(new_n351), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n590), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n502), .A2(G264), .A3(new_n271), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n227), .A2(new_n259), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n232), .A2(G1698), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n264), .A2(new_n600), .A3(new_n266), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(G33), .A2(G294), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n271), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n599), .A2(new_n604), .A3(new_n499), .ZN(new_n605));
  OR2_X1    g0405(.A1(new_n605), .A2(new_n287), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT90), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n599), .B2(new_n604), .ZN(new_n608));
  NOR2_X1   g0408(.A1(G250), .A2(G1698), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n609), .B1(new_n232), .B2(G1698), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n610), .A2(new_n258), .B1(G33), .B2(G294), .ZN(new_n611));
  OAI211_X1 g0411(.A(KEYINPUT90), .B(new_n598), .C1(new_n611), .C2(new_n271), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n608), .A2(new_n612), .A3(G179), .A4(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT91), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n606), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n597), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n590), .A2(new_n596), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n608), .A2(new_n613), .A3(new_n612), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n443), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n605), .A2(new_n322), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(G116), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n299), .A2(new_n256), .B1(G20), .B2(new_n626), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n484), .B(new_n212), .C1(G33), .C2(new_n231), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT20), .ZN(new_n630));
  OR2_X1    g0430(.A1(new_n630), .A2(KEYINPUT88), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(KEYINPUT88), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n627), .A2(KEYINPUT88), .A3(new_n628), .A4(new_n630), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n296), .A2(new_n626), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n626), .B1(new_n211), .B2(G33), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n308), .A2(new_n310), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT87), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT87), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n308), .A2(new_n640), .A3(new_n310), .A4(new_n637), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n636), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n502), .A2(G270), .A3(new_n271), .ZN(new_n643));
  MUX2_X1   g0443(.A(G257), .B(G264), .S(G1698), .Z(new_n644));
  NOR2_X1   g0444(.A1(new_n644), .A2(new_n267), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n257), .B1(new_n258), .B2(G303), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n613), .B(new_n643), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(G200), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n642), .B(new_n648), .C1(new_n322), .C2(new_n647), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT21), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n647), .A2(G169), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n650), .B1(new_n642), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n639), .A2(new_n641), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n651), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(KEYINPUT21), .A3(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n647), .A2(new_n292), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n649), .A2(new_n652), .A3(new_n657), .A4(new_n659), .ZN(new_n660));
  NOR4_X1   g0460(.A1(new_n457), .A2(new_n574), .A3(new_n625), .A4(new_n660), .ZN(G372));
  NAND3_X1  g0461(.A1(new_n557), .A2(new_n565), .A3(new_n561), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n571), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n663), .B1(new_n619), .B2(new_n623), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n664), .A2(new_n525), .A3(new_n527), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n652), .A2(new_n657), .A3(new_n659), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n608), .A2(new_n612), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n667), .A2(KEYINPUT91), .A3(G179), .A4(new_n613), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n614), .A2(new_n615), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(new_n669), .A3(new_n606), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n666), .B1(new_n597), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT26), .B1(new_n527), .B2(new_n572), .ZN(new_n674));
  INV_X1    g0474(.A(new_n663), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n518), .A2(new_n519), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT26), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n675), .A2(new_n676), .A3(new_n677), .A4(new_n517), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n674), .A2(new_n678), .A3(new_n662), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n457), .B1(new_n673), .B2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n437), .B1(new_n436), .B2(new_n402), .ZN(new_n682));
  AOI211_X1 g0482(.A(KEYINPUT18), .B(new_n401), .C1(new_n435), .C2(new_n429), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n371), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n323), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n320), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(KEYINPUT17), .B1(new_n450), .B2(new_n445), .ZN(new_n689));
  AND4_X1   g0489(.A1(KEYINPUT17), .A2(new_n435), .A3(new_n429), .A4(new_n445), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n685), .B1(new_n688), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n383), .A2(new_n385), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n347), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n681), .A2(new_n694), .ZN(G369));
  NAND3_X1  g0495(.A1(new_n211), .A2(new_n212), .A3(G13), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT92), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(G213), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(G343), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n655), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT93), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n704), .A2(new_n666), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n660), .ZN(new_n706));
  OAI21_X1  g0506(.A(G330), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  XOR2_X1   g0507(.A(new_n707), .B(KEYINPUT94), .Z(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n618), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n702), .ZN(new_n711));
  INV_X1    g0511(.A(new_n702), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n618), .B(new_n624), .C1(new_n619), .C2(new_n712), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n709), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n666), .A2(new_n712), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n625), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n718), .B1(new_n710), .B2(new_n712), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n716), .A2(new_n719), .ZN(G399));
  INV_X1    g0520(.A(new_n215), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT95), .B1(new_n721), .B2(G41), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n721), .A2(KEYINPUT95), .A3(G41), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n475), .A2(new_n226), .A3(new_n626), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n725), .A2(new_n211), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n727), .B1(new_n221), .B2(new_n725), .ZN(new_n728));
  XOR2_X1   g0528(.A(new_n728), .B(KEYINPUT28), .Z(new_n729));
  NAND3_X1  g0529(.A1(new_n520), .A2(new_n677), .A3(new_n573), .ZN(new_n730));
  OAI21_X1  g0530(.A(KEYINPUT26), .B1(new_n527), .B2(new_n663), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(new_n662), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n672), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT29), .B1(new_n733), .B2(new_n702), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n702), .B1(new_n673), .B2(new_n680), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n734), .B1(new_n736), .B2(KEYINPUT29), .ZN(new_n737));
  INV_X1    g0537(.A(G330), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n564), .A2(new_n647), .A3(new_n345), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n739), .A2(new_n620), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n608), .A2(new_n540), .A3(new_n612), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n645), .A2(new_n646), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(G179), .A3(new_n613), .A4(new_n643), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  AND3_X1   g0544(.A1(new_n494), .A2(new_n507), .A3(KEYINPUT30), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n740), .A2(new_n511), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT30), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n658), .A2(new_n540), .A3(new_n608), .A4(new_n612), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n747), .B1(new_n748), .B2(new_n511), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n712), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(KEYINPUT97), .B1(new_n750), .B2(KEYINPUT31), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n744), .A2(new_n745), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n739), .A2(new_n511), .A3(new_n620), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n749), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n702), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT97), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT31), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n712), .A2(new_n757), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n749), .A2(new_n753), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT96), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n749), .A2(KEYINPUT96), .A3(new_n753), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n762), .A2(new_n763), .A3(new_n752), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n751), .A2(new_n758), .B1(new_n759), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n618), .A2(new_n624), .A3(new_n712), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n660), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n529), .A2(new_n767), .A3(new_n573), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n738), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n737), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n729), .B1(new_n770), .B2(G1), .ZN(G364));
  INV_X1    g0571(.A(G13), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n211), .B1(new_n773), .B2(G45), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n725), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n705), .A2(new_n706), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n776), .B(new_n709), .C1(new_n738), .C2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n256), .B1(G20), .B2(new_n287), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n212), .A2(G179), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n780), .A2(G190), .A3(G200), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n267), .B1(new_n782), .B2(G87), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n783), .A2(KEYINPUT101), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G190), .A2(G200), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n780), .A2(new_n785), .ZN(new_n786));
  OR2_X1    g0586(.A1(new_n786), .A2(KEYINPUT100), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(KEYINPUT100), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G159), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n345), .A2(new_n212), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G200), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n322), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n791), .A2(KEYINPUT32), .B1(new_n207), .B2(new_n795), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n784), .B(new_n796), .C1(KEYINPUT32), .C2(new_n791), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n792), .A2(new_n785), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n780), .A2(new_n322), .A3(G200), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n799), .A2(G77), .B1(G107), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(KEYINPUT101), .B2(new_n783), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT99), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n322), .A2(G200), .ZN(new_n805));
  AND3_X1   g0605(.A1(new_n792), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n804), .B1(new_n792), .B2(new_n805), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n803), .B1(new_n809), .B2(G58), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n805), .A2(new_n292), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G20), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G97), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n792), .A2(new_n322), .A3(G200), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n814), .B2(new_n202), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT102), .ZN(new_n816));
  AND3_X1   g0616(.A1(new_n797), .A2(new_n810), .A3(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n812), .ZN(new_n818));
  INV_X1    g0618(.A(G294), .ZN(new_n819));
  INV_X1    g0619(.A(G283), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n818), .A2(new_n819), .B1(new_n800), .B2(new_n820), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n258), .B(new_n821), .C1(G303), .C2(new_n782), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n809), .A2(G322), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n790), .A2(G329), .B1(G311), .B2(new_n799), .ZN(new_n824));
  INV_X1    g0624(.A(new_n814), .ZN(new_n825));
  XNOR2_X1  g0625(.A(KEYINPUT33), .B(G317), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G326), .A2(new_n794), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n822), .A2(new_n823), .A3(new_n824), .A4(new_n827), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT103), .Z(new_n829));
  OAI21_X1  g0629(.A(new_n779), .B1(new_n817), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n776), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n721), .A2(new_n267), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n832), .A2(G355), .B1(new_n626), .B2(new_n721), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n721), .A2(new_n258), .ZN(new_n834));
  INV_X1    g0634(.A(new_n221), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n834), .B1(new_n835), .B2(G45), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n254), .A2(new_n273), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n833), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OR3_X1    g0638(.A1(KEYINPUT98), .A2(G13), .A3(G33), .ZN(new_n839));
  OAI21_X1  g0639(.A(KEYINPUT98), .B1(G13), .B2(G33), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n842), .A2(G20), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n843), .A2(new_n779), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n831), .B1(new_n838), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n830), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n843), .B(KEYINPUT104), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n846), .B1(new_n777), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n778), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(G396));
  NOR2_X1   g0651(.A1(new_n371), .A2(new_n702), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n369), .A2(new_n702), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n374), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n852), .B1(new_n371), .B2(new_n854), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n735), .B(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n769), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n776), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n857), .B2(new_n856), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n813), .B1(new_n808), .B2(new_n819), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT105), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n800), .A2(new_n226), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n258), .B(new_n862), .C1(G107), .C2(new_n782), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n790), .A2(G311), .B1(G116), .B2(new_n799), .ZN(new_n864));
  AOI22_X1  g0664(.A1(G303), .A2(new_n794), .B1(new_n825), .B2(G283), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n861), .A2(new_n863), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n794), .A2(G137), .B1(new_n799), .B2(G159), .ZN(new_n867));
  INV_X1    g0667(.A(G143), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n867), .B1(new_n326), .B2(new_n814), .C1(new_n808), .C2(new_n868), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n869), .B(KEYINPUT106), .Z(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT34), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n790), .A2(G132), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n267), .B1(new_n812), .B2(G58), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n782), .A2(G50), .B1(new_n801), .B2(G68), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n871), .A2(new_n872), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n870), .A2(KEYINPUT34), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n866), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n779), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n841), .A2(new_n779), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n831), .B1(new_n337), .B2(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n878), .B(new_n880), .C1(new_n842), .C2(new_n855), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n859), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(G384));
  NOR2_X1   g0683(.A1(new_n773), .A2(new_n211), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT37), .ZN(new_n886));
  INV_X1    g0686(.A(new_n700), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n427), .B2(new_n430), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n886), .B1(new_n888), .B2(KEYINPUT107), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n889), .A2(new_n431), .A3(new_n446), .A4(new_n888), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n700), .B1(new_n435), .B2(new_n429), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT107), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT37), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n431), .A2(new_n888), .A3(new_n446), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n888), .B1(new_n684), .B2(new_n691), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n885), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n452), .A2(new_n891), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n899), .A2(KEYINPUT38), .A3(new_n895), .A4(new_n890), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n712), .B(new_n855), .C1(new_n672), .C2(new_n679), .ZN(new_n903));
  INV_X1    g0703(.A(new_n852), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n319), .A2(new_n702), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n293), .B1(new_n286), .B2(new_n290), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n906), .B(new_n323), .C1(new_n907), .C2(new_n318), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n295), .A2(new_n319), .A3(new_n702), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n902), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n685), .B2(new_n700), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n898), .A2(KEYINPUT39), .A3(new_n900), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n886), .B1(new_n436), .B2(new_n402), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n446), .A2(KEYINPUT108), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT108), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n450), .A2(new_n917), .A3(new_n445), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n915), .A2(new_n916), .A3(new_n918), .A4(new_n888), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n894), .A2(new_n886), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n885), .B1(new_n897), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT39), .B1(new_n922), .B2(new_n900), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n914), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n320), .A2(new_n702), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n913), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n694), .B1(new_n456), .B2(new_n737), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n927), .B(new_n928), .Z(new_n929));
  NAND2_X1  g0729(.A1(new_n910), .A2(new_n855), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n529), .A2(new_n767), .A3(new_n573), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n754), .A2(new_n759), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT109), .B1(new_n755), .B2(new_n757), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT109), .ZN(new_n934));
  AOI211_X1 g0734(.A(new_n934), .B(KEYINPUT31), .C1(new_n754), .C2(new_n702), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n932), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(KEYINPUT110), .B1(new_n931), .B2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n932), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n934), .B1(new_n750), .B2(KEYINPUT31), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n755), .A2(KEYINPUT109), .A3(new_n757), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT110), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n941), .A2(new_n942), .A3(new_n768), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n930), .B1(new_n937), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT40), .B1(new_n944), .B2(new_n901), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT40), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n922), .B2(new_n900), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n945), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n457), .B1(new_n943), .B2(new_n937), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n738), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n948), .B2(new_n949), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n884), .B1(new_n929), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n929), .B2(new_n951), .ZN(new_n953));
  INV_X1    g0753(.A(new_n472), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n954), .A2(KEYINPUT35), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(KEYINPUT35), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n955), .A2(G116), .A3(new_n220), .A4(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT36), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n410), .A2(G77), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n250), .B1(new_n835), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n960), .A2(G1), .A3(new_n772), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n953), .A2(new_n958), .A3(new_n961), .ZN(G367));
  OAI211_X1 g0762(.A(new_n525), .B(new_n527), .C1(new_n480), .C2(new_n712), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n520), .A2(new_n702), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n718), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n969), .A2(KEYINPUT42), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT111), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n527), .B1(new_n963), .B2(new_n618), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n969), .A2(KEYINPUT42), .B1(new_n972), .B2(new_n712), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n712), .B1(new_n567), .B2(new_n569), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n975), .A2(new_n663), .ZN(new_n976));
  INV_X1    g0776(.A(new_n662), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT43), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n979), .A2(KEYINPUT43), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n974), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n971), .A2(new_n981), .A3(new_n980), .A4(new_n973), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n716), .A2(new_n966), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n986), .B(new_n987), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n725), .B(KEYINPUT41), .Z(new_n989));
  NAND2_X1  g0789(.A1(new_n719), .A2(new_n965), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT45), .Z(new_n991));
  NOR2_X1   g0791(.A1(new_n719), .A2(new_n965), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT44), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(new_n716), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n714), .A2(new_n717), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n967), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT112), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n997), .B1(new_n708), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n998), .B2(new_n708), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n709), .A2(KEYINPUT112), .A3(new_n997), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n995), .A2(new_n1002), .A3(new_n770), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n989), .B1(new_n1003), .B2(new_n770), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n988), .B1(new_n1004), .B2(new_n775), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n779), .B(new_n843), .C1(new_n721), .C2(new_n555), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n834), .A2(new_n245), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n831), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT46), .ZN(new_n1009));
  NOR3_X1   g0809(.A1(new_n781), .A2(new_n1009), .A3(new_n626), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1009), .B1(new_n781), .B2(new_n626), .ZN(new_n1011));
  INV_X1    g0811(.A(G317), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1011), .B1(new_n789), .B2(new_n1012), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1010), .B(new_n1013), .C1(G283), .C2(new_n799), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n258), .B1(new_n812), .B2(G107), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n801), .A2(G97), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1015), .B(new_n1016), .C1(new_n814), .C2(new_n819), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(G311), .B2(new_n794), .ZN(new_n1018));
  INV_X1    g0818(.A(G303), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1014), .B(new_n1018), .C1(new_n1019), .C2(new_n808), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n808), .A2(new_n326), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n790), .A2(G137), .B1(G50), .B2(new_n799), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n267), .B1(new_n801), .B2(G77), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n818), .A2(new_n202), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G58), .B2(new_n782), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G143), .A2(new_n794), .B1(new_n825), .B2(G159), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1022), .A2(new_n1023), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1020), .B1(new_n1021), .B2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT47), .Z(new_n1029));
  INV_X1    g0829(.A(new_n779), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1008), .B1(new_n847), .B2(new_n979), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1005), .A2(new_n1031), .ZN(G387));
  OAI21_X1  g0832(.A(KEYINPUT116), .B1(new_n1002), .B2(new_n770), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n725), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n1002), .B2(new_n770), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n770), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT116), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1000), .A2(new_n1036), .A3(new_n1037), .A4(new_n1001), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1033), .A2(new_n1035), .A3(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n832), .A2(new_n726), .B1(new_n351), .B2(new_n721), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n242), .A2(KEYINPUT113), .A3(G45), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n834), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n328), .A2(G50), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT50), .ZN(new_n1044));
  AOI211_X1 g0844(.A(G45), .B(new_n726), .C1(G68), .C2(G77), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1042), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT114), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1041), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(KEYINPUT113), .B1(new_n242), .B2(G45), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1040), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n831), .B1(new_n1050), .B2(new_n844), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n715), .B2(new_n847), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n790), .A2(G150), .B1(G68), .B2(new_n799), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n818), .A2(new_n360), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G77), .B2(new_n782), .ZN(new_n1055));
  AND4_X1   g0855(.A1(new_n258), .A2(new_n1053), .A3(new_n1016), .A4(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n329), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G159), .A2(new_n794), .B1(new_n1057), .B2(new_n825), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1056), .B(new_n1058), .C1(new_n207), .C2(new_n808), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n825), .A2(G311), .B1(new_n799), .B2(G303), .ZN(new_n1060));
  INV_X1    g0860(.A(G322), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1060), .B1(new_n795), .B2(new_n1061), .C1(new_n1012), .C2(new_n808), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT115), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT48), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n782), .A2(G294), .B1(new_n812), .B2(G283), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT49), .Z(new_n1069));
  NAND2_X1  g0869(.A1(new_n790), .A2(G326), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n258), .B1(new_n801), .B2(G116), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1059), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1052), .B1(new_n1073), .B2(new_n779), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n1002), .B2(new_n775), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1039), .A2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1076), .A2(KEYINPUT117), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1076), .A2(KEYINPUT117), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(G393));
  INV_X1    g0880(.A(new_n995), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n774), .B1(new_n1081), .B2(KEYINPUT118), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(KEYINPUT118), .B2(new_n1081), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1042), .A2(new_n249), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n779), .B(new_n843), .C1(G97), .C2(new_n721), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n831), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n809), .A2(G311), .B1(G317), .B2(new_n794), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT52), .Z(new_n1088));
  AOI22_X1  g0888(.A1(new_n782), .A2(G283), .B1(new_n812), .B2(G116), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1089), .B(new_n267), .C1(new_n351), .C2(new_n800), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n789), .A2(new_n1061), .B1(new_n819), .B2(new_n798), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1090), .B(new_n1091), .C1(G303), .C2(new_n825), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n407), .A2(new_n808), .B1(new_n795), .B2(new_n326), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT51), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n862), .A2(new_n267), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n812), .A2(G77), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1095), .B(new_n1096), .C1(new_n202), .C2(new_n781), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n789), .A2(new_n868), .B1(new_n328), .B2(new_n798), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n1097), .B(new_n1098), .C1(G50), .C2(new_n825), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1088), .A2(new_n1092), .B1(new_n1094), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n843), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n1086), .B1(new_n1100), .B2(new_n1030), .C1(new_n1101), .C2(new_n965), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1083), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1003), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n995), .B1(new_n770), .B2(new_n1002), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n1104), .A2(new_n1105), .A3(new_n1034), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(G390));
  AND3_X1   g0908(.A1(new_n941), .A2(new_n942), .A3(new_n768), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n942), .B1(new_n941), .B2(new_n768), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n456), .B(G330), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1111), .A2(new_n928), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n910), .A2(new_n855), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1113), .B(G330), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n765), .A2(new_n768), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1115), .A2(G330), .A3(new_n855), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n910), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1114), .A2(new_n1118), .B1(new_n904), .B2(new_n903), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1115), .A2(G330), .A3(new_n855), .A4(new_n910), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n854), .A2(new_n371), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n712), .B(new_n1121), .C1(new_n672), .C2(new_n732), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n904), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1120), .A2(new_n1124), .ZN(new_n1125));
  OAI211_X1 g0925(.A(G330), .B(new_n855), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1125), .B1(new_n1117), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1112), .B1(new_n1119), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1114), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n925), .B1(new_n905), .B2(new_n910), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT39), .ZN(new_n1131));
  AND4_X1   g0931(.A1(KEYINPUT38), .A2(new_n899), .A3(new_n895), .A4(new_n890), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n916), .A2(new_n918), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n431), .A2(new_n888), .A3(KEYINPUT37), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1133), .A2(new_n1134), .B1(new_n886), .B2(new_n894), .ZN(new_n1135));
  AOI21_X1  g0935(.A(KEYINPUT38), .B1(new_n1135), .B2(new_n899), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1131), .B1(new_n1132), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n898), .A2(KEYINPUT39), .A3(new_n900), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1130), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1123), .A2(new_n910), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n922), .A2(new_n900), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n925), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1129), .B1(new_n1139), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n911), .A2(new_n1142), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n914), .B2(new_n923), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1147), .A2(new_n1143), .A3(new_n1120), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1128), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n905), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1126), .A2(new_n1117), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1125), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1156), .A2(new_n1148), .A3(new_n1145), .A4(new_n1112), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1150), .A2(new_n725), .A3(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1145), .A2(new_n1148), .A3(new_n775), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n782), .A2(G150), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT53), .ZN(new_n1161));
  INV_X1    g0961(.A(G128), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n795), .A2(new_n1162), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1161), .B(new_n1163), .C1(G137), .C2(new_n825), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT54), .B(G143), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n798), .A2(new_n1165), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n258), .B1(new_n800), .B2(new_n207), .C1(new_n818), .C2(new_n407), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(G125), .C2(new_n790), .ZN(new_n1168));
  INV_X1    g0968(.A(G132), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1164), .B(new_n1168), .C1(new_n1169), .C2(new_n808), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1096), .B1(new_n202), .B2(new_n800), .C1(new_n789), .C2(new_n819), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G97), .B2(new_n799), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n267), .B1(new_n781), .B2(new_n226), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT119), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(G283), .A2(new_n794), .B1(new_n825), .B2(G107), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n809), .A2(G116), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1172), .A2(new_n1174), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1030), .B1(new_n1170), .B2(new_n1177), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n831), .B(new_n1178), .C1(new_n329), .C2(new_n879), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n924), .B2(new_n842), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1158), .A2(new_n1159), .A3(new_n1180), .ZN(G378));
  INV_X1    g0981(.A(new_n693), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n335), .A2(new_n887), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n1182), .A2(new_n347), .A3(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1183), .B1(new_n1182), .B2(new_n347), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  OR3_X1    g0987(.A1(new_n1184), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1187), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n841), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n258), .A2(G41), .ZN(new_n1193));
  AOI211_X1 g0993(.A(G50), .B(new_n1193), .C1(new_n263), .C2(new_n272), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n789), .A2(new_n820), .B1(new_n360), .B2(new_n798), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1193), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n801), .A2(G58), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n337), .B2(new_n781), .ZN(new_n1198));
  NOR4_X1   g0998(.A1(new_n1195), .A2(new_n1024), .A3(new_n1196), .A4(new_n1198), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G116), .A2(new_n794), .B1(new_n825), .B2(G97), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(new_n351), .C2(new_n808), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT58), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1194), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n818), .A2(new_n326), .B1(new_n781), .B2(new_n1165), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n799), .A2(G137), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1204), .B(new_n1205), .C1(G125), .C2(new_n794), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n1162), .B2(new_n808), .C1(new_n1169), .C2(new_n814), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(KEYINPUT59), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n790), .A2(G124), .ZN(new_n1209));
  AOI211_X1 g1009(.A(G33), .B(G41), .C1(new_n801), .C2(G159), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1207), .A2(KEYINPUT59), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1203), .B1(new_n1202), .B2(new_n1201), .C1(new_n1211), .C2(new_n1212), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1213), .A2(new_n779), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n831), .B(new_n1214), .C1(new_n207), .C2(new_n879), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1192), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT120), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1113), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n947), .ZN(new_n1219));
  OAI21_X1  g1019(.A(G330), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1217), .B1(new_n1220), .B2(new_n945), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n946), .B1(new_n1218), .B2(new_n902), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n738), .B1(new_n944), .B2(new_n947), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1222), .A2(new_n1223), .A3(KEYINPUT120), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1221), .A2(new_n1224), .A3(new_n1190), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1191), .A2(KEYINPUT120), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n927), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1225), .A2(new_n926), .A3(new_n913), .A4(new_n1226), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1216), .B1(new_n1230), .B2(new_n774), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT121), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n1157), .B2(new_n1112), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1127), .A2(new_n1119), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1232), .B(new_n1112), .C1(new_n1149), .C2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1229), .B(new_n1228), .C1(new_n1233), .C2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT57), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1034), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1112), .B1(new_n1149), .B2(new_n1234), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(KEYINPUT121), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1235), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1242), .A2(KEYINPUT57), .A3(new_n1229), .A4(new_n1228), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1231), .B1(new_n1239), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(G375));
  NAND2_X1  g1045(.A1(new_n1111), .A2(new_n928), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1234), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n989), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(new_n1128), .A3(new_n1248), .ZN(new_n1249));
  XOR2_X1   g1049(.A(new_n1249), .B(KEYINPUT122), .Z(new_n1250));
  XOR2_X1   g1050(.A(new_n774), .B(KEYINPUT123), .Z(new_n1251));
  NOR2_X1   g1051(.A1(new_n910), .A2(new_n842), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n795), .A2(new_n819), .B1(new_n626), .B2(new_n814), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n267), .B1(new_n800), .B2(new_n337), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1254), .B(new_n1054), .C1(G97), .C2(new_n782), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1255), .B1(new_n351), .B2(new_n798), .C1(new_n1019), .C2(new_n789), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1253), .B(new_n1256), .C1(G283), .C2(new_n809), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n795), .A2(new_n1169), .B1(new_n814), .B2(new_n1165), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n790), .A2(G128), .B1(G150), .B2(new_n799), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n782), .A2(G159), .B1(new_n812), .B2(G50), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1259), .A2(new_n258), .A3(new_n1197), .A4(new_n1260), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n1258), .B(new_n1261), .C1(G137), .C2(new_n809), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n779), .B1(new_n1257), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n879), .A2(new_n202), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1263), .A2(new_n776), .A3(new_n1264), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n1234), .A2(new_n1251), .B1(new_n1252), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1250), .A2(new_n1267), .ZN(G381));
  NOR2_X1   g1068(.A1(G375), .A2(G378), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1078), .A2(new_n850), .A3(new_n1079), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT124), .ZN(new_n1271));
  OR3_X1    g1071(.A1(new_n1270), .A2(new_n1271), .A3(G384), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1271), .B1(new_n1270), .B2(G384), .ZN(new_n1273));
  NOR3_X1   g1073(.A1(G390), .A2(G381), .A3(G387), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1269), .A2(new_n1272), .A3(new_n1273), .A4(new_n1274), .ZN(G407));
  NAND2_X1  g1075(.A1(new_n1269), .A2(new_n701), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(G407), .A2(G213), .A3(new_n1276), .ZN(G409));
  NAND2_X1  g1077(.A1(new_n1128), .A2(KEYINPUT60), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1034), .B1(new_n1278), .B2(new_n1247), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT125), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1234), .A2(KEYINPUT60), .A3(new_n1246), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1246), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT60), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1247), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1285), .A2(new_n1281), .A3(new_n725), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(KEYINPUT125), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1282), .A2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(G384), .B1(new_n1288), .B2(new_n1267), .ZN(new_n1289));
  AOI211_X1 g1089(.A(new_n882), .B(new_n1266), .C1(new_n1282), .C2(new_n1287), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(G213), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1292), .A2(G343), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(G378), .ZN(new_n1295));
  AOI211_X1 g1095(.A(new_n1295), .B(new_n1231), .C1(new_n1239), .C2(new_n1243), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n989), .B1(new_n1241), .B2(new_n1235), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1251), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1229), .B(new_n1228), .C1(new_n1297), .C2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(G378), .B1(new_n1299), .B2(new_n1216), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1291), .B(new_n1294), .C1(new_n1296), .C2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(KEYINPUT62), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT61), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1288), .A2(new_n1267), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n882), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1288), .A2(G384), .A3(new_n1267), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1293), .A2(G2897), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1305), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1307), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1309), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1300), .B1(new_n1244), .B2(G378), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1308), .B(new_n1310), .C1(new_n1311), .C2(new_n1293), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1313), .A2(new_n725), .A3(new_n1243), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1231), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1314), .A2(G378), .A3(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1300), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT62), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1318), .A2(new_n1319), .A3(new_n1291), .A4(new_n1294), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1302), .A2(new_n1303), .A3(new_n1312), .A4(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1079), .ZN(new_n1322));
  OAI21_X1  g1122(.A(G396), .B1(new_n1322), .B2(new_n1077), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1323), .A2(new_n1270), .A3(G387), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT126), .ZN(new_n1326));
  AOI22_X1  g1126(.A1(new_n1270), .A2(new_n1323), .B1(G387), .B2(new_n1326), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1107), .B1(new_n1325), .B2(new_n1327), .ZN(new_n1328));
  AND2_X1   g1128(.A1(new_n1323), .A2(new_n1270), .ZN(new_n1329));
  AOI21_X1  g1129(.A(KEYINPUT126), .B1(new_n1005), .B2(new_n1031), .ZN(new_n1330));
  OAI211_X1 g1130(.A(G390), .B(new_n1324), .C1(new_n1329), .C2(new_n1330), .ZN(new_n1331));
  AND2_X1   g1131(.A1(new_n1328), .A2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1321), .A2(new_n1332), .ZN(new_n1333));
  AND2_X1   g1133(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1318), .A2(new_n1294), .ZN(new_n1335));
  AOI21_X1  g1135(.A(KEYINPUT61), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT63), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1301), .A2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1328), .A2(new_n1331), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1318), .A2(KEYINPUT63), .A3(new_n1291), .A4(new_n1294), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1336), .A2(new_n1338), .A3(new_n1339), .A4(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1333), .A2(new_n1341), .ZN(G405));
  NOR2_X1   g1142(.A1(new_n1244), .A2(G378), .ZN(new_n1343));
  NOR2_X1   g1143(.A1(new_n1343), .A2(new_n1296), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1291), .A2(KEYINPUT127), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  OAI211_X1 g1146(.A(KEYINPUT127), .B(new_n1291), .C1(new_n1343), .C2(new_n1296), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  XNOR2_X1  g1148(.A(new_n1348), .B(new_n1332), .ZN(G402));
endmodule


