

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U324 ( .A(n300), .B(n299), .ZN(n314) );
  XNOR2_X1 U325 ( .A(n478), .B(n477), .ZN(n499) );
  XNOR2_X1 U326 ( .A(n309), .B(n308), .ZN(n526) );
  XNOR2_X1 U327 ( .A(n443), .B(n323), .ZN(n517) );
  XOR2_X1 U328 ( .A(n383), .B(n382), .Z(n292) );
  INV_X1 U329 ( .A(KEYINPUT98), .ZN(n463) );
  XNOR2_X1 U330 ( .A(n298), .B(G183GAT), .ZN(n299) );
  XNOR2_X1 U331 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n405) );
  INV_X1 U332 ( .A(KEYINPUT94), .ZN(n315) );
  XNOR2_X1 U333 ( .A(n406), .B(n405), .ZN(n565) );
  OR2_X1 U334 ( .A1(n581), .A2(n576), .ZN(n474) );
  XNOR2_X1 U335 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U336 ( .A(n384), .B(n292), .ZN(n385) );
  OR2_X1 U337 ( .A1(n484), .A2(n474), .ZN(n475) );
  XNOR2_X1 U338 ( .A(n318), .B(n317), .ZN(n322) );
  XNOR2_X1 U339 ( .A(n386), .B(n385), .ZN(n387) );
  NOR2_X1 U340 ( .A1(n526), .A2(n449), .ZN(n561) );
  INV_X1 U341 ( .A(G43GAT), .ZN(n479) );
  XNOR2_X1 U342 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U343 ( .A(n479), .B(KEYINPUT40), .ZN(n480) );
  XNOR2_X1 U344 ( .A(n456), .B(n455), .ZN(G1351GAT) );
  XNOR2_X1 U345 ( .A(n481), .B(n480), .ZN(G1330GAT) );
  XOR2_X1 U346 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n294) );
  NAND2_X1 U347 ( .A1(G227GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U348 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U349 ( .A(n295), .B(KEYINPUT84), .Z(n305) );
  XOR2_X1 U350 ( .A(KEYINPUT83), .B(KEYINPUT19), .Z(n297) );
  XNOR2_X1 U351 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n296) );
  XNOR2_X1 U352 ( .A(n297), .B(n296), .ZN(n300) );
  XOR2_X1 U353 ( .A(G169GAT), .B(G176GAT), .Z(n298) );
  XOR2_X1 U354 ( .A(G99GAT), .B(G134GAT), .Z(n302) );
  XNOR2_X1 U355 ( .A(G43GAT), .B(G190GAT), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U357 ( .A(n314), .B(n303), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n305), .B(n304), .ZN(n307) );
  XNOR2_X1 U359 ( .A(G127GAT), .B(KEYINPUT82), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n306), .B(KEYINPUT0), .ZN(n415) );
  XOR2_X1 U361 ( .A(n307), .B(n415), .Z(n309) );
  XOR2_X1 U362 ( .A(G113GAT), .B(G15GAT), .Z(n362) );
  XOR2_X1 U363 ( .A(G120GAT), .B(G71GAT), .Z(n381) );
  XNOR2_X1 U364 ( .A(n362), .B(n381), .ZN(n308) );
  XOR2_X1 U365 ( .A(KEYINPUT88), .B(G204GAT), .Z(n311) );
  XNOR2_X1 U366 ( .A(G197GAT), .B(G211GAT), .ZN(n310) );
  XNOR2_X1 U367 ( .A(n311), .B(n310), .ZN(n313) );
  XOR2_X1 U368 ( .A(KEYINPUT21), .B(KEYINPUT87), .Z(n312) );
  XNOR2_X1 U369 ( .A(n313), .B(n312), .ZN(n443) );
  XOR2_X1 U370 ( .A(G8GAT), .B(G64GAT), .Z(n342) );
  XOR2_X1 U371 ( .A(n342), .B(n314), .Z(n318) );
  NAND2_X1 U372 ( .A1(G226GAT), .A2(G233GAT), .ZN(n316) );
  XOR2_X1 U373 ( .A(G92GAT), .B(G218GAT), .Z(n320) );
  XNOR2_X1 U374 ( .A(G36GAT), .B(G190GAT), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n333) );
  XNOR2_X1 U376 ( .A(n333), .B(KEYINPUT95), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U378 ( .A(n517), .B(KEYINPUT118), .Z(n404) );
  XOR2_X1 U379 ( .A(KEYINPUT9), .B(KEYINPUT74), .Z(n325) );
  XNOR2_X1 U380 ( .A(KEYINPUT76), .B(KEYINPUT66), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U382 ( .A(n326), .B(KEYINPUT10), .Z(n328) );
  XOR2_X1 U383 ( .A(G134GAT), .B(G162GAT), .Z(n416) );
  XNOR2_X1 U384 ( .A(n416), .B(KEYINPUT77), .ZN(n327) );
  XNOR2_X1 U385 ( .A(n328), .B(n327), .ZN(n337) );
  XOR2_X1 U386 ( .A(KEYINPUT11), .B(KEYINPUT75), .Z(n330) );
  NAND2_X1 U387 ( .A1(G232GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U389 ( .A(n331), .B(KEYINPUT78), .Z(n335) );
  XNOR2_X1 U390 ( .A(G99GAT), .B(G106GAT), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n332), .B(G85GAT), .ZN(n377) );
  XNOR2_X1 U392 ( .A(n333), .B(n377), .ZN(n334) );
  XNOR2_X1 U393 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U394 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U395 ( .A(KEYINPUT8), .B(G50GAT), .Z(n339) );
  XNOR2_X1 U396 ( .A(G43GAT), .B(G29GAT), .ZN(n338) );
  XNOR2_X1 U397 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U398 ( .A(KEYINPUT7), .B(n340), .ZN(n373) );
  XNOR2_X1 U399 ( .A(n341), .B(n373), .ZN(n555) );
  XOR2_X1 U400 ( .A(KEYINPUT13), .B(G57GAT), .Z(n380) );
  XOR2_X1 U401 ( .A(n342), .B(n380), .Z(n344) );
  XNOR2_X1 U402 ( .A(G22GAT), .B(G155GAT), .ZN(n343) );
  XNOR2_X1 U403 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U404 ( .A(KEYINPUT81), .B(KEYINPUT12), .Z(n346) );
  NAND2_X1 U405 ( .A1(G231GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U406 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U407 ( .A(n348), .B(n347), .Z(n350) );
  XOR2_X1 U408 ( .A(KEYINPUT69), .B(G1GAT), .Z(n361) );
  XNOR2_X1 U409 ( .A(n361), .B(KEYINPUT14), .ZN(n349) );
  XNOR2_X1 U410 ( .A(n350), .B(n349), .ZN(n358) );
  XOR2_X1 U411 ( .A(G78GAT), .B(G211GAT), .Z(n352) );
  XNOR2_X1 U412 ( .A(G15GAT), .B(G71GAT), .ZN(n351) );
  XNOR2_X1 U413 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U414 ( .A(KEYINPUT80), .B(KEYINPUT15), .Z(n354) );
  XNOR2_X1 U415 ( .A(G183GAT), .B(G127GAT), .ZN(n353) );
  XNOR2_X1 U416 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U417 ( .A(n356), .B(n355), .Z(n357) );
  XNOR2_X1 U418 ( .A(n358), .B(n357), .ZN(n576) );
  XOR2_X1 U419 ( .A(KEYINPUT67), .B(KEYINPUT29), .Z(n360) );
  XNOR2_X1 U420 ( .A(G169GAT), .B(KEYINPUT30), .ZN(n359) );
  XNOR2_X1 U421 ( .A(n360), .B(n359), .ZN(n372) );
  XOR2_X1 U422 ( .A(G197GAT), .B(G36GAT), .Z(n364) );
  XNOR2_X1 U423 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U424 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U425 ( .A(G141GAT), .B(G22GAT), .Z(n431) );
  XOR2_X1 U426 ( .A(n365), .B(n431), .Z(n370) );
  XOR2_X1 U427 ( .A(KEYINPUT70), .B(G8GAT), .Z(n367) );
  NAND2_X1 U428 ( .A1(G229GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U430 ( .A(KEYINPUT68), .B(n368), .ZN(n369) );
  XNOR2_X1 U431 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U432 ( .A(n372), .B(n371), .ZN(n374) );
  XNOR2_X1 U433 ( .A(n374), .B(n373), .ZN(n569) );
  XOR2_X1 U434 ( .A(KEYINPUT33), .B(G92GAT), .Z(n376) );
  XNOR2_X1 U435 ( .A(G176GAT), .B(G204GAT), .ZN(n375) );
  XNOR2_X1 U436 ( .A(n376), .B(n375), .ZN(n388) );
  XOR2_X1 U437 ( .A(G148GAT), .B(G78GAT), .Z(n430) );
  XOR2_X1 U438 ( .A(n377), .B(n430), .Z(n379) );
  NAND2_X1 U439 ( .A1(G230GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U440 ( .A(n379), .B(n378), .ZN(n386) );
  XNOR2_X1 U441 ( .A(n381), .B(n380), .ZN(n384) );
  XOR2_X1 U442 ( .A(KEYINPUT72), .B(KEYINPUT31), .Z(n383) );
  XNOR2_X1 U443 ( .A(G64GAT), .B(KEYINPUT32), .ZN(n382) );
  XOR2_X1 U444 ( .A(n388), .B(n387), .Z(n573) );
  XOR2_X1 U445 ( .A(KEYINPUT41), .B(KEYINPUT65), .Z(n389) );
  XNOR2_X1 U446 ( .A(n573), .B(n389), .ZN(n545) );
  NOR2_X1 U447 ( .A1(n569), .A2(n545), .ZN(n390) );
  XNOR2_X1 U448 ( .A(n390), .B(KEYINPUT46), .ZN(n391) );
  NOR2_X1 U449 ( .A1(n576), .A2(n391), .ZN(n392) );
  NAND2_X1 U450 ( .A1(n555), .A2(n392), .ZN(n393) );
  XNOR2_X1 U451 ( .A(n393), .B(KEYINPUT47), .ZN(n394) );
  XNOR2_X1 U452 ( .A(n394), .B(KEYINPUT109), .ZN(n401) );
  INV_X1 U453 ( .A(n576), .ZN(n551) );
  XNOR2_X1 U454 ( .A(KEYINPUT79), .B(n555), .ZN(n538) );
  XNOR2_X1 U455 ( .A(KEYINPUT36), .B(KEYINPUT101), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n538), .B(n395), .ZN(n581) );
  NOR2_X1 U457 ( .A1(n551), .A2(n581), .ZN(n396) );
  XOR2_X1 U458 ( .A(n396), .B(KEYINPUT45), .Z(n397) );
  XNOR2_X1 U459 ( .A(KEYINPUT110), .B(n397), .ZN(n398) );
  NOR2_X1 U460 ( .A1(n573), .A2(n398), .ZN(n399) );
  XNOR2_X1 U461 ( .A(KEYINPUT71), .B(n569), .ZN(n558) );
  INV_X1 U462 ( .A(n558), .ZN(n529) );
  NAND2_X1 U463 ( .A1(n399), .A2(n529), .ZN(n400) );
  NAND2_X1 U464 ( .A1(n401), .A2(n400), .ZN(n403) );
  XNOR2_X1 U465 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n402) );
  XNOR2_X1 U466 ( .A(n403), .B(n402), .ZN(n524) );
  NAND2_X1 U467 ( .A1(n404), .A2(n524), .ZN(n406) );
  XOR2_X1 U468 ( .A(KEYINPUT1), .B(KEYINPUT93), .Z(n408) );
  XNOR2_X1 U469 ( .A(KEYINPUT92), .B(KEYINPUT6), .ZN(n407) );
  XNOR2_X1 U470 ( .A(n408), .B(n407), .ZN(n427) );
  XOR2_X1 U471 ( .A(G57GAT), .B(G120GAT), .Z(n410) );
  XNOR2_X1 U472 ( .A(G113GAT), .B(G1GAT), .ZN(n409) );
  XNOR2_X1 U473 ( .A(n410), .B(n409), .ZN(n414) );
  XOR2_X1 U474 ( .A(G85GAT), .B(G148GAT), .Z(n412) );
  XNOR2_X1 U475 ( .A(G29GAT), .B(G141GAT), .ZN(n411) );
  XNOR2_X1 U476 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U477 ( .A(n414), .B(n413), .ZN(n425) );
  XOR2_X1 U478 ( .A(n416), .B(n415), .Z(n418) );
  NAND2_X1 U479 ( .A1(G225GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U481 ( .A(n419), .B(KEYINPUT4), .Z(n423) );
  XOR2_X1 U482 ( .A(G155GAT), .B(KEYINPUT89), .Z(n421) );
  XNOR2_X1 U483 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n421), .B(n420), .ZN(n435) );
  XNOR2_X1 U485 ( .A(n435), .B(KEYINPUT5), .ZN(n422) );
  XNOR2_X1 U486 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U488 ( .A(n427), .B(n426), .ZN(n564) );
  XOR2_X1 U489 ( .A(KEYINPUT91), .B(KEYINPUT23), .Z(n429) );
  XNOR2_X1 U490 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n429), .B(n428), .ZN(n442) );
  XOR2_X1 U492 ( .A(G106GAT), .B(G162GAT), .Z(n433) );
  XNOR2_X1 U493 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U494 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U495 ( .A(n434), .B(G218GAT), .Z(n440) );
  XOR2_X1 U496 ( .A(n435), .B(KEYINPUT90), .Z(n437) );
  NAND2_X1 U497 ( .A1(G228GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U498 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U499 ( .A(G50GAT), .B(n438), .ZN(n439) );
  XNOR2_X1 U500 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U501 ( .A(n442), .B(n441), .ZN(n444) );
  XNOR2_X1 U502 ( .A(n444), .B(n443), .ZN(n467) );
  INV_X1 U503 ( .A(n467), .ZN(n445) );
  AND2_X1 U504 ( .A1(n564), .A2(n445), .ZN(n446) );
  AND2_X1 U505 ( .A1(n565), .A2(n446), .ZN(n448) );
  XNOR2_X1 U506 ( .A(KEYINPUT120), .B(KEYINPUT55), .ZN(n447) );
  XNOR2_X1 U507 ( .A(n448), .B(n447), .ZN(n449) );
  INV_X1 U508 ( .A(n545), .ZN(n501) );
  NAND2_X1 U509 ( .A1(n561), .A2(n501), .ZN(n452) );
  XOR2_X1 U510 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n450) );
  XNOR2_X1 U511 ( .A(n450), .B(G176GAT), .ZN(n451) );
  XNOR2_X1 U512 ( .A(n452), .B(n451), .ZN(G1349GAT) );
  NAND2_X1 U513 ( .A1(n561), .A2(n538), .ZN(n456) );
  XOR2_X1 U514 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n454) );
  XNOR2_X1 U515 ( .A(G190GAT), .B(KEYINPUT123), .ZN(n453) );
  NOR2_X1 U516 ( .A1(n526), .A2(n517), .ZN(n457) );
  NOR2_X1 U517 ( .A1(n467), .A2(n457), .ZN(n458) );
  XOR2_X1 U518 ( .A(KEYINPUT25), .B(n458), .Z(n462) );
  XOR2_X1 U519 ( .A(KEYINPUT97), .B(KEYINPUT26), .Z(n460) );
  NAND2_X1 U520 ( .A1(n526), .A2(n467), .ZN(n459) );
  XNOR2_X1 U521 ( .A(n460), .B(n459), .ZN(n566) );
  XNOR2_X1 U522 ( .A(KEYINPUT27), .B(n517), .ZN(n468) );
  NOR2_X1 U523 ( .A1(n566), .A2(n468), .ZN(n461) );
  NOR2_X1 U524 ( .A1(n462), .A2(n461), .ZN(n464) );
  XNOR2_X1 U525 ( .A(n464), .B(n463), .ZN(n465) );
  NAND2_X1 U526 ( .A1(n465), .A2(n564), .ZN(n466) );
  XNOR2_X1 U527 ( .A(KEYINPUT99), .B(n466), .ZN(n473) );
  XNOR2_X1 U528 ( .A(KEYINPUT28), .B(n467), .ZN(n492) );
  XNOR2_X1 U529 ( .A(n526), .B(KEYINPUT86), .ZN(n469) );
  NOR2_X1 U530 ( .A1(n564), .A2(n468), .ZN(n525) );
  NAND2_X1 U531 ( .A1(n469), .A2(n525), .ZN(n470) );
  NOR2_X1 U532 ( .A1(n492), .A2(n470), .ZN(n471) );
  XNOR2_X1 U533 ( .A(n471), .B(KEYINPUT96), .ZN(n472) );
  NOR2_X1 U534 ( .A1(n473), .A2(n472), .ZN(n484) );
  XNOR2_X1 U535 ( .A(KEYINPUT37), .B(n475), .ZN(n514) );
  NOR2_X1 U536 ( .A1(n573), .A2(n529), .ZN(n476) );
  XOR2_X1 U537 ( .A(KEYINPUT73), .B(n476), .Z(n486) );
  NAND2_X1 U538 ( .A1(n514), .A2(n486), .ZN(n478) );
  XNOR2_X1 U539 ( .A(KEYINPUT38), .B(KEYINPUT102), .ZN(n477) );
  NOR2_X1 U540 ( .A1(n526), .A2(n499), .ZN(n481) );
  NOR2_X1 U541 ( .A1(n551), .A2(n538), .ZN(n482) );
  XOR2_X1 U542 ( .A(KEYINPUT16), .B(n482), .Z(n483) );
  NOR2_X1 U543 ( .A1(n484), .A2(n483), .ZN(n485) );
  XNOR2_X1 U544 ( .A(KEYINPUT100), .B(n485), .ZN(n502) );
  NAND2_X1 U545 ( .A1(n486), .A2(n502), .ZN(n493) );
  NOR2_X1 U546 ( .A1(n564), .A2(n493), .ZN(n487) );
  XOR2_X1 U547 ( .A(n487), .B(KEYINPUT34), .Z(n488) );
  XNOR2_X1 U548 ( .A(G1GAT), .B(n488), .ZN(G1324GAT) );
  NOR2_X1 U549 ( .A1(n517), .A2(n493), .ZN(n489) );
  XOR2_X1 U550 ( .A(G8GAT), .B(n489), .Z(G1325GAT) );
  NOR2_X1 U551 ( .A1(n526), .A2(n493), .ZN(n491) );
  XNOR2_X1 U552 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(G1326GAT) );
  INV_X1 U554 ( .A(n492), .ZN(n527) );
  NOR2_X1 U555 ( .A1(n527), .A2(n493), .ZN(n494) );
  XOR2_X1 U556 ( .A(G22GAT), .B(n494), .Z(G1327GAT) );
  NOR2_X1 U557 ( .A1(n499), .A2(n564), .ZN(n496) );
  XNOR2_X1 U558 ( .A(KEYINPUT39), .B(KEYINPUT103), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U560 ( .A(G29GAT), .B(n497), .Z(G1328GAT) );
  NOR2_X1 U561 ( .A1(n517), .A2(n499), .ZN(n498) );
  XOR2_X1 U562 ( .A(G36GAT), .B(n498), .Z(G1329GAT) );
  NOR2_X1 U563 ( .A1(n527), .A2(n499), .ZN(n500) );
  XOR2_X1 U564 ( .A(G50GAT), .B(n500), .Z(G1331GAT) );
  AND2_X1 U565 ( .A1(n501), .A2(n569), .ZN(n513) );
  NAND2_X1 U566 ( .A1(n502), .A2(n513), .ZN(n503) );
  XNOR2_X1 U567 ( .A(KEYINPUT104), .B(n503), .ZN(n509) );
  NOR2_X1 U568 ( .A1(n509), .A2(n564), .ZN(n505) );
  XNOR2_X1 U569 ( .A(KEYINPUT42), .B(KEYINPUT105), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U571 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  NOR2_X1 U572 ( .A1(n517), .A2(n509), .ZN(n507) );
  XOR2_X1 U573 ( .A(G64GAT), .B(n507), .Z(G1333GAT) );
  NOR2_X1 U574 ( .A1(n526), .A2(n509), .ZN(n508) );
  XOR2_X1 U575 ( .A(G71GAT), .B(n508), .Z(G1334GAT) );
  NOR2_X1 U576 ( .A1(n509), .A2(n527), .ZN(n511) );
  XNOR2_X1 U577 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(n512), .ZN(G1335GAT) );
  NAND2_X1 U580 ( .A1(n514), .A2(n513), .ZN(n521) );
  NOR2_X1 U581 ( .A1(n564), .A2(n521), .ZN(n516) );
  XNOR2_X1 U582 ( .A(G85GAT), .B(KEYINPUT107), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n516), .B(n515), .ZN(G1336GAT) );
  NOR2_X1 U584 ( .A1(n517), .A2(n521), .ZN(n518) );
  XOR2_X1 U585 ( .A(KEYINPUT108), .B(n518), .Z(n519) );
  XNOR2_X1 U586 ( .A(G92GAT), .B(n519), .ZN(G1337GAT) );
  NOR2_X1 U587 ( .A1(n526), .A2(n521), .ZN(n520) );
  XOR2_X1 U588 ( .A(G99GAT), .B(n520), .Z(G1338GAT) );
  NOR2_X1 U589 ( .A1(n527), .A2(n521), .ZN(n522) );
  XOR2_X1 U590 ( .A(KEYINPUT44), .B(n522), .Z(n523) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  NAND2_X1 U592 ( .A1(n525), .A2(n524), .ZN(n543) );
  NOR2_X1 U593 ( .A1(n526), .A2(n543), .ZN(n528) );
  NAND2_X1 U594 ( .A1(n528), .A2(n527), .ZN(n537) );
  NOR2_X1 U595 ( .A1(n529), .A2(n537), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n530), .B(KEYINPUT111), .ZN(n531) );
  XNOR2_X1 U597 ( .A(G113GAT), .B(n531), .ZN(G1340GAT) );
  NOR2_X1 U598 ( .A1(n545), .A2(n537), .ZN(n533) );
  XNOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  NOR2_X1 U601 ( .A1(n551), .A2(n537), .ZN(n535) );
  XNOR2_X1 U602 ( .A(KEYINPUT50), .B(KEYINPUT112), .ZN(n534) );
  XNOR2_X1 U603 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U604 ( .A(G127GAT), .B(n536), .Z(G1342GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n541) );
  INV_X1 U606 ( .A(n537), .ZN(n539) );
  NAND2_X1 U607 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U609 ( .A(G134GAT), .B(n542), .Z(G1343GAT) );
  OR2_X1 U610 ( .A1(n566), .A2(n543), .ZN(n554) );
  NOR2_X1 U611 ( .A1(n569), .A2(n554), .ZN(n544) );
  XOR2_X1 U612 ( .A(G141GAT), .B(n544), .Z(G1344GAT) );
  NOR2_X1 U613 ( .A1(n545), .A2(n554), .ZN(n550) );
  XOR2_X1 U614 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n547) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n546) );
  XNOR2_X1 U616 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U617 ( .A(KEYINPUT53), .B(n548), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(G1345GAT) );
  NOR2_X1 U619 ( .A1(n551), .A2(n554), .ZN(n552) );
  XOR2_X1 U620 ( .A(KEYINPUT116), .B(n552), .Z(n553) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(n553), .ZN(G1346GAT) );
  NOR2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G162GAT), .B(KEYINPUT117), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1347GAT) );
  NAND2_X1 U625 ( .A1(n558), .A2(n561), .ZN(n560) );
  XOR2_X1 U626 ( .A(G169GAT), .B(KEYINPUT121), .Z(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1348GAT) );
  NAND2_X1 U628 ( .A1(n576), .A2(n561), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(KEYINPUT122), .ZN(n563) );
  XNOR2_X1 U630 ( .A(G183GAT), .B(n563), .ZN(G1350GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n567) );
  NOR2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(n568), .B(KEYINPUT125), .ZN(n582) );
  NOR2_X1 U634 ( .A1(n569), .A2(n582), .ZN(n571) );
  XNOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT61), .Z(n575) );
  INV_X1 U639 ( .A(n582), .ZN(n577) );
  NAND2_X1 U640 ( .A1(n577), .A2(n573), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(G1353GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n579) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(KEYINPUT62), .B(n583), .Z(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

