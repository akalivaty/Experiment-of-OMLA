//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1273,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n208));
  INV_X1    g0008(.A(G232), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n208), .B1(new_n202), .B2(new_n209), .C1(new_n203), .C2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n207), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT65), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT1), .ZN(new_n217));
  AND2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n216), .A2(new_n217), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT64), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g0022(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  NOR3_X1   g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n207), .A2(G13), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT0), .Z(new_n230));
  NOR4_X1   g0030(.A1(new_n218), .A2(new_n219), .A3(new_n227), .A4(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n209), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT66), .ZN(new_n243));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XOR2_X1   g0044(.A(G50), .B(G58), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  AND2_X1   g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NOR2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n250), .B1(G223), .B2(G1698), .ZN(new_n251));
  INV_X1    g0051(.A(G222), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT68), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n251), .B1(new_n252), .B2(new_n257), .ZN(new_n258));
  AND3_X1   g0058(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n259));
  AOI21_X1  g0059(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n260));
  AND2_X1   g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  OR2_X1    g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n258), .B(new_n262), .C1(G77), .C2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  INV_X1    g0067(.A(G41), .ZN(new_n268));
  INV_X1    g0068(.A(G45), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AND2_X1   g0070(.A1(G1), .A2(G13), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n267), .A2(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  XOR2_X1   g0073(.A(KEYINPUT67), .B(G226), .Z(new_n274));
  INV_X1    g0074(.A(G274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(new_n271), .B2(new_n272), .ZN(new_n276));
  AOI21_X1  g0076(.A(G1), .B1(new_n268), .B2(new_n269), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n273), .A2(new_n274), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n266), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G179), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n283), .B1(new_n259), .B2(new_n260), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT69), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT69), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n224), .A2(new_n286), .A3(new_n283), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n267), .A2(G13), .A3(G20), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n267), .A2(G20), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(G50), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G33), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT70), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT8), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G58), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n225), .A2(G33), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT70), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n296), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(G20), .A2(G33), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n288), .A2(new_n307), .B1(new_n201), .B2(new_n290), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n293), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G169), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n279), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n282), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n309), .A2(KEYINPUT9), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT9), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n293), .A2(new_n315), .A3(new_n308), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n314), .A2(new_n316), .B1(new_n280), .B2(G190), .ZN(new_n317));
  INV_X1    g0117(.A(G200), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n317), .A2(KEYINPUT75), .B1(new_n318), .B2(new_n280), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n317), .A2(KEYINPUT75), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT10), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n280), .A2(new_n318), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT74), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT10), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n324), .B(new_n317), .C1(new_n323), .C2(new_n322), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n313), .B1(new_n321), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n255), .A2(G226), .A3(new_n256), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n209), .A2(new_n254), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n250), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G97), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n294), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n262), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT13), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n273), .A2(G238), .B1(new_n276), .B2(new_n277), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n336), .B(KEYINPUT78), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT77), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n333), .A2(new_n335), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n338), .B1(new_n339), .B2(KEYINPUT13), .ZN(new_n340));
  AOI211_X1 g0140(.A(KEYINPUT77), .B(new_n334), .C1(new_n333), .C2(new_n335), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n337), .A2(new_n342), .A3(G190), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT72), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n289), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n267), .A2(KEYINPUT72), .A3(G13), .A4(G20), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n203), .A2(KEYINPUT12), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n347), .A2(new_n348), .B1(KEYINPUT12), .B2(new_n290), .ZN(new_n349));
  INV_X1    g0149(.A(new_n207), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n222), .A2(new_n223), .B1(new_n350), .B2(G33), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n347), .A2(new_n351), .A3(new_n292), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT12), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n349), .B1(new_n353), .B2(G68), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n296), .A2(G77), .A3(new_n303), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n305), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n288), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT11), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n288), .A2(KEYINPUT11), .A3(new_n357), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n354), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT79), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT79), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n354), .A2(new_n364), .A3(new_n360), .A4(new_n361), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n262), .ZN(new_n367));
  AND2_X1   g0167(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n368));
  NOR2_X1   g0168(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n369));
  INV_X1    g0169(.A(G226), .ZN(new_n370));
  NOR3_X1   g0170(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n265), .B1(new_n371), .B2(new_n328), .ZN(new_n372));
  INV_X1    g0172(.A(new_n332), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n367), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n335), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT13), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT76), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(new_n377), .A3(new_n336), .ZN(new_n378));
  OAI211_X1 g0178(.A(KEYINPUT76), .B(KEYINPUT13), .C1(new_n374), .C2(new_n375), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(G200), .A3(new_n379), .ZN(new_n380));
  AND3_X1   g0180(.A1(new_n343), .A2(new_n366), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n366), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n378), .A2(G169), .A3(new_n379), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT14), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n337), .A2(new_n342), .A3(G179), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT14), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n378), .A2(new_n386), .A3(G169), .A4(new_n379), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n381), .B1(new_n382), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n255), .A2(G223), .A3(new_n256), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G226), .A2(G1698), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n250), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G87), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n262), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n273), .A2(G232), .B1(new_n276), .B2(new_n277), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(new_n281), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT82), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n395), .A2(KEYINPUT82), .A3(new_n281), .A4(new_n396), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n395), .A2(new_n396), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n310), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n202), .A2(new_n203), .ZN(new_n404));
  NOR2_X1   g0204(.A1(G58), .A2(G68), .ZN(new_n405));
  OAI21_X1  g0205(.A(G20), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n305), .A2(G159), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n263), .A2(new_n225), .A3(new_n264), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT7), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n263), .A2(KEYINPUT7), .A3(new_n225), .A4(new_n264), .ZN(new_n413));
  AND3_X1   g0213(.A1(new_n412), .A2(KEYINPUT80), .A3(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(G68), .B1(new_n413), .B2(KEYINPUT80), .ZN(new_n415));
  OAI211_X1 g0215(.A(KEYINPUT16), .B(new_n409), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  XNOR2_X1  g0216(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n203), .B1(new_n412), .B2(new_n413), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n417), .B1(new_n418), .B2(new_n408), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n416), .A2(new_n284), .A3(new_n419), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n300), .A2(new_n292), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n285), .A2(new_n421), .A3(new_n287), .A4(new_n289), .ZN(new_n422));
  INV_X1    g0222(.A(new_n300), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n290), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT18), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n403), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT7), .B1(new_n250), .B2(new_n225), .ZN(new_n430));
  INV_X1    g0230(.A(new_n413), .ZN(new_n431));
  OAI21_X1  g0231(.A(G68), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n409), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n351), .B1(new_n433), .B2(new_n417), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n425), .B1(new_n434), .B2(new_n416), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT18), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n429), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT83), .ZN(new_n439));
  INV_X1    g0239(.A(G190), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n395), .A2(new_n440), .A3(new_n396), .ZN(new_n441));
  AOI21_X1  g0241(.A(G200), .B1(new_n395), .B2(new_n396), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n395), .A2(new_n440), .A3(new_n396), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n273), .A2(G232), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n276), .A2(new_n277), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n368), .A2(new_n369), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n448), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n393), .B1(new_n449), .B2(new_n250), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n447), .B1(new_n450), .B2(new_n262), .ZN(new_n451));
  OAI211_X1 g0251(.A(KEYINPUT83), .B(new_n444), .C1(new_n451), .C2(G200), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n443), .A2(new_n452), .A3(new_n420), .A4(new_n426), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT17), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT17), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n435), .A2(new_n455), .A3(new_n452), .A4(new_n443), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n438), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n300), .A2(new_n305), .B1(G20), .B2(G77), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT71), .ZN(new_n461));
  XNOR2_X1  g0261(.A(KEYINPUT15), .B(G87), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n461), .B1(new_n462), .B2(new_n301), .ZN(new_n463));
  INV_X1    g0263(.A(G87), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n464), .A2(KEYINPUT15), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n464), .A2(KEYINPUT15), .ZN(new_n466));
  OAI211_X1 g0266(.A(KEYINPUT71), .B(new_n295), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n460), .A2(new_n463), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G77), .ZN(new_n469));
  INV_X1    g0269(.A(new_n347), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n468), .A2(new_n284), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n347), .A2(new_n351), .A3(G77), .A4(new_n292), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT73), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n472), .A2(new_n473), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G107), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n250), .A2(new_n477), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n368), .A2(new_n369), .A3(new_n209), .ZN(new_n479));
  OAI22_X1  g0279(.A1(new_n248), .A2(new_n249), .B1(new_n210), .B2(new_n254), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n478), .B(new_n262), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n273), .A2(G244), .B1(new_n276), .B2(new_n277), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n481), .A2(new_n281), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(G169), .B1(new_n481), .B2(new_n482), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n476), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g0286(.A(new_n472), .B(new_n473), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n481), .A2(G190), .A3(new_n482), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n481), .A2(new_n482), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G200), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n487), .A2(new_n488), .A3(new_n471), .A4(new_n490), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n326), .A2(new_n389), .A3(new_n459), .A4(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT21), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n347), .A2(new_n351), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n267), .A2(G33), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G116), .ZN(new_n498));
  OAI22_X1  g0298(.A1(new_n496), .A2(new_n498), .B1(G116), .B2(new_n347), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT20), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G283), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT85), .ZN(new_n502));
  XNOR2_X1  g0302(.A(new_n501), .B(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(G20), .B1(new_n294), .B2(G97), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(G116), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G20), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n284), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n500), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g0310(.A(new_n501), .B(KEYINPUT85), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n504), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n512), .A2(KEYINPUT20), .A3(new_n284), .A4(new_n508), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n499), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(G303), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n250), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(G257), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n368), .A2(new_n369), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(G264), .ZN(new_n519));
  OAI22_X1  g0319(.A1(new_n248), .A2(new_n249), .B1(new_n519), .B2(new_n254), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n516), .B(new_n262), .C1(new_n518), .C2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT86), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n522), .A2(new_n268), .A3(KEYINPUT5), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT5), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(KEYINPUT86), .B2(G41), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n269), .A2(G1), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n272), .A2(G1), .A3(G13), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n527), .A2(G270), .A3(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n276), .A2(new_n526), .A3(new_n523), .A4(new_n525), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n521), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G169), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n495), .B1(new_n514), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n510), .A2(new_n513), .ZN(new_n534));
  INV_X1    g0334(.A(new_n499), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n531), .A2(G169), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n536), .A2(new_n537), .A3(KEYINPUT21), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n521), .A2(G179), .A3(new_n529), .A4(new_n530), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n533), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n531), .A2(G200), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n514), .B(new_n543), .C1(new_n440), .C2(new_n531), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n265), .A2(new_n448), .A3(G244), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT4), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n265), .A2(new_n448), .A3(KEYINPUT4), .A4(G244), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n265), .A2(G250), .A3(G1698), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n548), .A2(new_n511), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n262), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n527), .A2(new_n528), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n530), .B1(new_n553), .B2(new_n517), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT87), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT87), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n552), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G200), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT6), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n331), .A2(new_n477), .ZN(new_n562));
  NOR2_X1   g0362(.A1(G97), .A2(G107), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n477), .A2(KEYINPUT84), .A3(KEYINPUT6), .A4(G97), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT84), .ZN(new_n566));
  NAND2_X1  g0366(.A1(KEYINPUT6), .A2(G97), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n566), .B1(new_n567), .B2(G107), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n564), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n569), .A2(G20), .B1(G77), .B2(new_n305), .ZN(new_n570));
  OAI21_X1  g0370(.A(G107), .B1(new_n430), .B2(new_n431), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n351), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n290), .A2(new_n331), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n285), .A2(new_n287), .A3(new_n289), .A4(new_n497), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n573), .B1(new_n574), .B2(new_n331), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n554), .B1(new_n551), .B2(new_n262), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G190), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n560), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  OR2_X1    g0379(.A1(new_n572), .A2(new_n575), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n552), .A2(new_n555), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n310), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n552), .A2(new_n556), .A3(new_n281), .A4(new_n558), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n580), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n517), .A2(new_n254), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(G294), .ZN(new_n588));
  OAI22_X1  g0388(.A1(new_n587), .A2(new_n250), .B1(new_n294), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(G250), .B1(new_n248), .B2(new_n249), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n590), .A2(new_n257), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n262), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n527), .A2(G264), .A3(new_n528), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(new_n530), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n318), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n592), .A2(KEYINPUT89), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT89), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n597), .B(new_n262), .C1(new_n589), .C2(new_n591), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n593), .A2(new_n530), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n596), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n595), .B1(new_n600), .B2(G190), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n225), .B(G87), .C1(new_n248), .C2(new_n249), .ZN(new_n602));
  XNOR2_X1  g0402(.A(new_n602), .B(KEYINPUT22), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT24), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT23), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n225), .B2(G107), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n477), .A2(KEYINPUT23), .A3(G20), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n294), .A2(new_n507), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n606), .A2(new_n607), .B1(new_n608), .B2(new_n225), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n603), .A2(new_n604), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n604), .B1(new_n603), .B2(new_n609), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n284), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n290), .A2(new_n477), .ZN(new_n613));
  XOR2_X1   g0413(.A(new_n613), .B(KEYINPUT25), .Z(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(new_n574), .B2(new_n477), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n601), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n600), .A2(G169), .ZN(new_n618));
  OR2_X1    g0418(.A1(new_n594), .A2(new_n281), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n618), .A2(new_n619), .B1(new_n612), .B2(new_n616), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n528), .A2(G274), .A3(new_n526), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT88), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT88), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n276), .A2(new_n623), .A3(new_n526), .ZN(new_n624));
  INV_X1    g0424(.A(G250), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n526), .A2(new_n625), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n622), .A2(new_n624), .B1(new_n528), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n255), .A2(G238), .A3(new_n256), .ZN(new_n628));
  NAND2_X1  g0428(.A1(G244), .A2(G1698), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n250), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n262), .B1(new_n630), .B2(new_n608), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n310), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n464), .A2(new_n331), .A3(new_n477), .ZN(new_n634));
  OAI211_X1 g0434(.A(KEYINPUT19), .B(new_n634), .C1(new_n332), .C2(G20), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n225), .B(G68), .C1(new_n248), .C2(new_n249), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT19), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(new_n301), .B2(new_n331), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n635), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n639), .A2(new_n284), .B1(new_n470), .B2(new_n462), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n462), .B2(new_n574), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n633), .B(new_n641), .C1(G179), .C2(new_n632), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n640), .B1(new_n464), .B2(new_n574), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n632), .A2(G200), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n627), .A2(new_n631), .A3(G190), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n642), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n617), .A2(new_n620), .A3(new_n647), .ZN(new_n648));
  AND4_X1   g0448(.A1(new_n494), .A2(new_n545), .A3(new_n585), .A4(new_n648), .ZN(G372));
  AND3_X1   g0449(.A1(new_n429), .A2(new_n437), .A3(KEYINPUT92), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT92), .B1(new_n429), .B2(new_n437), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n343), .A2(new_n380), .A3(new_n366), .ZN(new_n654));
  INV_X1    g0454(.A(new_n486), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n382), .A2(new_n388), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n457), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n653), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n321), .A2(new_n325), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n313), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT90), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n574), .A2(new_n464), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n639), .A2(new_n284), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n470), .A2(new_n462), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n662), .B1(new_n663), .B2(new_n666), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n640), .B(KEYINPUT90), .C1(new_n464), .C2(new_n574), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n667), .A2(new_n645), .A3(new_n644), .A4(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n642), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n661), .B1(new_n670), .B2(new_n584), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT91), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT91), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n673), .B(new_n661), .C1(new_n670), .C2(new_n584), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n647), .A2(new_n584), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(KEYINPUT26), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n672), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n642), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n603), .A2(new_n609), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(KEYINPUT24), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n603), .A2(new_n604), .A3(new_n609), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n615), .B1(new_n682), .B2(new_n284), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n601), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n684), .A2(new_n579), .A3(new_n584), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n618), .A2(new_n619), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n612), .A2(new_n616), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n670), .B1(new_n542), .B2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n678), .B1(new_n685), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n677), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n660), .B1(new_n493), .B2(new_n692), .ZN(G369));
  NAND3_X1  g0493(.A1(new_n267), .A2(new_n225), .A3(G13), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n694), .A2(KEYINPUT93), .A3(KEYINPUT27), .ZN(new_n695));
  AOI21_X1  g0495(.A(KEYINPUT93), .B1(new_n694), .B2(KEYINPUT27), .ZN(new_n696));
  OAI221_X1 g0496(.A(G213), .B1(KEYINPUT27), .B2(new_n694), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G343), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n536), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n545), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n542), .B2(new_n700), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G330), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT94), .ZN(new_n704));
  INV_X1    g0504(.A(new_n699), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n704), .B1(new_n683), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n687), .A2(KEYINPUT94), .A3(new_n699), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n706), .A2(new_n688), .A3(new_n684), .A4(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT95), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n620), .A2(new_n699), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n709), .B1(new_n708), .B2(new_n710), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n703), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n688), .A2(new_n699), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n708), .A2(new_n710), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(KEYINPUT95), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n542), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n705), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n716), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n715), .A2(new_n724), .ZN(G399));
  NOR2_X1   g0525(.A1(new_n634), .A2(G116), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n228), .A2(new_n268), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n726), .A2(new_n727), .A3(G1), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(new_n226), .B2(new_n727), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT28), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n675), .A2(new_n661), .ZN(new_n731));
  OAI21_X1  g0531(.A(KEYINPUT26), .B1(new_n670), .B2(new_n584), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n733), .A2(new_n690), .ZN(new_n734));
  OAI21_X1  g0534(.A(KEYINPUT29), .B1(new_n734), .B2(new_n699), .ZN(new_n735));
  AND4_X1   g0535(.A1(new_n631), .A2(new_n627), .A3(new_n592), .A4(new_n593), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n539), .A2(KEYINPUT96), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n539), .A2(KEYINPUT96), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n577), .B(new_n736), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT30), .ZN(new_n740));
  AND4_X1   g0540(.A1(new_n281), .A2(new_n594), .A3(new_n632), .A4(new_n531), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n739), .A2(new_n740), .B1(new_n559), .B2(new_n741), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n736), .A2(new_n577), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n743), .B(KEYINPUT30), .C1(new_n738), .C2(new_n737), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n705), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n745), .A2(KEYINPUT31), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(KEYINPUT31), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n648), .A2(new_n545), .A3(new_n585), .A4(new_n705), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G330), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n699), .B1(new_n677), .B2(new_n690), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT29), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n735), .A2(new_n750), .A3(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n730), .B1(new_n755), .B2(G1), .ZN(G364));
  INV_X1    g0556(.A(G13), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G45), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n727), .A2(G1), .A3(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n265), .A2(new_n228), .ZN(new_n762));
  INV_X1    g0562(.A(G355), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n762), .A2(new_n763), .B1(G116), .B2(new_n228), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n246), .A2(G45), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n250), .A2(new_n228), .ZN(new_n766));
  INV_X1    g0566(.A(new_n226), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n766), .B1(new_n269), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n764), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n224), .B1(G20), .B2(new_n310), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G13), .A2(G33), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n761), .B1(new_n769), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n225), .A2(G190), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n777), .A2(new_n281), .A3(new_n318), .ZN(new_n778));
  INV_X1    g0578(.A(G159), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT32), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT99), .Z(new_n782));
  NAND2_X1  g0582(.A1(G20), .A2(G179), .ZN(new_n783));
  OR3_X1    g0583(.A1(new_n783), .A2(new_n318), .A3(KEYINPUT98), .ZN(new_n784));
  OAI21_X1  g0584(.A(KEYINPUT98), .B1(new_n783), .B2(new_n318), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n784), .A2(G190), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n784), .A2(new_n440), .A3(new_n785), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n782), .B1(new_n201), .B2(new_n786), .C1(new_n203), .C2(new_n787), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n783), .A2(G190), .A3(G200), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n265), .B1(new_n790), .B2(new_n469), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n440), .A2(G179), .A3(G200), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n225), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n791), .B1(G97), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT100), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(new_n318), .B2(G179), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n281), .A2(KEYINPUT100), .A3(G200), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n797), .A2(new_n777), .A3(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G107), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n225), .A2(new_n440), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n797), .A2(new_n802), .A3(new_n798), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G87), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n783), .A2(new_n440), .A3(G200), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT97), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G58), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n795), .A2(new_n801), .A3(new_n805), .A4(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n786), .B(KEYINPUT101), .ZN(new_n810));
  INV_X1    g0610(.A(G326), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n806), .ZN(new_n813));
  INV_X1    g0613(.A(G322), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G311), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n250), .B1(new_n790), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n778), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n815), .B(new_n817), .C1(G329), .C2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n787), .ZN(new_n820));
  XNOR2_X1  g0620(.A(KEYINPUT33), .B(G317), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n794), .A2(G294), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G303), .A2(new_n804), .B1(new_n800), .B2(G283), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n819), .A2(new_n822), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n788), .A2(new_n809), .B1(new_n812), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n776), .B1(new_n826), .B2(new_n770), .ZN(new_n827));
  INV_X1    g0627(.A(new_n773), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n827), .B1(new_n702), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n703), .A2(new_n760), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n702), .A2(G330), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(G396));
  NAND2_X1  g0632(.A1(new_n486), .A2(KEYINPUT102), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT102), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n476), .A2(new_n485), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n476), .A2(new_n699), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n833), .A2(new_n491), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT103), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n836), .A2(new_n491), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n840), .A2(KEYINPUT103), .A3(new_n833), .A4(new_n835), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n839), .A2(new_n841), .B1(new_n655), .B2(new_n699), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n751), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n839), .A2(new_n841), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n844), .B1(new_n751), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n750), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n847), .A2(new_n848), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n849), .A2(new_n760), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n770), .A2(new_n771), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n760), .B1(new_n852), .B2(new_n469), .ZN(new_n853));
  INV_X1    g0653(.A(new_n770), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n818), .A2(G311), .B1(new_n789), .B2(G116), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n265), .B1(G294), .B2(new_n806), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n855), .B(new_n856), .C1(new_n331), .C2(new_n793), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n803), .A2(new_n477), .B1(new_n799), .B2(new_n464), .ZN(new_n858));
  INV_X1    g0658(.A(G283), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n859), .A2(new_n787), .B1(new_n786), .B2(new_n515), .ZN(new_n860));
  NOR3_X1   g0660(.A1(new_n857), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n807), .A2(G143), .B1(G159), .B2(new_n789), .ZN(new_n862));
  INV_X1    g0662(.A(G137), .ZN(new_n863));
  INV_X1    g0663(.A(G150), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n862), .B1(new_n863), .B2(new_n786), .C1(new_n864), .C2(new_n787), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT34), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n799), .A2(new_n203), .ZN(new_n867));
  INV_X1    g0667(.A(G132), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n265), .B1(new_n778), .B2(new_n868), .C1(new_n793), .C2(new_n202), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n867), .B(new_n869), .C1(G50), .C2(new_n804), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n861), .B1(new_n866), .B2(new_n870), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n853), .B1(new_n854), .B2(new_n871), .C1(new_n843), .C2(new_n772), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n851), .A2(new_n872), .ZN(G384));
  NOR2_X1   g0673(.A1(new_n758), .A2(new_n267), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT31), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT107), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n875), .B1(new_n745), .B2(new_n876), .ZN(new_n877));
  AOI211_X1 g0677(.A(KEYINPUT107), .B(new_n705), .C1(new_n742), .C2(new_n744), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n747), .B(new_n748), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n388), .A2(new_n382), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n382), .A2(new_n699), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n880), .A2(new_n654), .A3(new_n881), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n382), .B(new_n699), .C1(new_n381), .C2(new_n388), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n842), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT108), .B1(new_n879), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n416), .A2(new_n288), .ZN(new_n887));
  INV_X1    g0687(.A(new_n417), .ZN(new_n888));
  INV_X1    g0688(.A(new_n415), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n412), .A2(KEYINPUT80), .A3(new_n413), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n888), .B1(new_n891), .B2(new_n409), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n426), .B1(new_n887), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n697), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n458), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n893), .A2(new_n403), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n898), .A2(new_n895), .A3(new_n453), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT37), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n403), .A2(new_n427), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n427), .A2(new_n894), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT37), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n901), .A2(new_n902), .A3(new_n453), .A4(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n897), .A2(KEYINPUT38), .A3(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n901), .A2(new_n902), .A3(new_n453), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n904), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n457), .A2(KEYINPUT105), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT105), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n454), .A2(new_n913), .A3(new_n456), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n912), .B(new_n914), .C1(new_n650), .C2(new_n651), .ZN(new_n915));
  INV_X1    g0715(.A(new_n902), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n911), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n907), .B1(new_n917), .B2(KEYINPUT38), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n879), .A2(new_n884), .A3(KEYINPUT108), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n886), .A2(new_n918), .A3(KEYINPUT40), .A4(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT40), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT38), .B1(new_n897), .B2(new_n905), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n906), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n879), .A2(new_n884), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n920), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n494), .A2(new_n879), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n928), .A2(G330), .A3(new_n929), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(KEYINPUT109), .Z(new_n931));
  NOR2_X1   g0731(.A1(new_n880), .A2(new_n699), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n458), .A2(new_n896), .B1(new_n900), .B2(new_n904), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT39), .B1(new_n933), .B2(KEYINPUT38), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n917), .B2(KEYINPUT38), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT39), .B1(new_n906), .B2(new_n922), .ZN(new_n936));
  AND3_X1   g0736(.A1(new_n935), .A2(KEYINPUT106), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT106), .B1(new_n935), .B2(new_n936), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n932), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n833), .A2(new_n835), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n940), .A2(new_n699), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n751), .B2(new_n846), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n882), .A2(new_n883), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n942), .A2(new_n923), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n652), .B2(new_n697), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n939), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n493), .B1(new_n735), .B2(new_n753), .ZN(new_n948));
  INV_X1    g0748(.A(new_n660), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n947), .B(new_n950), .Z(new_n951));
  AOI21_X1  g0751(.A(new_n874), .B1(new_n931), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n931), .B2(new_n951), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n569), .A2(KEYINPUT35), .ZN(new_n954));
  NOR3_X1   g0754(.A1(new_n224), .A2(new_n225), .A3(new_n507), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n569), .B2(KEYINPUT35), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT104), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(new_n957), .B2(new_n956), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT36), .Z(new_n960));
  NOR3_X1   g0760(.A1(new_n404), .A2(new_n226), .A3(new_n469), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n203), .A2(G50), .ZN(new_n962));
  OAI211_X1 g0762(.A(G1), .B(new_n757), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n953), .A2(new_n960), .A3(new_n963), .ZN(G367));
  AOI21_X1  g0764(.A(new_n722), .B1(new_n718), .B2(new_n719), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n585), .B1(new_n576), .B2(new_n705), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n584), .A2(new_n705), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n969), .A2(KEYINPUT42), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n966), .A2(new_n688), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n699), .B1(new_n971), .B2(new_n584), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(new_n969), .B2(KEYINPUT42), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n667), .A2(new_n668), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n699), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n975), .A2(new_n642), .A3(new_n669), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n976), .A2(KEYINPUT110), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(KEYINPUT110), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n977), .B(new_n978), .C1(new_n642), .C2(new_n975), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n970), .A2(new_n973), .B1(KEYINPUT43), .B2(new_n979), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n979), .A2(KEYINPUT43), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n980), .B(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n714), .A2(new_n968), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n982), .B(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n759), .A2(G1), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n727), .B(KEYINPUT41), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n723), .B1(new_n711), .B2(new_n712), .ZN(new_n989));
  INV_X1    g0789(.A(new_n716), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n989), .A2(new_n990), .A3(new_n968), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT45), .ZN(new_n992));
  OAI21_X1  g0792(.A(KEYINPUT44), .B1(new_n724), .B2(new_n968), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT44), .ZN(new_n994));
  INV_X1    g0794(.A(new_n968), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(new_n965), .C2(new_n716), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n714), .B1(new_n992), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT111), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n713), .A2(new_n722), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n1000), .A2(G330), .A3(new_n702), .A4(new_n989), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n720), .A2(new_n723), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n703), .B1(new_n1002), .B2(new_n965), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n755), .A2(new_n999), .A3(new_n1001), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1001), .ZN(new_n1005));
  OAI21_X1  g0805(.A(KEYINPUT111), .B1(new_n1005), .B2(new_n754), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n724), .A2(KEYINPUT45), .A3(new_n968), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT45), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n991), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1010), .A2(new_n715), .A3(new_n993), .A4(new_n996), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n998), .A2(new_n1004), .A3(new_n1006), .A4(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n988), .B1(new_n1012), .B2(new_n755), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n987), .B1(new_n1013), .B2(KEYINPUT112), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT112), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1015), .B(new_n988), .C1(new_n1012), .C2(new_n755), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n985), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n774), .B1(new_n228), .B2(new_n462), .ZN(new_n1018));
  AND3_X1   g0818(.A1(new_n238), .A2(new_n228), .A3(new_n250), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n761), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n803), .A2(new_n202), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G50), .A2(new_n789), .B1(new_n806), .B2(G150), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n203), .B2(new_n793), .C1(new_n863), .C2(new_n778), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1021), .B(new_n1023), .C1(G159), .C2(new_n820), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n265), .B1(new_n799), .B2(new_n469), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT115), .Z(new_n1026));
  INV_X1    g0826(.A(G143), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1024), .B(new_n1026), .C1(new_n1027), .C2(new_n810), .ZN(new_n1028));
  AOI21_X1  g0828(.A(KEYINPUT46), .B1(new_n804), .B2(G116), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT114), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n820), .A2(G294), .ZN(new_n1031));
  INV_X1    g0831(.A(G317), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n250), .B1(new_n778), .B2(new_n1032), .C1(new_n790), .C2(new_n859), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G107), .B2(new_n794), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n807), .A2(G303), .B1(G97), .B2(new_n800), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1030), .A2(new_n1031), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n804), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT113), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n816), .B2(new_n810), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1028), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT47), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1020), .B1(new_n1041), .B2(new_n770), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n828), .B2(new_n979), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1017), .A2(new_n1043), .ZN(G387));
  NAND2_X1  g0844(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n727), .B1(new_n1005), .B2(new_n754), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n720), .A2(new_n828), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n762), .A2(new_n726), .B1(G107), .B2(new_n228), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n235), .A2(G45), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n726), .ZN(new_n1051));
  AOI211_X1 g0851(.A(G45), .B(new_n1051), .C1(G68), .C2(G77), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n300), .A2(new_n201), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT50), .Z(new_n1054));
  AOI21_X1  g0854(.A(new_n766), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1049), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n250), .B1(G68), .B2(new_n789), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n201), .B2(new_n813), .C1(new_n864), .C2(new_n778), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n804), .A2(G77), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n331), .B2(new_n799), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n779), .A2(new_n786), .B1(new_n787), .B2(new_n423), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n793), .A2(new_n462), .ZN(new_n1062));
  NOR4_X1   g0862(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n250), .B1(new_n778), .B2(new_n811), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n807), .A2(G317), .B1(G303), .B2(new_n789), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n816), .B2(new_n787), .C1(new_n810), .C2(new_n814), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT48), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G283), .A2(new_n794), .B1(new_n804), .B2(G294), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT49), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1064), .B(new_n1073), .C1(G116), .C2(new_n800), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1063), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n761), .B1(new_n775), .B2(new_n1056), .C1(new_n1076), .C2(new_n854), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1047), .B1(new_n1005), .B2(new_n987), .C1(new_n1048), .C2(new_n1077), .ZN(G393));
  OAI21_X1  g0878(.A(new_n774), .B1(new_n331), .B2(new_n228), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n242), .A2(new_n766), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n761), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n820), .A2(G303), .B1(G116), .B2(new_n794), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1082), .A2(KEYINPUT116), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(KEYINPUT116), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n804), .A2(G283), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n250), .B1(new_n778), .B2(new_n814), .C1(new_n790), .C2(new_n588), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(G107), .B2(new_n800), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .A4(new_n1087), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n786), .A2(new_n1032), .B1(new_n816), .B2(new_n813), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT52), .Z(new_n1090));
  OAI22_X1  g0890(.A1(new_n786), .A2(new_n864), .B1(new_n779), .B2(new_n813), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT51), .Z(new_n1092));
  OAI21_X1  g0892(.A(new_n265), .B1(new_n778), .B2(new_n1027), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n793), .A2(new_n469), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1093), .B(new_n1094), .C1(new_n300), .C2(new_n789), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(G68), .A2(new_n804), .B1(new_n800), .B2(G87), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1095), .B(new_n1096), .C1(new_n201), .C2(new_n787), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n1088), .A2(new_n1090), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1081), .B1(new_n1098), .B2(new_n770), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT117), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n968), .B2(new_n828), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n998), .A2(new_n1011), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1101), .B1(new_n1102), .B2(new_n987), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1045), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT118), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1102), .A2(KEYINPUT118), .A3(new_n1045), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n727), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n1012), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1103), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(G390));
  NAND3_X1  g0912(.A1(new_n749), .A2(G330), .A3(new_n843), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n1113), .A2(new_n944), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n879), .A2(G330), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n944), .B1(new_n1115), .B2(new_n842), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n699), .B1(new_n733), .B2(new_n690), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n941), .B1(new_n1117), .B2(new_n846), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1114), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1115), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1120), .A2(new_n884), .B1(new_n944), .B2(new_n1113), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1119), .B1(new_n942), .B2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n493), .A2(new_n1115), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n948), .A2(new_n949), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n935), .A2(new_n936), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT106), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n935), .A2(new_n936), .A3(KEYINPUT106), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n932), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n942), .B2(new_n944), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1128), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n1118), .A2(new_n944), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1133), .A2(new_n918), .A3(new_n1130), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n1132), .A2(new_n1134), .A3(new_n1114), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1120), .A2(new_n884), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1125), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1136), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n691), .A2(new_n705), .A3(new_n846), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n941), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n932), .B1(new_n1142), .B2(new_n943), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n937), .A2(new_n938), .A3(new_n1143), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1133), .A2(new_n918), .A3(new_n1130), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1139), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1132), .A2(new_n1134), .A3(new_n1114), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1123), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n735), .A2(new_n753), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1148), .B(new_n660), .C1(new_n1149), .C2(new_n493), .ZN(new_n1150));
  OR2_X1    g0950(.A1(new_n1121), .A2(new_n942), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1150), .B1(new_n1151), .B2(new_n1119), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1146), .A2(new_n1147), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1138), .A2(new_n1109), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n852), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n805), .A2(new_n250), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT120), .Z(new_n1157));
  AOI22_X1  g0957(.A1(new_n818), .A2(G294), .B1(new_n806), .B2(G116), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n331), .B2(new_n790), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n477), .A2(new_n787), .B1(new_n786), .B2(new_n859), .ZN(new_n1160));
  NOR4_X1   g0960(.A1(new_n1159), .A2(new_n1160), .A3(new_n867), .A4(new_n1094), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(KEYINPUT54), .B(G143), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT119), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n1163), .A2(new_n790), .B1(new_n201), .B2(new_n799), .ZN(new_n1164));
  INV_X1    g0964(.A(G128), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n1165), .A2(new_n786), .B1(new_n787), .B2(new_n863), .ZN(new_n1166));
  INV_X1    g0966(.A(G125), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n265), .B1(new_n778), .B2(new_n1167), .C1(new_n813), .C2(new_n868), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n793), .A2(new_n779), .ZN(new_n1169));
  NOR4_X1   g0969(.A1(new_n1164), .A2(new_n1166), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n803), .A2(new_n864), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT53), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1157), .A2(new_n1161), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n761), .B1(new_n300), .B2(new_n1155), .C1(new_n1173), .C2(new_n854), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n937), .A2(new_n938), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1174), .B1(new_n1175), .B2(new_n771), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1176), .B1(new_n1177), .B2(new_n986), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1154), .A2(new_n1178), .ZN(G378));
  NAND2_X1  g0979(.A1(new_n1153), .A2(new_n1124), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n912), .A2(new_n914), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n916), .B1(new_n1181), .B2(new_n652), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT38), .B1(new_n1182), .B2(new_n910), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n919), .B(KEYINPUT40), .C1(new_n1183), .C2(new_n906), .ZN(new_n1184));
  OAI211_X1 g0984(.A(G330), .B(new_n925), .C1(new_n1184), .C2(new_n885), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n309), .A2(new_n894), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n326), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n326), .A2(new_n1188), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1186), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1191), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1186), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1193), .A2(new_n1194), .A3(new_n1189), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1192), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1185), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1192), .A2(new_n1195), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1198), .A2(new_n920), .A3(G330), .A4(new_n925), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n947), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1197), .A2(new_n1199), .A3(new_n939), .A4(new_n946), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1180), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT57), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1153), .A2(new_n1124), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(KEYINPUT57), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1206), .A2(new_n1109), .A3(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT123), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n265), .A2(G41), .ZN(new_n1211));
  AOI211_X1 g1011(.A(G50), .B(new_n1211), .C1(new_n294), .C2(new_n268), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n800), .A2(G58), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n818), .A2(G283), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1059), .A2(new_n1213), .A3(new_n1211), .A4(new_n1214), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT121), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n806), .A2(G107), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n790), .B2(new_n462), .C1(new_n203), .C2(new_n793), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G97), .B2(new_n820), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1216), .B(new_n1219), .C1(new_n507), .C2(new_n786), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT58), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1212), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G128), .A2(new_n806), .B1(new_n789), .B2(G137), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n1163), .B2(new_n803), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n786), .A2(new_n1167), .B1(new_n864), .B2(new_n793), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT122), .Z(new_n1226));
  AOI211_X1 g1026(.A(new_n1224), .B(new_n1226), .C1(G132), .C2(new_n820), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n800), .A2(G159), .ZN(new_n1230));
  AOI211_X1 g1030(.A(G33), .B(G41), .C1(new_n818), .C2(G124), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1222), .B1(new_n1221), .B2(new_n1220), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n770), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n760), .B1(new_n852), .B2(new_n201), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1235), .B(new_n1236), .C1(new_n1198), .C2(new_n772), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n1203), .B2(new_n986), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1209), .A2(new_n1210), .A3(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1210), .B1(new_n1209), .B2(new_n1239), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(G375));
  NAND2_X1  g1043(.A1(new_n944), .A2(new_n771), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n761), .B1(new_n1155), .B2(G68), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n265), .B1(new_n778), .B2(new_n1165), .C1(new_n790), .C2(new_n864), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(G50), .B2(new_n794), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n1247), .B1(new_n868), .B2(new_n786), .C1(new_n787), .C2(new_n1163), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n807), .A2(G137), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1249), .B(new_n1213), .C1(new_n779), .C2(new_n803), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n790), .A2(new_n477), .B1(new_n778), .B2(new_n515), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n265), .B(new_n1251), .C1(G283), .C2(new_n806), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(G97), .A2(new_n804), .B1(new_n800), .B2(G77), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1252), .B(new_n1253), .C1(new_n462), .C2(new_n793), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n507), .A2(new_n787), .B1(new_n786), .B2(new_n588), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n1248), .A2(new_n1250), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1245), .B1(new_n1256), .B2(new_n770), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1122), .A2(new_n986), .B1(new_n1244), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n988), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1125), .A2(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1258), .B1(new_n1260), .B2(new_n1261), .ZN(G381));
  OAI21_X1  g1062(.A(new_n1109), .B1(new_n1207), .B2(KEYINPUT57), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1180), .A2(KEYINPUT57), .A3(new_n1203), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1239), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(KEYINPUT123), .ZN(new_n1266));
  AOI21_X1  g1066(.A(G378), .B1(new_n1266), .B2(new_n1240), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1017), .A2(new_n1043), .A3(new_n1111), .ZN(new_n1268));
  NOR4_X1   g1068(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1267), .A2(new_n1271), .ZN(G407));
  OAI21_X1  g1072(.A(new_n1267), .B1(new_n1271), .B2(new_n698), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(G213), .ZN(G409));
  XOR2_X1   g1074(.A(G393), .B(G396), .Z(new_n1275));
  AOI21_X1  g1075(.A(new_n1111), .B1(new_n1017), .B2(new_n1043), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1275), .B1(new_n1268), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(G387), .A2(G390), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1017), .A2(new_n1043), .A3(new_n1111), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1275), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1278), .A2(new_n1279), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1277), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(G213), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1283), .A2(G343), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1154), .A2(new_n1178), .A3(new_n1237), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1180), .A2(new_n1259), .A3(new_n1203), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1203), .A2(KEYINPUT124), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT124), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1289), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1290));
  OR3_X1    g1090(.A1(new_n1288), .A2(new_n987), .A3(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1284), .B1(new_n1287), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1265), .A2(G378), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT60), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1294), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1151), .A2(new_n1150), .A3(KEYINPUT60), .A4(new_n1119), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1295), .A2(new_n1296), .A3(new_n1109), .A4(new_n1125), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1297), .A2(G384), .A3(new_n1258), .ZN(new_n1298));
  AOI21_X1  g1098(.A(G384), .B1(new_n1297), .B2(new_n1258), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1292), .A2(new_n1293), .A3(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(KEYINPUT125), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT62), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT125), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1292), .A2(new_n1293), .A3(new_n1304), .A4(new_n1300), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1302), .A2(new_n1303), .A3(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1284), .A2(G2897), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1300), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(new_n1283), .A2(KEYINPUT126), .A3(G343), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1307), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1300), .A2(KEYINPUT126), .A3(G2897), .A4(new_n1284), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(G378), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1313), .B1(new_n1209), .B2(new_n1239), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1180), .A2(new_n1259), .A3(new_n1203), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1315), .A2(new_n1154), .A3(new_n1178), .A4(new_n1237), .ZN(new_n1316));
  NOR3_X1   g1116(.A1(new_n1288), .A2(new_n987), .A3(new_n1290), .ZN(new_n1317));
  OAI22_X1  g1117(.A1(new_n1316), .A2(new_n1317), .B1(new_n1283), .B2(G343), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1312), .B1(new_n1314), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT61), .ZN(new_n1320));
  NOR3_X1   g1120(.A1(new_n1314), .A2(new_n1318), .A3(new_n1308), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n1319), .B(new_n1320), .C1(new_n1321), .C2(new_n1303), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1282), .B1(new_n1306), .B2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT63), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1314), .A2(new_n1318), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1304), .B1(new_n1325), .B2(new_n1300), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1305), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1324), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1277), .A2(new_n1281), .A3(new_n1320), .ZN(new_n1329));
  AOI22_X1  g1129(.A1(new_n1292), .A2(new_n1293), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1329), .B1(KEYINPUT127), .B2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT127), .ZN(new_n1332));
  AOI22_X1  g1132(.A1(new_n1319), .A2(new_n1332), .B1(new_n1321), .B2(KEYINPUT63), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1328), .A2(new_n1331), .A3(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1323), .A2(new_n1334), .ZN(G405));
  INV_X1    g1135(.A(new_n1267), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1336), .A2(new_n1282), .A3(new_n1293), .ZN(new_n1337));
  OAI211_X1 g1137(.A(new_n1277), .B(new_n1281), .C1(new_n1267), .C2(new_n1314), .ZN(new_n1338));
  AND3_X1   g1138(.A1(new_n1337), .A2(new_n1300), .A3(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1300), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1339), .A2(new_n1340), .ZN(G402));
endmodule


