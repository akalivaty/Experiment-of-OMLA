//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XOR2_X1   g002(.A(KEYINPUT2), .B(G113), .Z(new_n189));
  XNOR2_X1  g003(.A(G116), .B(G119), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT82), .A3(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT3), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n192), .A2(G104), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n197), .A2(new_n192), .A3(KEYINPUT82), .A4(G104), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(new_n196), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT83), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n194), .A2(new_n196), .A3(KEYINPUT83), .A4(new_n198), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(G101), .A3(new_n202), .ZN(new_n203));
  OR2_X1    g017(.A1(new_n199), .A2(G101), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(KEYINPUT4), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT4), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n201), .A2(new_n206), .A3(G101), .A4(new_n202), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT84), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n207), .A2(new_n208), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n191), .B(new_n205), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G104), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(G107), .ZN(new_n213));
  OAI21_X1  g027(.A(G101), .B1(new_n213), .B2(new_n195), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n204), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G113), .ZN(new_n217));
  INV_X1    g031(.A(G119), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n218), .A2(G116), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT5), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n217), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n190), .A2(KEYINPUT5), .ZN(new_n222));
  AOI22_X1  g036(.A1(new_n221), .A2(new_n222), .B1(new_n190), .B2(new_n189), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n216), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n211), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g039(.A(G110), .B(G122), .Z(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n226), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n211), .A2(new_n228), .A3(new_n224), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n227), .A2(KEYINPUT6), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G143), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(G146), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  XOR2_X1   g047(.A(KEYINPUT64), .B(G146), .Z(new_n234));
  OAI21_X1  g048(.A(new_n233), .B1(new_n234), .B2(G143), .ZN(new_n235));
  NAND2_X1  g049(.A1(KEYINPUT0), .A2(G128), .ZN(new_n236));
  NOR2_X1   g050(.A1(KEYINPUT0), .A2(G128), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n235), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n234), .A2(G143), .ZN(new_n240));
  INV_X1    g054(.A(G146), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n241), .A2(G143), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n236), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n240), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n239), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G125), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT64), .B(G146), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(new_n231), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT1), .ZN(new_n250));
  OAI21_X1  g064(.A(G128), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n235), .ZN(new_n252));
  INV_X1    g066(.A(G125), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n240), .A2(new_n250), .A3(G128), .A4(new_n243), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n247), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G953), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G224), .ZN(new_n258));
  XOR2_X1   g072(.A(new_n256), .B(new_n258), .Z(new_n259));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n225), .A2(new_n260), .A3(new_n226), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n230), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G902), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n215), .A2(new_n223), .ZN(new_n264));
  XOR2_X1   g078(.A(new_n226), .B(KEYINPUT8), .Z(new_n265));
  XOR2_X1   g079(.A(new_n222), .B(KEYINPUT87), .Z(new_n266));
  AOI22_X1  g080(.A1(new_n266), .A2(new_n221), .B1(new_n190), .B2(new_n189), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n264), .B(new_n265), .C1(new_n267), .C2(new_n215), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n256), .A2(G224), .A3(new_n257), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n247), .A2(new_n255), .A3(KEYINPUT7), .A4(new_n258), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n256), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n271), .B(new_n229), .C1(KEYINPUT7), .C2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n262), .A2(new_n263), .A3(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(G210), .B1(G237), .B2(G902), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n262), .A2(new_n263), .A3(new_n275), .A4(new_n273), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n188), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(G234), .A2(G237), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(G952), .A3(new_n257), .ZN(new_n281));
  XOR2_X1   g095(.A(KEYINPUT21), .B(G898), .Z(new_n282));
  NAND3_X1  g096(.A1(new_n280), .A2(G902), .A3(G953), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n279), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G469), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT66), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n288), .A2(G137), .ZN(new_n289));
  INV_X1    g103(.A(G137), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(KEYINPUT66), .ZN(new_n291));
  OAI211_X1 g105(.A(KEYINPUT11), .B(G134), .C1(new_n289), .C2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT67), .B1(new_n290), .B2(G134), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT67), .ZN(new_n294));
  INV_X1    g108(.A(G134), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(new_n295), .A3(G137), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n290), .A2(G134), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT11), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n293), .A2(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n292), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT68), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(new_n301), .A3(G131), .ZN(new_n302));
  INV_X1    g116(.A(G131), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n292), .B(new_n299), .C1(KEYINPUT68), .C2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n215), .A2(new_n252), .A3(new_n254), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(G128), .B1(new_n232), .B2(new_n250), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n308), .B1(new_n249), .B2(new_n242), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n215), .B1(new_n254), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n305), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT12), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT85), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n305), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n254), .A2(new_n309), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n216), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n314), .B1(new_n316), .B2(new_n306), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT85), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT12), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n311), .A2(KEYINPUT86), .A3(new_n312), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT86), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n321), .B1(new_n317), .B2(KEYINPUT12), .ZN(new_n322));
  AOI22_X1  g136(.A1(new_n313), .A2(new_n319), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT72), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n246), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n239), .A2(KEYINPUT72), .A3(new_n245), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n327), .B(new_n205), .C1(new_n209), .C2(new_n210), .ZN(new_n328));
  OR2_X1    g142(.A1(new_n310), .A2(KEYINPUT10), .ZN(new_n329));
  INV_X1    g143(.A(G128), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n330), .B1(new_n240), .B2(KEYINPUT1), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n232), .B1(new_n248), .B2(new_n231), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n254), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n216), .A2(new_n333), .A3(KEYINPUT10), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n328), .A2(new_n329), .A3(new_n314), .A4(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(G110), .B(G140), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n257), .A2(G227), .ZN(new_n337));
  XOR2_X1   g151(.A(new_n336), .B(new_n337), .Z(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n323), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n328), .A2(new_n329), .A3(new_n334), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n305), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n338), .B1(new_n342), .B2(new_n335), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n287), .B(new_n263), .C1(new_n340), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(G469), .A2(G902), .ZN(new_n345));
  INV_X1    g159(.A(new_n338), .ZN(new_n346));
  INV_X1    g160(.A(new_n335), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n346), .B1(new_n323), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n342), .A2(new_n335), .A3(new_n338), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(G469), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n344), .A2(new_n345), .A3(new_n350), .ZN(new_n351));
  XOR2_X1   g165(.A(KEYINPUT9), .B(G234), .Z(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(KEYINPUT81), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n263), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n354), .A2(G221), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(G475), .A2(G902), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G237), .ZN(new_n361));
  AND4_X1   g175(.A1(G143), .A2(new_n361), .A3(new_n257), .A4(G214), .ZN(new_n362));
  NOR2_X1   g176(.A1(G237), .A2(G953), .ZN(new_n363));
  AOI21_X1  g177(.A(G143), .B1(new_n363), .B2(G214), .ZN(new_n364));
  OAI21_X1  g178(.A(G131), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT17), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n361), .A2(new_n257), .A3(G214), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n231), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n363), .A2(G143), .A3(G214), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n303), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n365), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G140), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G125), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n253), .A2(G140), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT16), .ZN(new_n375));
  OR3_X1    g189(.A1(new_n253), .A2(KEYINPUT16), .A3(G140), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(G146), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n376), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n241), .ZN(new_n379));
  OAI211_X1 g193(.A(KEYINPUT17), .B(G131), .C1(new_n362), .C2(new_n364), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n371), .A2(new_n377), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(G113), .B(G122), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(new_n212), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n362), .A2(new_n364), .ZN(new_n384));
  NAND2_X1  g198(.A1(KEYINPUT18), .A2(G131), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI211_X1 g200(.A(KEYINPUT18), .B(G131), .C1(new_n362), .C2(new_n364), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n373), .A2(new_n374), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(KEYINPUT78), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT78), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n373), .A2(new_n374), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n248), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n388), .A2(G146), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n386), .B(new_n387), .C1(new_n392), .C2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n381), .A2(new_n383), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT89), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT89), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n381), .A2(new_n395), .A3(new_n398), .A4(new_n383), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT19), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n373), .A2(new_n374), .A3(new_n390), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n390), .B1(new_n373), .B2(new_n374), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n388), .A2(KEYINPUT19), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n234), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT77), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n377), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n375), .A2(new_n376), .A3(KEYINPUT77), .A4(G146), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n365), .A2(new_n370), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n406), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n395), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT88), .ZN(new_n414));
  INV_X1    g228(.A(new_n383), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n408), .A2(new_n409), .B1(new_n365), .B2(new_n370), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n234), .B1(new_n402), .B2(new_n403), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n418), .A2(new_n393), .B1(new_n384), .B2(new_n385), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n406), .A2(new_n417), .B1(new_n419), .B2(new_n387), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT88), .B1(new_n420), .B2(new_n383), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n400), .A2(new_n416), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT90), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n414), .B1(new_n413), .B2(new_n415), .ZN(new_n424));
  AOI211_X1 g238(.A(KEYINPUT88), .B(new_n383), .C1(new_n412), .C2(new_n395), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT90), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n427), .A3(new_n400), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n360), .B1(new_n423), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT20), .ZN(new_n430));
  OAI21_X1  g244(.A(KEYINPUT91), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n427), .B1(new_n426), .B2(new_n400), .ZN(new_n432));
  AND4_X1   g246(.A1(new_n427), .A2(new_n400), .A3(new_n416), .A4(new_n421), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n359), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT91), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n435), .A3(KEYINPUT20), .ZN(new_n436));
  XOR2_X1   g250(.A(new_n359), .B(KEYINPUT92), .Z(new_n437));
  NAND3_X1  g251(.A1(new_n422), .A2(new_n430), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT93), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n438), .B(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n431), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n383), .B1(new_n381), .B2(new_n395), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n442), .B1(new_n397), .B2(new_n399), .ZN(new_n443));
  OAI21_X1  g257(.A(G475), .B1(new_n443), .B2(G902), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G122), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n446), .A2(G116), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(G116), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n192), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n330), .A2(G143), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n231), .A2(G128), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(new_n295), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT14), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n449), .B1(new_n447), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT94), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n457), .B(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n459), .B1(new_n456), .B2(new_n447), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n451), .B(new_n455), .C1(new_n460), .C2(new_n192), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n450), .B(new_n192), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n454), .A2(new_n295), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n453), .B1(KEYINPUT13), .B2(new_n452), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(KEYINPUT13), .B2(new_n452), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(G134), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n462), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n353), .A2(G217), .A3(new_n257), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(KEYINPUT95), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n468), .A2(new_n470), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(G902), .ZN(new_n475));
  INV_X1    g289(.A(G478), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(KEYINPUT15), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n475), .B(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n445), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n286), .A2(new_n358), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(G217), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n483), .B1(G234), .B2(new_n263), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT25), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n257), .A2(G221), .A3(G234), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(KEYINPUT80), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT22), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n488), .B(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(G137), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n218), .A2(G128), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n330), .A2(G119), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT24), .B(G110), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT76), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT76), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n494), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT23), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n330), .A2(KEYINPUT23), .A3(G119), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n492), .A3(new_n502), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n497), .B(new_n499), .C1(G110), .C2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(new_n410), .A3(new_n418), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT79), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n505), .B(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT74), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT74), .A4(new_n492), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(G110), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n379), .A2(new_n377), .ZN(new_n512));
  OR2_X1    g326(.A1(new_n494), .A2(new_n495), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT75), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT75), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n511), .A2(new_n512), .A3(new_n516), .A4(new_n513), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n491), .B1(new_n507), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n505), .B(KEYINPUT79), .ZN(new_n520));
  INV_X1    g334(.A(new_n518), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n490), .B(new_n290), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n486), .B1(new_n524), .B2(G902), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n519), .A2(new_n523), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(KEYINPUT25), .A3(new_n263), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n485), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n484), .A2(G902), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n528), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT65), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n332), .A2(new_n244), .A3(new_n237), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n249), .A2(new_n242), .A3(new_n236), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n239), .A2(KEYINPUT65), .A3(new_n245), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n535), .A2(new_n305), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n292), .A2(new_n299), .A3(new_n303), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n290), .A2(KEYINPUT66), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n288), .A2(G137), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n541), .A3(new_n295), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n297), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(G131), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT69), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT69), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n539), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT70), .B1(new_n549), .B2(new_n333), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n539), .A2(new_n547), .A3(new_n544), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n547), .B1(new_n539), .B2(new_n544), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n333), .B(KEYINPUT70), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n538), .B1(new_n550), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT71), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT30), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n333), .B1(new_n551), .B2(new_n552), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT70), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n537), .B1(new_n561), .B2(new_n553), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT71), .B1(new_n562), .B2(KEYINPUT30), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n327), .A2(new_n305), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n333), .A2(new_n544), .A3(new_n539), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(KEYINPUT30), .A3(new_n565), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n558), .A2(new_n563), .A3(new_n191), .A4(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n191), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n564), .A2(new_n568), .A3(new_n565), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n363), .A2(G210), .ZN(new_n570));
  XOR2_X1   g384(.A(new_n570), .B(KEYINPUT27), .Z(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(KEYINPUT26), .ZN(new_n572));
  INV_X1    g386(.A(G101), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n572), .B(new_n573), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n567), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT31), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT28), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n569), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n564), .A2(KEYINPUT28), .A3(new_n568), .A4(new_n565), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n579), .B(new_n580), .C1(new_n568), .C2(new_n562), .ZN(new_n581));
  INV_X1    g395(.A(new_n574), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT31), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n567), .A2(new_n585), .A3(new_n575), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n577), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(G472), .A2(G902), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT32), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G472), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n567), .A2(new_n569), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n582), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT29), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n581), .A2(new_n582), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n314), .B1(new_n326), .B2(new_n325), .ZN(new_n597));
  INV_X1    g411(.A(new_n565), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n191), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n599), .A2(new_n569), .A3(KEYINPUT73), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT73), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n564), .A2(new_n601), .A3(new_n568), .A4(new_n565), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n600), .A2(KEYINPUT28), .A3(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n603), .A2(KEYINPUT29), .A3(new_n574), .A4(new_n579), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n263), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n590), .B1(new_n596), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n589), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n587), .A2(KEYINPUT32), .A3(new_n588), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n531), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n482), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  AND3_X1   g426(.A1(new_n567), .A2(new_n585), .A3(new_n575), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n585), .B1(new_n567), .B2(new_n575), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n613), .A2(new_n614), .A3(new_n583), .ZN(new_n615));
  OAI21_X1  g429(.A(KEYINPUT96), .B1(new_n615), .B2(G902), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT96), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n587), .A2(new_n617), .A3(new_n263), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n616), .A2(G472), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT97), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n587), .A2(new_n588), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n357), .A2(new_n531), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n616), .A2(KEYINPUT97), .A3(G472), .A4(new_n618), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n621), .A2(new_n622), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n626), .B1(new_n472), .B2(new_n473), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n461), .A2(new_n467), .ZN(new_n628));
  INV_X1    g442(.A(new_n470), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(KEYINPUT33), .A3(new_n471), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n627), .A2(G478), .A3(new_n263), .A4(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n476), .B1(new_n474), .B2(G902), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n441), .B2(new_n444), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n637), .A2(new_n285), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n625), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(new_n212), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT98), .B(KEYINPUT34), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  OAI211_X1 g457(.A(new_n431), .B(new_n436), .C1(KEYINPUT20), .C2(new_n434), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n644), .A2(new_n444), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n286), .A2(new_n479), .A3(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n625), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT99), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT35), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G107), .ZN(G9));
  INV_X1    g464(.A(KEYINPUT101), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n507), .A2(new_n518), .A3(KEYINPUT100), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n522), .A2(KEYINPUT36), .ZN(new_n654));
  OAI21_X1  g468(.A(KEYINPUT100), .B1(new_n507), .B2(new_n518), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n520), .B2(new_n521), .ZN(new_n658));
  OAI22_X1  g472(.A1(new_n652), .A2(new_n658), .B1(KEYINPUT36), .B2(new_n522), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n656), .A2(new_n659), .A3(new_n529), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n651), .B1(new_n528), .B2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n527), .ZN(new_n663));
  AOI21_X1  g477(.A(KEYINPUT25), .B1(new_n526), .B2(new_n263), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n484), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n665), .A2(KEYINPUT101), .A3(new_n660), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n621), .A2(new_n622), .A3(new_n624), .A4(new_n667), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n668), .A2(KEYINPUT102), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(KEYINPUT102), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n669), .A2(new_n670), .A3(new_n481), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT37), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G110), .ZN(G12));
  INV_X1    g487(.A(KEYINPUT32), .ZN(new_n674));
  INV_X1    g488(.A(new_n588), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n674), .B1(new_n615), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n574), .B1(new_n567), .B2(new_n569), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n677), .A2(new_n594), .A3(KEYINPUT29), .ZN(new_n678));
  OAI21_X1  g492(.A(G472), .B1(new_n678), .B2(new_n605), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n676), .A2(new_n609), .A3(new_n679), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n667), .A2(new_n279), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n680), .A2(new_n681), .A3(new_n358), .ZN(new_n682));
  INV_X1    g496(.A(new_n281), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT103), .B(G900), .Z(new_n684));
  INV_X1    g498(.A(new_n283), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n645), .A2(new_n479), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n682), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT104), .B(G128), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G30));
  INV_X1    g506(.A(new_n445), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n693), .A2(new_n188), .A3(new_n478), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n665), .A3(new_n660), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT105), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n574), .B1(new_n600), .B2(new_n602), .ZN(new_n697));
  AOI211_X1 g511(.A(G902), .B(new_n697), .C1(new_n591), .C2(new_n574), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n676), .B(new_n609), .C1(new_n590), .C2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n277), .A2(new_n278), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT38), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n696), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n703));
  OR2_X1    g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n686), .B(KEYINPUT39), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n357), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT40), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n704), .A2(new_n705), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G143), .ZN(G45));
  AND2_X1   g524(.A1(new_n680), .A2(new_n681), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n712));
  AND4_X1   g526(.A1(KEYINPUT107), .A2(new_n445), .A3(new_n634), .A4(new_n687), .ZN(new_n713));
  AOI21_X1  g527(.A(KEYINPUT107), .B1(new_n636), .B2(new_n687), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n711), .A2(new_n712), .A3(new_n358), .A4(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n445), .A2(new_n634), .A3(new_n687), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n636), .A2(KEYINPUT107), .A3(new_n687), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(KEYINPUT108), .B1(new_n682), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n716), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G146), .ZN(G48));
  OR2_X1    g538(.A1(new_n340), .A2(new_n343), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n263), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(G469), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n344), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n355), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n610), .A2(new_n638), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT41), .B(G113), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G15));
  NAND2_X1  g546(.A1(new_n610), .A2(new_n729), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n646), .ZN(new_n734));
  XOR2_X1   g548(.A(KEYINPUT109), .B(G116), .Z(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G18));
  NAND4_X1  g550(.A1(new_n711), .A2(new_n284), .A3(new_n480), .A4(new_n729), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G119), .ZN(G21));
  OAI21_X1  g552(.A(G472), .B1(new_n615), .B2(G902), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n574), .B1(new_n603), .B2(new_n579), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n613), .A2(new_n614), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n740), .B1(new_n742), .B2(new_n675), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n577), .A2(new_n586), .ZN(new_n744));
  OAI211_X1 g558(.A(KEYINPUT110), .B(new_n588), .C1(new_n744), .C2(new_n741), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n739), .A2(new_n743), .A3(new_n530), .A4(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n693), .A2(new_n478), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n747), .A2(new_n286), .A3(new_n748), .A4(new_n729), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G122), .ZN(G24));
  NAND2_X1  g564(.A1(new_n665), .A2(new_n660), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n739), .A2(new_n743), .A3(new_n751), .A4(new_n745), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n753), .A2(new_n715), .A3(new_n279), .A4(new_n729), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n721), .A2(new_n752), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n757), .A2(KEYINPUT111), .A3(new_n279), .A4(new_n729), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G125), .ZN(G27));
  NAND2_X1  g574(.A1(new_n609), .A2(KEYINPUT113), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n587), .A2(new_n762), .A3(KEYINPUT32), .A4(new_n588), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n531), .B1(new_n764), .B2(new_n608), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n277), .A2(new_n187), .A3(new_n278), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n357), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n765), .A2(KEYINPUT42), .A3(new_n715), .A4(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n715), .A2(new_n680), .A3(new_n530), .A4(new_n767), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT42), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT112), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n680), .A2(new_n767), .A3(new_n530), .ZN(new_n772));
  OAI211_X1 g586(.A(KEYINPUT112), .B(new_n770), .C1(new_n772), .C2(new_n721), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n768), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G131), .ZN(G33));
  NAND3_X1  g590(.A1(new_n610), .A2(new_n688), .A3(new_n767), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  NAND2_X1  g592(.A1(new_n348), .A2(new_n349), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT45), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(G469), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT46), .B1(new_n781), .B2(new_n345), .ZN(new_n782));
  INV_X1    g596(.A(new_n344), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n781), .A2(KEYINPUT46), .A3(new_n345), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n355), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n621), .A2(new_n624), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n622), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n693), .A2(new_n634), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT43), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n789), .A2(new_n751), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT44), .ZN(new_n794));
  AOI211_X1 g608(.A(new_n706), .B(new_n787), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n766), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G137), .ZN(G39));
  NAND2_X1  g613(.A1(new_n787), .A2(KEYINPUT47), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n721), .A2(new_n530), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT47), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n786), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n680), .A2(new_n766), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n800), .A2(new_n801), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G140), .ZN(G42));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n792), .A2(new_n683), .ZN(new_n808));
  INV_X1    g622(.A(new_n729), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n808), .A2(new_n809), .A3(new_n766), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n753), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n699), .A2(new_n281), .ZN(new_n812));
  INV_X1    g626(.A(new_n766), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n812), .A2(new_n530), .A3(new_n729), .A4(new_n813), .ZN(new_n814));
  OR3_X1    g628(.A1(new_n814), .A2(new_n445), .A3(new_n634), .ZN(new_n815));
  NOR4_X1   g629(.A1(new_n808), .A2(new_n187), .A3(new_n746), .A4(new_n809), .ZN(new_n816));
  INV_X1    g630(.A(new_n701), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(KEYINPUT50), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT50), .B1(new_n816), .B2(new_n817), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n811), .B(new_n815), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n820), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n818), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n825), .A2(KEYINPUT116), .A3(new_n811), .A4(new_n815), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n800), .A2(new_n803), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n827), .B1(new_n356), .B2(new_n728), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n808), .A2(new_n766), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n747), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n823), .A2(new_n826), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT51), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n807), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n810), .A2(new_n765), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT48), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n257), .A2(G952), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n808), .A2(new_n809), .A3(new_n746), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n836), .B1(new_n837), .B2(new_n279), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n821), .A2(new_n832), .ZN(new_n839));
  INV_X1    g653(.A(new_n830), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n835), .B(new_n838), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n833), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n843));
  INV_X1    g657(.A(new_n734), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n844), .A2(new_n730), .A3(new_n737), .A4(new_n749), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT115), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n625), .A2(new_n639), .ZN(new_n847));
  OR3_X1    g661(.A1(new_n445), .A2(KEYINPUT114), .A3(new_n478), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT114), .B1(new_n445), .B2(new_n478), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n285), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n788), .A2(new_n622), .A3(new_n623), .A4(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n847), .A2(new_n851), .A3(new_n611), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n846), .B1(new_n671), .B2(new_n852), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n668), .A2(KEYINPUT102), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n668), .A2(KEYINPUT102), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n854), .A2(new_n482), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n850), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n611), .B1(new_n625), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(new_n640), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n856), .A2(new_n859), .A3(KEYINPUT115), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n845), .B1(new_n853), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n479), .A2(new_n686), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n680), .A2(new_n645), .A3(new_n667), .A4(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n767), .B1(new_n757), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n775), .A2(new_n777), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n690), .B1(new_n716), .B2(new_n722), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n694), .A2(new_n700), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n751), .A2(new_n686), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n867), .A2(new_n358), .A3(new_n699), .A4(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n759), .A2(new_n866), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT52), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n759), .A2(new_n866), .A3(KEYINPUT52), .A4(new_n869), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n865), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n861), .A2(new_n874), .A3(KEYINPUT53), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT53), .B1(new_n861), .B2(new_n874), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n843), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n872), .A2(new_n873), .ZN(new_n879));
  INV_X1    g693(.A(new_n865), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n845), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n856), .A2(new_n859), .A3(KEYINPUT115), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT115), .B1(new_n856), .B2(new_n859), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n878), .B1(new_n881), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n861), .A2(new_n874), .A3(KEYINPUT53), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n886), .A2(KEYINPUT54), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n877), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n831), .A2(new_n832), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n842), .B(new_n889), .C1(KEYINPUT117), .C2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n814), .A2(new_n637), .ZN(new_n892));
  OAI22_X1  g706(.A1(new_n891), .A2(new_n892), .B1(G952), .B2(G953), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n531), .B1(new_n728), .B2(KEYINPUT49), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n894), .B1(KEYINPUT49), .B2(new_n728), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n895), .A2(new_n701), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n699), .A2(new_n355), .A3(new_n790), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n896), .A2(new_n187), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n893), .A2(new_n898), .ZN(G75));
  AOI21_X1  g713(.A(new_n263), .B1(new_n886), .B2(new_n887), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(G210), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n230), .A2(new_n261), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT118), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT55), .Z(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(new_n259), .ZN(new_n905));
  XOR2_X1   g719(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n906));
  AND3_X1   g720(.A1(new_n901), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT56), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n905), .B1(new_n901), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n257), .A2(G952), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n907), .A2(new_n909), .A3(new_n910), .ZN(G51));
  XNOR2_X1  g725(.A(new_n345), .B(KEYINPUT57), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n725), .B1(new_n889), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n900), .A2(G469), .A3(new_n780), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n910), .B1(new_n913), .B2(new_n914), .ZN(G54));
  NAND3_X1  g729(.A1(new_n900), .A2(KEYINPUT58), .A3(G475), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n916), .A2(new_n423), .A3(new_n428), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n916), .B1(new_n423), .B2(new_n428), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n917), .A2(new_n918), .A3(new_n910), .ZN(G60));
  NAND2_X1  g733(.A1(G478), .A2(G902), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT59), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n877), .A2(new_n888), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n627), .A2(new_n631), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n923), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n877), .A2(new_n888), .A3(new_n927), .A4(new_n921), .ZN(new_n928));
  INV_X1    g742(.A(new_n910), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n922), .A2(KEYINPUT120), .A3(new_n923), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n926), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(KEYINPUT121), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT121), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n926), .A2(new_n930), .A3(new_n934), .A4(new_n931), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n933), .A2(new_n935), .ZN(G63));
  NAND2_X1  g750(.A1(new_n886), .A2(new_n887), .ZN(new_n937));
  NAND2_X1  g751(.A1(G217), .A2(G902), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT60), .Z(new_n939));
  NAND4_X1  g753(.A1(new_n937), .A2(new_n656), .A3(new_n659), .A4(new_n939), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n937), .A2(new_n939), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n940), .B(new_n929), .C1(new_n526), .C2(new_n941), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g757(.A(new_n257), .B1(new_n282), .B2(G224), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n885), .B2(new_n257), .ZN(new_n945));
  INV_X1    g759(.A(G898), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n903), .B1(new_n946), .B2(G953), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n945), .B(new_n947), .ZN(G69));
  NAND3_X1  g762(.A1(new_n558), .A2(new_n563), .A3(new_n566), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n404), .A2(new_n405), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n949), .B(new_n950), .Z(new_n951));
  INV_X1    g765(.A(new_n805), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n797), .B2(new_n795), .ZN(new_n953));
  AOI211_X1 g767(.A(new_n355), .B(new_n706), .C1(new_n784), .C2(new_n785), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n954), .A2(KEYINPUT122), .A3(new_n765), .A4(new_n867), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n955), .A2(new_n759), .A3(new_n866), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT123), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n775), .A2(new_n777), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n775), .A2(KEYINPUT123), .A3(new_n777), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n954), .A2(new_n765), .A3(new_n867), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT122), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n953), .A2(new_n959), .A3(new_n960), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n257), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n257), .A2(G900), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n965), .A2(KEYINPUT124), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(KEYINPUT124), .B1(new_n965), .B2(new_n966), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n951), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n709), .A2(new_n759), .A3(new_n866), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT62), .Z(new_n971));
  NAND3_X1  g785(.A1(new_n848), .A2(new_n637), .A3(new_n849), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n610), .A2(new_n972), .A3(new_n707), .A4(new_n813), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n971), .A2(new_n953), .A3(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n951), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n974), .A2(new_n257), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(G227), .A2(G900), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(G953), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n969), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n978), .B1(new_n969), .B2(new_n976), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(new_n980), .ZN(G72));
  NAND2_X1  g795(.A1(new_n591), .A2(new_n574), .ZN(new_n982));
  NAND2_X1  g796(.A1(G472), .A2(G902), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT126), .Z(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT125), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT63), .Z(new_n986));
  NAND3_X1  g800(.A1(new_n567), .A2(new_n582), .A3(new_n569), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n937), .A2(new_n982), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT127), .Z(new_n989));
  NAND4_X1  g803(.A1(new_n971), .A2(new_n861), .A3(new_n953), .A4(new_n973), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n982), .B1(new_n990), .B2(new_n986), .ZN(new_n991));
  OR2_X1    g805(.A1(new_n964), .A2(new_n885), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n992), .A2(new_n986), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n929), .B1(new_n993), .B2(new_n987), .ZN(new_n994));
  NOR3_X1   g808(.A1(new_n989), .A2(new_n991), .A3(new_n994), .ZN(G57));
endmodule


