//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1254, new_n1255,
    new_n1256, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1322, new_n1323;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  AND2_X1   g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G20), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n203), .A2(G50), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n213), .B1(new_n202), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n201), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n206), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n209), .B1(new_n211), .B2(new_n212), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XOR2_X1   g0025(.A(G250), .B(G257), .Z(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT64), .ZN(new_n227));
  XOR2_X1   g0027(.A(G264), .B(G270), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(new_n219), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n229), .B(new_n233), .Z(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT65), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  INV_X1    g0042(.A(G20), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G33), .ZN(new_n244));
  INV_X1    g0044(.A(G77), .ZN(new_n245));
  OAI22_X1  g0045(.A1(new_n244), .A2(new_n245), .B1(new_n243), .B2(G68), .ZN(new_n246));
  INV_X1    g0046(.A(G33), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n243), .A2(new_n247), .A3(KEYINPUT69), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT69), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n249), .B1(G20), .B2(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n246), .B1(G50), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G1), .A2(G13), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT68), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT68), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n253), .A2(new_n257), .A3(new_n254), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n252), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT11), .ZN(new_n261));
  INV_X1    g0061(.A(G13), .ZN(new_n262));
  NOR3_X1   g0062(.A1(new_n262), .A2(new_n243), .A3(G1), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n263), .B1(new_n256), .B2(new_n258), .ZN(new_n264));
  OAI21_X1  g0064(.A(KEYINPUT70), .B1(new_n243), .B2(G1), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT70), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(new_n267), .A3(G20), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n264), .A2(G68), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n261), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n263), .A2(new_n202), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n272), .B(KEYINPUT12), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n273), .B1(new_n260), .B2(KEYINPUT11), .ZN(new_n274));
  OAI21_X1  g0074(.A(KEYINPUT74), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT12), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n272), .B(new_n276), .ZN(new_n277));
  AND3_X1   g0077(.A1(new_n253), .A2(new_n257), .A3(new_n254), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n257), .B1(new_n253), .B2(new_n254), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n248), .A2(new_n250), .ZN(new_n281));
  INV_X1    g0081(.A(G50), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n280), .B1(new_n283), .B2(new_n246), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT11), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n277), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT74), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n286), .A2(new_n287), .A3(new_n261), .A4(new_n270), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n275), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n219), .A2(G1698), .ZN(new_n290));
  AND2_X1   g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NOR2_X1   g0091(.A1(KEYINPUT3), .A2(G33), .ZN(new_n292));
  OAI221_X1 g0092(.A(new_n290), .B1(G226), .B2(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G97), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n254), .B1(G33), .B2(G41), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G274), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G33), .A2(G41), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n301), .B1(new_n210), .B2(new_n302), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n300), .A2(G238), .B1(new_n299), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT13), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n297), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n210), .A2(new_n302), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n307), .B1(new_n293), .B2(new_n294), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n303), .A2(new_n299), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n307), .A2(new_n298), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n309), .B1(new_n310), .B2(new_n214), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT13), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT14), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n314), .A2(KEYINPUT75), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n313), .A2(G169), .A3(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n306), .A2(new_n312), .A3(G179), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n316), .B1(new_n313), .B2(G169), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT76), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n305), .B1(new_n297), .B2(new_n304), .ZN(new_n322));
  NOR3_X1   g0122(.A1(new_n308), .A2(new_n311), .A3(KEYINPUT13), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G169), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n315), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT76), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n326), .A2(new_n327), .A3(new_n318), .A4(new_n317), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n289), .B1(new_n321), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G190), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n289), .B1(new_n330), .B2(new_n313), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n313), .A2(G200), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT73), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n332), .B(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n329), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT8), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G58), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G150), .ZN(new_n343));
  OAI221_X1 g0143(.A(new_n337), .B1(new_n342), .B2(new_n244), .C1(new_n281), .C2(new_n343), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n344), .A2(new_n280), .B1(new_n282), .B2(new_n263), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n269), .A2(G50), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n346), .B(KEYINPUT71), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n264), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n349), .B(KEYINPUT9), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT3), .B(G33), .ZN(new_n351));
  INV_X1    g0151(.A(G1698), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(G222), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(G223), .A3(G1698), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n353), .B(new_n354), .C1(new_n245), .C2(new_n351), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT67), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n356), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n307), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n309), .ZN(new_n360));
  XOR2_X1   g0160(.A(KEYINPUT66), .B(G226), .Z(new_n361));
  AOI21_X1  g0161(.A(new_n360), .B1(new_n300), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G190), .ZN(new_n365));
  OAI21_X1  g0165(.A(G200), .B1(new_n359), .B2(new_n363), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n350), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT10), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT10), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n350), .A2(new_n369), .A3(new_n365), .A4(new_n366), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n281), .A2(new_n342), .ZN(new_n372));
  XNOR2_X1  g0172(.A(KEYINPUT15), .B(G87), .ZN(new_n373));
  OAI22_X1  g0173(.A1(new_n373), .A2(new_n244), .B1(new_n243), .B2(new_n245), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n280), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n264), .A2(G77), .A3(new_n269), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n262), .A2(G1), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G20), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n375), .B(new_n376), .C1(G77), .C2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n351), .A2(G232), .A3(new_n352), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n351), .A2(G238), .A3(G1698), .ZN(new_n381));
  INV_X1    g0181(.A(G107), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n380), .B(new_n381), .C1(new_n382), .C2(new_n351), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n296), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n360), .B1(G244), .B2(new_n300), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n379), .B1(new_n386), .B2(G200), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n330), .B2(new_n386), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n325), .ZN(new_n389));
  INV_X1    g0189(.A(G179), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n384), .A2(new_n385), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n389), .A2(new_n391), .A3(new_n379), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n364), .A2(new_n390), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n325), .B1(new_n359), .B2(new_n363), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(new_n349), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT72), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT72), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n394), .A2(new_n398), .A3(new_n395), .A4(new_n349), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n393), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g0200(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT7), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n351), .B2(G20), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n291), .A2(new_n292), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n404), .A2(KEYINPUT7), .A3(new_n243), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n202), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  XNOR2_X1  g0206(.A(G58), .B(G68), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n251), .A2(G159), .B1(new_n407), .B2(G20), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n401), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT7), .B1(new_n404), .B2(new_n243), .ZN(new_n411));
  NOR4_X1   g0211(.A1(new_n291), .A2(new_n292), .A3(new_n402), .A4(G20), .ZN(new_n412));
  OAI21_X1  g0212(.A(G68), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n413), .A2(KEYINPUT16), .A3(new_n408), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n410), .A2(new_n414), .A3(new_n280), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT79), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT78), .ZN(new_n417));
  AND3_X1   g0217(.A1(new_n269), .A2(new_n417), .A3(new_n341), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n378), .B1(new_n278), .B2(new_n279), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n417), .B1(new_n269), .B2(new_n341), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n378), .A2(new_n341), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n416), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n420), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n269), .A2(new_n417), .A3(new_n341), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n424), .A2(new_n264), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n422), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(KEYINPUT79), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n415), .A2(new_n423), .A3(new_n428), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n352), .A2(G226), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n351), .B(new_n430), .C1(G223), .C2(G1698), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G87), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n307), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n309), .B1(new_n310), .B2(new_n219), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(G179), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n325), .B2(new_n435), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n429), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT18), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT18), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n429), .A2(new_n440), .A3(new_n437), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n423), .A2(new_n428), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n431), .A2(new_n432), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n296), .ZN(new_n444));
  INV_X1    g0244(.A(new_n434), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(new_n330), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(G200), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(new_n433), .B2(new_n434), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n442), .A2(KEYINPUT17), .A3(new_n415), .A4(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n449), .A2(new_n415), .A3(new_n423), .A4(new_n428), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT17), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n439), .A2(new_n441), .A3(new_n450), .A4(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  AND4_X1   g0255(.A1(new_n336), .A2(new_n371), .A3(new_n400), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G283), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n457), .B(new_n243), .C1(G33), .C2(new_n220), .ZN(new_n458));
  INV_X1    g0258(.A(G116), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G20), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n458), .A2(new_n255), .A3(new_n460), .ZN(new_n461));
  XOR2_X1   g0261(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n462));
  AOI22_X1  g0262(.A1(new_n461), .A2(new_n462), .B1(new_n459), .B2(new_n263), .ZN(new_n463));
  NOR2_X1   g0263(.A1(KEYINPUT83), .A2(KEYINPUT20), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n458), .A2(new_n255), .A3(new_n460), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n267), .A2(G33), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n378), .B(new_n466), .C1(new_n278), .C2(new_n279), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n463), .B(new_n465), .C1(new_n459), .C2(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(G264), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n469));
  OAI211_X1 g0269(.A(G257), .B(new_n352), .C1(new_n291), .C2(new_n292), .ZN(new_n470));
  XNOR2_X1  g0270(.A(KEYINPUT82), .B(G303), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n469), .B(new_n470), .C1(new_n351), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n296), .ZN(new_n473));
  XNOR2_X1  g0273(.A(KEYINPUT5), .B(G41), .ZN(new_n474));
  INV_X1    g0274(.A(G45), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(G1), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n474), .A2(new_n476), .B1(new_n210), .B2(new_n302), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n267), .A2(G45), .ZN(new_n478));
  NOR2_X1   g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(KEYINPUT5), .A2(G41), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n477), .A2(G270), .B1(new_n303), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n473), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n468), .A2(new_n484), .A3(KEYINPUT21), .A4(G169), .ZN(new_n485));
  AND2_X1   g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n476), .B1(new_n486), .B2(new_n479), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(G270), .A3(new_n307), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n303), .A2(new_n476), .A3(new_n474), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n490), .B1(new_n296), .B2(new_n472), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n468), .A2(new_n491), .A3(G179), .ZN(new_n492));
  AND2_X1   g0292(.A1(new_n485), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n325), .B1(new_n473), .B2(new_n483), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n468), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT21), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n463), .A2(new_n465), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n467), .A2(new_n459), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n501), .B(KEYINPUT84), .C1(new_n447), .C2(new_n491), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT84), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n447), .B1(new_n473), .B2(new_n483), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n503), .B1(new_n504), .B2(new_n468), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n491), .A2(G190), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n502), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT85), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT85), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n502), .A2(new_n505), .A3(new_n509), .A4(new_n506), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n498), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n263), .A2(KEYINPUT80), .A3(new_n220), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT80), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n378), .B2(G97), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n512), .B(new_n514), .C1(new_n467), .C2(new_n220), .ZN(new_n515));
  XNOR2_X1  g0315(.A(G97), .B(G107), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT6), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n382), .A2(KEYINPUT6), .A3(G97), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n521), .A2(G20), .B1(G77), .B2(new_n251), .ZN(new_n522));
  OAI21_X1  g0322(.A(G107), .B1(new_n411), .B2(new_n412), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n515), .B1(new_n524), .B2(new_n280), .ZN(new_n525));
  OAI211_X1 g0325(.A(G244), .B(new_n352), .C1(new_n291), .C2(new_n292), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT4), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n351), .A2(KEYINPUT4), .A3(G244), .A4(new_n352), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n351), .A2(G250), .A3(G1698), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n528), .A2(new_n529), .A3(new_n457), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n296), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n487), .A2(new_n307), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n489), .B1(new_n533), .B2(new_n221), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT81), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n489), .B(KEYINPUT81), .C1(new_n533), .C2(new_n221), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n532), .A2(new_n536), .A3(G190), .A4(new_n537), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n532), .A2(new_n536), .A3(new_n537), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n525), .B(new_n538), .C1(new_n539), .C2(new_n447), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n532), .A2(new_n536), .A3(new_n390), .A4(new_n537), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n519), .B1(new_n516), .B2(new_n517), .ZN(new_n542));
  OAI22_X1  g0342(.A1(new_n542), .A2(new_n243), .B1(new_n245), .B2(new_n281), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n382), .B1(new_n403), .B2(new_n405), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n280), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n514), .A2(new_n512), .ZN(new_n546));
  INV_X1    g0346(.A(new_n467), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n546), .B1(new_n547), .B2(G97), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n541), .B(new_n549), .C1(new_n539), .C2(G169), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n540), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n243), .B(G87), .C1(new_n291), .C2(new_n292), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT22), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT22), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n351), .A2(new_n554), .A3(new_n243), .A4(G87), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n382), .A2(KEYINPUT23), .A3(G20), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT23), .B1(new_n382), .B2(G20), .ZN(new_n558));
  NAND2_X1  g0358(.A1(G33), .A2(G116), .ZN(new_n559));
  OAI22_X1  g0359(.A1(new_n557), .A2(new_n558), .B1(G20), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT24), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n560), .B1(new_n553), .B2(new_n555), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT24), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n280), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT86), .ZN(new_n568));
  OR2_X1    g0368(.A1(new_n568), .A2(KEYINPUT25), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n243), .A2(G107), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(KEYINPUT25), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n569), .A2(new_n377), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n377), .A2(new_n570), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n572), .B1(new_n573), .B2(new_n571), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n547), .B2(G107), .ZN(new_n575));
  OAI211_X1 g0375(.A(G257), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n576));
  OAI211_X1 g0376(.A(G250), .B(new_n352), .C1(new_n291), .C2(new_n292), .ZN(new_n577));
  NAND2_X1  g0377(.A1(G33), .A2(G294), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n579), .A2(new_n296), .B1(new_n477), .B2(G264), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n580), .A2(new_n330), .A3(new_n489), .ZN(new_n581));
  AOI21_X1  g0381(.A(G200), .B1(new_n580), .B2(new_n489), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n567), .B(new_n575), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n280), .B1(new_n565), .B2(KEYINPUT24), .ZN(new_n584));
  AOI211_X1 g0384(.A(new_n563), .B(new_n560), .C1(new_n553), .C2(new_n555), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n575), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n580), .A2(new_n390), .A3(new_n489), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n580), .A2(new_n489), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n325), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n583), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n373), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n259), .A2(new_n378), .A3(new_n592), .A4(new_n466), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT19), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n243), .B1(new_n294), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n215), .A2(new_n220), .A3(new_n382), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n243), .B(G68), .C1(new_n291), .C2(new_n292), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n594), .B1(new_n244), .B2(new_n220), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n280), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n373), .A2(new_n263), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n593), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n303), .A2(new_n476), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n216), .B1(new_n267), .B2(G45), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n307), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n214), .A2(new_n352), .ZN(new_n608));
  INV_X1    g0408(.A(G244), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(G1698), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n608), .B(new_n610), .C1(new_n291), .C2(new_n292), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n307), .B1(new_n611), .B2(new_n559), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n325), .B1(new_n607), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n559), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n296), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n303), .A2(new_n476), .B1(new_n307), .B2(new_n605), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n390), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n603), .A2(new_n613), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(G200), .B1(new_n607), .B2(new_n612), .ZN(new_n619));
  NOR2_X1   g0419(.A1(G238), .A2(G1698), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n620), .B1(new_n609), .B2(G1698), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n621), .A2(new_n351), .B1(G33), .B2(G116), .ZN(new_n622));
  OAI211_X1 g0422(.A(G190), .B(new_n616), .C1(new_n622), .C2(new_n307), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n600), .A2(new_n280), .B1(new_n263), .B2(new_n373), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n264), .A2(G87), .A3(new_n466), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n619), .A2(new_n623), .A3(new_n624), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n618), .A2(new_n626), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n551), .A2(new_n591), .A3(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n456), .A2(new_n511), .A3(new_n628), .ZN(G372));
  INV_X1    g0429(.A(KEYINPUT87), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n618), .A2(new_n630), .A3(new_n626), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n630), .B1(new_n618), .B2(new_n626), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n633), .A2(new_n583), .A3(new_n550), .A4(new_n540), .ZN(new_n634));
  INV_X1    g0434(.A(new_n590), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n485), .A2(new_n492), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT21), .B1(new_n494), .B2(new_n468), .ZN(new_n637));
  OAI21_X1  g0437(.A(KEYINPUT88), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT88), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n497), .A2(new_n639), .A3(new_n492), .A4(new_n485), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n635), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n634), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(KEYINPUT26), .B1(new_n550), .B2(new_n627), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n627), .A2(KEYINPUT87), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n532), .A2(new_n536), .A3(new_n537), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n645), .A2(new_n325), .B1(new_n545), .B2(new_n548), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n618), .A2(new_n630), .A3(new_n626), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n644), .A2(new_n541), .A3(new_n646), .A4(new_n647), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n618), .B(new_n643), .C1(new_n648), .C2(KEYINPUT26), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n642), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n456), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g0451(.A(new_n651), .B(KEYINPUT89), .Z(new_n652));
  NOR2_X1   g0452(.A1(new_n335), .A2(new_n392), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n453), .B(new_n450), .C1(new_n653), .C2(new_n329), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n654), .A2(new_n439), .A3(new_n441), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n655), .A2(new_n371), .B1(new_n397), .B2(new_n399), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n652), .A2(new_n656), .ZN(G369));
  INV_X1    g0457(.A(G330), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n377), .A2(new_n243), .ZN(new_n659));
  AOI21_X1  g0459(.A(KEYINPUT90), .B1(new_n659), .B2(KEYINPUT27), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n659), .A2(KEYINPUT90), .A3(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(G213), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g0465(.A(KEYINPUT91), .B(G343), .Z(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(new_n501), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n511), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n638), .A2(new_n640), .A3(new_n669), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n658), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n586), .A2(new_n667), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n583), .A2(new_n590), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT92), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n583), .A2(new_n590), .A3(KEYINPUT92), .A4(new_n674), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n635), .A2(new_n667), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n673), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n635), .A2(new_n668), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n667), .B1(new_n493), .B2(new_n497), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n677), .A2(new_n678), .A3(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n682), .A2(new_n683), .A3(new_n685), .ZN(G399));
  INV_X1    g0486(.A(new_n207), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(G41), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n596), .A2(G116), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G1), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n212), .B2(new_n689), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT28), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT29), .ZN(new_n694));
  OAI211_X1 g0494(.A(new_n694), .B(new_n668), .C1(new_n642), .C2(new_n649), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n618), .A2(new_n626), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT26), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n696), .A2(new_n646), .A3(new_n697), .A4(new_n541), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n618), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n699), .B1(KEYINPUT26), .B2(new_n648), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n549), .B1(G200), .B2(new_n645), .ZN(new_n701));
  AOI22_X1  g0501(.A1(new_n701), .A2(new_n538), .B1(new_n646), .B2(new_n541), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n493), .A2(new_n497), .A3(new_n590), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n702), .A2(new_n703), .A3(new_n633), .A4(new_n583), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n667), .B1(new_n700), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n695), .B1(new_n705), .B2(new_n694), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT93), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n390), .B1(new_n607), .B2(new_n612), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n707), .B1(new_n491), .B2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(G179), .B1(new_n615), .B2(new_n616), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n484), .A2(new_n710), .A3(KEYINPUT93), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n709), .A2(new_n588), .A3(new_n645), .A4(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n607), .A2(new_n612), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n491), .A2(G179), .A3(new_n580), .A4(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n713), .B1(new_n715), .B2(new_n645), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n484), .A2(new_n390), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n580), .A2(new_n714), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n539), .A2(KEYINPUT30), .A3(new_n717), .A4(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n712), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n667), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT31), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n720), .A2(KEYINPUT31), .A3(new_n667), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n628), .A2(new_n511), .A3(new_n668), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n658), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT94), .B1(new_n706), .B2(new_n728), .ZN(new_n729));
  AND3_X1   g0529(.A1(new_n628), .A2(new_n511), .A3(new_n668), .ZN(new_n730));
  OAI21_X1  g0530(.A(G330), .B1(new_n730), .B2(new_n725), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n698), .A2(new_n618), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n648), .A2(KEYINPUT26), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n704), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n668), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT29), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT94), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n731), .A2(new_n736), .A3(new_n737), .A4(new_n695), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n729), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n693), .B1(new_n739), .B2(G1), .ZN(G364));
  NOR2_X1   g0540(.A1(new_n262), .A2(G20), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n267), .B1(new_n741), .B2(G45), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n688), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n673), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n672), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(new_n511), .B2(new_n670), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n745), .B1(G330), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G13), .A2(G33), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n254), .B1(G20), .B2(new_n325), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n241), .A2(G45), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT95), .Z(new_n757));
  NOR2_X1   g0557(.A1(new_n687), .A2(new_n351), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n757), .B(new_n758), .C1(G45), .C2(new_n212), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n687), .A2(new_n404), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n760), .A2(G355), .B1(new_n459), .B2(new_n687), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n755), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n753), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n390), .A2(G200), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n764), .A2(G20), .A3(G190), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n351), .B1(new_n765), .B2(new_n201), .ZN(new_n766));
  NOR4_X1   g0566(.A1(new_n243), .A2(new_n330), .A3(new_n447), .A4(G179), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n330), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n768), .A2(new_n215), .B1(new_n282), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n243), .A2(G190), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(new_n764), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n766), .B(new_n772), .C1(G77), .C2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G179), .A2(G200), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n243), .B1(new_n777), .B2(G190), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT97), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G97), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n773), .A2(new_n777), .ZN(new_n781));
  INV_X1    g0581(.A(G159), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  XOR2_X1   g0584(.A(KEYINPUT96), .B(KEYINPUT32), .Z(new_n785));
  NOR4_X1   g0585(.A1(new_n243), .A2(new_n447), .A3(G179), .A4(G190), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n784), .A2(new_n785), .B1(G107), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n785), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n769), .A2(G190), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n783), .A2(new_n788), .B1(G68), .B2(new_n789), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n776), .A2(new_n780), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G322), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n765), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G311), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n404), .B1(new_n774), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n781), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n793), .B(new_n795), .C1(G329), .C2(new_n796), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT98), .B(G326), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n771), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(KEYINPUT33), .B(G317), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n767), .A2(G303), .B1(new_n789), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n778), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n802), .A2(G294), .B1(new_n786), .B2(G283), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n797), .A2(new_n799), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n763), .B1(new_n791), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n744), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n762), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n752), .B(KEYINPUT99), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n748), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n749), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(G396));
  NAND2_X1  g0611(.A1(new_n650), .A2(new_n668), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n667), .A2(new_n379), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n388), .A2(new_n392), .A3(new_n813), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n389), .A2(new_n667), .A3(new_n391), .A4(new_n379), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(KEYINPUT102), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n815), .A2(KEYINPUT102), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n814), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n812), .A2(new_n820), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n668), .B(new_n819), .C1(new_n642), .C2(new_n649), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n744), .B1(new_n823), .B2(new_n731), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n731), .B2(new_n823), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n774), .A2(new_n459), .B1(new_n781), .B2(new_n794), .ZN(new_n826));
  INV_X1    g0626(.A(new_n765), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n351), .B(new_n826), .C1(G294), .C2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n786), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(new_n215), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(G303), .B2(new_n770), .ZN(new_n831));
  XNOR2_X1  g0631(.A(KEYINPUT100), .B(G283), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G107), .A2(new_n767), .B1(new_n833), .B2(new_n789), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n828), .A2(new_n780), .A3(new_n831), .A4(new_n834), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n827), .A2(G143), .B1(new_n775), .B2(G159), .ZN(new_n836));
  INV_X1    g0636(.A(G137), .ZN(new_n837));
  INV_X1    g0637(.A(new_n789), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n836), .B1(new_n771), .B2(new_n837), .C1(new_n343), .C2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT34), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(G132), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n351), .B1(new_n781), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G68), .B2(new_n786), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n767), .A2(G50), .B1(new_n802), .B2(G58), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n841), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n839), .A2(new_n840), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n835), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT101), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n763), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n849), .B2(new_n848), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n753), .A2(new_n750), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n806), .B1(new_n245), .B2(new_n852), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n851), .B(new_n853), .C1(new_n819), .C2(new_n751), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n825), .A2(new_n854), .ZN(G384));
  NOR2_X1   g0655(.A1(new_n741), .A2(new_n267), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n289), .A2(new_n668), .ZN(new_n857));
  NOR3_X1   g0657(.A1(new_n329), .A2(new_n335), .A3(new_n857), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n329), .A2(new_n667), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n819), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n724), .A2(KEYINPUT106), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT106), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n720), .A2(new_n862), .A3(KEYINPUT31), .A4(new_n667), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n727), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT105), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT31), .B1(new_n721), .B2(KEYINPUT104), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT104), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n720), .A2(new_n868), .A3(new_n667), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n866), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n867), .A2(new_n866), .A3(new_n869), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n860), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n421), .A2(new_n422), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n415), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n665), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n454), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n429), .A2(new_n876), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT37), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n438), .A2(new_n880), .A3(new_n881), .A4(new_n451), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n875), .A2(new_n437), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n883), .A2(new_n877), .A3(new_n451), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n882), .B1(new_n884), .B2(new_n881), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n879), .A2(KEYINPUT38), .A3(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n880), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n454), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n438), .A2(new_n880), .A3(new_n451), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT37), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n882), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT38), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT107), .B1(new_n886), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n879), .A2(KEYINPUT38), .A3(new_n885), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT107), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n454), .A2(new_n887), .B1(new_n890), .B2(new_n882), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n894), .B(new_n895), .C1(new_n896), .C2(KEYINPUT38), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n873), .A2(KEYINPUT40), .A3(new_n893), .A4(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT40), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n721), .A2(KEYINPUT104), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(new_n722), .A3(new_n869), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT105), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n902), .A2(new_n727), .A3(new_n872), .A4(new_n864), .ZN(new_n903));
  INV_X1    g0703(.A(new_n329), .ZN(new_n904));
  INV_X1    g0704(.A(new_n335), .ZN(new_n905));
  INV_X1    g0705(.A(new_n857), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n329), .A2(new_n667), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n820), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n903), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n879), .A2(new_n885), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT38), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n894), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n899), .B1(new_n910), .B2(new_n915), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n898), .A2(new_n916), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n903), .A2(new_n456), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n658), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n917), .B2(new_n918), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n858), .A2(new_n859), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n392), .A2(new_n667), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n921), .B1(new_n822), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n914), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT39), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n886), .B2(new_n892), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n913), .A2(KEYINPUT39), .A3(new_n894), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n329), .A2(new_n668), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n439), .ZN(new_n931));
  INV_X1    g0731(.A(new_n441), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n665), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n924), .A2(new_n930), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n706), .A2(new_n456), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n656), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n934), .B(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n856), .B1(new_n920), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n937), .B2(new_n920), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n521), .A2(KEYINPUT35), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n211), .A2(new_n459), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n521), .B2(KEYINPUT35), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT103), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n943), .B2(new_n942), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT36), .Z(new_n946));
  OAI21_X1  g0746(.A(G77), .B1(new_n201), .B2(new_n202), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n212), .A2(new_n947), .B1(G50), .B2(new_n202), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n948), .A2(G1), .A3(new_n262), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n939), .A2(new_n946), .A3(new_n949), .ZN(G367));
  NAND2_X1  g0750(.A1(new_n624), .A2(new_n625), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n667), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n952), .A2(new_n618), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n633), .B2(new_n952), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT43), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n702), .B(new_n635), .C1(new_n525), .C2(new_n668), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n667), .B1(new_n957), .B2(new_n550), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n668), .A2(new_n525), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n551), .A2(new_n959), .B1(new_n550), .B2(new_n668), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n960), .A2(new_n677), .A3(new_n678), .A4(new_n684), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n958), .B1(KEYINPUT42), .B2(new_n961), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n961), .A2(KEYINPUT42), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n956), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n954), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n964), .B1(KEYINPUT43), .B2(new_n965), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n962), .A2(new_n963), .A3(new_n955), .A4(new_n954), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n960), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n682), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n968), .B(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n688), .B(KEYINPUT41), .Z(new_n972));
  INV_X1    g0772(.A(new_n684), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n679), .A2(new_n680), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n685), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n673), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n685), .B(new_n974), .C1(new_n747), .C2(new_n658), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n729), .B2(new_n738), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n685), .A2(new_n683), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n969), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(KEYINPUT108), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT108), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n980), .A2(new_n983), .A3(new_n969), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n982), .A2(KEYINPUT44), .A3(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT44), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n983), .B1(new_n980), .B2(new_n969), .ZN(new_n987));
  AOI211_X1 g0787(.A(KEYINPUT108), .B(new_n960), .C1(new_n685), .C2(new_n683), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n685), .A2(new_n683), .A3(new_n960), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT45), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n985), .A2(new_n989), .A3(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n682), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n985), .A2(new_n989), .A3(new_n682), .A4(new_n992), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n979), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n972), .B1(new_n997), .B2(new_n739), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n971), .B1(new_n998), .B2(new_n743), .ZN(new_n999));
  INV_X1    g0799(.A(new_n758), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n229), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n754), .B1(new_n207), .B2(new_n373), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n744), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n774), .A2(new_n282), .B1(new_n781), .B2(new_n837), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n404), .B(new_n1004), .C1(G150), .C2(new_n827), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n779), .A2(G68), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n829), .A2(new_n245), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(G159), .B2(new_n789), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n767), .A2(G58), .B1(G143), .B2(new_n770), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1005), .A2(new_n1006), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n829), .A2(new_n220), .ZN(new_n1011));
  INV_X1    g0811(.A(G317), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n404), .B1(new_n781), .B2(new_n1012), .C1(new_n774), .C2(new_n832), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1011), .B(new_n1013), .C1(G107), .C2(new_n802), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT46), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n768), .B2(new_n459), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n767), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1017));
  INV_X1    g0817(.A(G294), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1016), .B(new_n1017), .C1(new_n1018), .C2(new_n838), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT110), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n771), .A2(new_n794), .B1(new_n765), .B2(new_n471), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1022), .A2(KEYINPUT109), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(KEYINPUT109), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1014), .A2(new_n1021), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1010), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT47), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1003), .B1(new_n1028), .B2(new_n753), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n808), .B2(new_n965), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n999), .A2(new_n1030), .ZN(G387));
  INV_X1    g0831(.A(new_n978), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n739), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n729), .A2(new_n738), .A3(new_n978), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n688), .B(KEYINPUT113), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n681), .A2(new_n808), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n690), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n760), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(G107), .B2(new_n207), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1000), .B1(new_n233), .B2(G45), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n475), .B1(new_n202), .B2(new_n245), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT111), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1042), .B1(new_n1038), .B2(new_n1043), .ZN(new_n1044));
  AND3_X1   g0844(.A1(new_n341), .A2(KEYINPUT50), .A3(new_n282), .ZN(new_n1045));
  AOI21_X1  g0845(.A(KEYINPUT50), .B1(new_n341), .B2(new_n282), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1044), .B1(new_n1043), .B2(new_n1038), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1040), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n744), .B1(new_n1048), .B2(new_n755), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n765), .A2(new_n282), .B1(new_n774), .B2(new_n202), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n404), .B(new_n1050), .C1(G150), .C2(new_n796), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n779), .A2(new_n592), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1011), .B1(G159), .B2(new_n770), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n767), .A2(G77), .B1(new_n341), .B2(new_n789), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT112), .Z(new_n1056));
  NOR2_X1   g0856(.A1(new_n774), .A2(new_n471), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G317), .B2(new_n827), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n794), .B2(new_n838), .C1(new_n792), .C2(new_n771), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT48), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n767), .A2(G294), .B1(new_n802), .B2(new_n833), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT49), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n404), .B1(new_n781), .B2(new_n798), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(G116), .B2(new_n786), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1056), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1049), .B1(new_n1070), .B2(new_n753), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1032), .A2(new_n743), .B1(new_n1037), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1036), .A2(new_n1072), .ZN(G393));
  NAND2_X1  g0873(.A1(new_n995), .A2(new_n996), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n1033), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1075), .A2(new_n997), .A3(new_n1035), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n995), .A2(new_n743), .A3(new_n996), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n238), .A2(new_n758), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n754), .B1(new_n220), .B2(new_n207), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n744), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n771), .A2(new_n1012), .B1(new_n765), .B2(new_n794), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1081), .B(new_n1082), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n404), .B1(new_n781), .B2(new_n792), .C1(new_n1018), .C2(new_n774), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n829), .A2(new_n382), .B1(new_n471), .B2(new_n838), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n768), .A2(new_n832), .B1(new_n459), .B2(new_n778), .ZN(new_n1086));
  NOR4_X1   g0886(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .A4(new_n1086), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT117), .Z(new_n1088));
  INV_X1    g0888(.A(G143), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n351), .B1(new_n781), .B2(new_n1089), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1090), .B(new_n830), .C1(G68), .C2(new_n767), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n771), .A2(new_n343), .B1(new_n765), .B2(new_n782), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT51), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n779), .A2(G77), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n342), .A2(new_n774), .B1(new_n838), .B2(new_n282), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT114), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1091), .A2(new_n1093), .A3(new_n1094), .A4(new_n1096), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n1097), .A2(KEYINPUT115), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(KEYINPUT115), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1088), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1080), .B1(new_n1100), .B2(new_n753), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n752), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1101), .B1(new_n1102), .B2(new_n960), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n1077), .A2(KEYINPUT118), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(KEYINPUT118), .B1(new_n1077), .B2(new_n1103), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1076), .B1(new_n1104), .B2(new_n1105), .ZN(G390));
  NAND2_X1  g0906(.A1(new_n926), .A2(new_n927), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n750), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1094), .B1(new_n459), .B2(new_n765), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT120), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n404), .B1(new_n781), .B2(new_n1018), .C1(new_n220), .C2(new_n774), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n768), .A2(new_n215), .B1(new_n829), .B2(new_n202), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n770), .A2(G283), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n838), .B2(new_n382), .ZN(new_n1114));
  NOR4_X1   g0914(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .A4(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(G128), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n771), .A2(new_n1116), .B1(new_n765), .B2(new_n842), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT119), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n779), .A2(G159), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n1118), .B2(new_n1117), .ZN(new_n1120));
  INV_X1    g0920(.A(G125), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT54), .B(G143), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n351), .B1(new_n781), .B2(new_n1121), .C1(new_n774), .C2(new_n1122), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n829), .A2(new_n282), .B1(new_n837), .B2(new_n838), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n767), .A2(G150), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT53), .ZN(new_n1126));
  NOR4_X1   g0926(.A1(new_n1120), .A2(new_n1123), .A3(new_n1124), .A4(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n753), .B1(new_n1115), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n806), .B1(new_n342), .B2(new_n852), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1108), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n903), .A2(G330), .A3(new_n909), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n734), .A2(new_n668), .A3(new_n819), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n922), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n907), .A2(new_n908), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AND4_X1   g0936(.A1(new_n928), .A2(new_n1136), .A3(new_n893), .A4(new_n897), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n822), .A2(new_n922), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n1135), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1139), .A2(new_n928), .B1(new_n926), .B2(new_n927), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1132), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1107), .B1(new_n923), .B2(new_n929), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1136), .A2(new_n893), .A3(new_n928), .A4(new_n897), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n731), .A2(new_n820), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n1135), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1142), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1141), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1130), .B1(new_n1147), .B2(new_n742), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n921), .B1(new_n731), .B2(new_n820), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1131), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n1138), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n903), .A2(G330), .A3(new_n819), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n921), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1134), .B1(new_n1144), .B2(new_n1135), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n903), .A2(new_n456), .A3(G330), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n656), .A2(new_n1157), .A3(new_n935), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1156), .A2(new_n1141), .A3(new_n1146), .A4(new_n1159), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n1160), .A2(new_n1035), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n1147), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1148), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(G378));
  AND2_X1   g0965(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1159), .B1(new_n1147), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n349), .A2(new_n876), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n371), .B2(new_n396), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n371), .A2(new_n396), .A3(new_n1168), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1172), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n371), .A2(new_n396), .A3(new_n1168), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1174), .B1(new_n1175), .B2(new_n1169), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n893), .A2(KEYINPUT40), .A3(new_n897), .ZN(new_n1178));
  OAI21_X1  g0978(.A(G330), .B1(new_n1178), .B2(new_n910), .ZN(new_n1179));
  AOI21_X1  g0979(.A(KEYINPUT40), .B1(new_n873), .B2(new_n914), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1177), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n898), .A2(new_n1182), .A3(new_n916), .A4(G330), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n934), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n934), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1181), .A2(new_n1183), .A3(new_n1186), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1167), .A2(new_n1185), .A3(KEYINPUT57), .A4(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n934), .A2(KEYINPUT122), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1184), .A2(new_n1189), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n934), .A2(KEYINPUT122), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1191), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1190), .A2(new_n1192), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1035), .B(new_n1188), .C1(new_n1193), .C2(KEYINPUT57), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1182), .A2(new_n750), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n852), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n744), .B1(G50), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n282), .B1(G33), .B2(G41), .ZN(new_n1199));
  INV_X1    g0999(.A(G41), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1199), .B1(new_n404), .B2(new_n1200), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n838), .A2(new_n220), .B1(new_n771), .B2(new_n459), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n829), .A2(new_n201), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1202), .B(new_n1203), .C1(G77), .C2(new_n767), .ZN(new_n1204));
  AOI211_X1 g1004(.A(G41), .B(new_n351), .C1(new_n796), .C2(G283), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n827), .A2(G107), .B1(new_n775), .B2(new_n592), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1204), .A2(new_n1006), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT58), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1201), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n768), .A2(new_n1122), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT121), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n838), .A2(new_n842), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n765), .A2(new_n1116), .B1(new_n774), .B2(new_n837), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(G125), .C2(new_n770), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n779), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1211), .B(new_n1214), .C1(new_n343), .C2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(KEYINPUT59), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n786), .A2(G159), .ZN(new_n1218));
  AOI211_X1 g1018(.A(G33), .B(G41), .C1(new_n796), .C2(G124), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1216), .A2(KEYINPUT59), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1209), .B1(new_n1208), .B2(new_n1207), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1198), .B1(new_n1222), .B2(new_n753), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1195), .A2(new_n743), .B1(new_n1196), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1194), .A2(new_n1224), .ZN(G375));
  INV_X1    g1025(.A(new_n972), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1151), .A2(new_n1155), .A3(new_n1158), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1162), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n768), .A2(new_n220), .B1(new_n1018), .B2(new_n771), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1007), .B(new_n1229), .C1(G116), .C2(new_n789), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n351), .B1(new_n827), .B2(G283), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n775), .A2(G107), .B1(new_n796), .B2(G303), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1230), .A2(new_n1052), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT123), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n842), .A2(new_n771), .B1(new_n838), .B2(new_n1122), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n1236), .B(new_n1203), .C1(G159), .C2(new_n767), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n765), .A2(new_n837), .B1(new_n781), .B2(new_n1116), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n404), .B(new_n1238), .C1(G150), .C2(new_n775), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1237), .B(new_n1239), .C1(new_n282), .C2(new_n1215), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1235), .A2(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n753), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1243), .B(new_n744), .C1(G68), .C2(new_n1197), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n921), .B2(new_n750), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(new_n1156), .B2(new_n743), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1228), .A2(new_n1246), .ZN(G381));
  NAND3_X1  g1047(.A1(new_n1036), .A2(new_n810), .A3(new_n1072), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(G384), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  OR3_X1    g1051(.A1(new_n1251), .A2(G381), .A3(G390), .ZN(new_n1252));
  OR4_X1    g1052(.A1(G387), .A2(G375), .A3(G378), .A4(new_n1252), .ZN(G407));
  NAND2_X1  g1053(.A1(new_n666), .A2(G213), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1164), .A2(new_n1255), .ZN(new_n1256));
  OAI211_X1 g1056(.A(G407), .B(G213), .C1(G375), .C2(new_n1256), .ZN(G409));
  NAND3_X1  g1057(.A1(G390), .A2(new_n999), .A3(new_n1030), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(KEYINPUT125), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n810), .B1(new_n1036), .B2(new_n1072), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT124), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(new_n1249), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G393), .A2(G396), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT124), .B1(new_n1263), .B2(new_n1248), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1259), .A2(new_n1265), .ZN(new_n1266));
  OR2_X1    g1066(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(G387), .A2(new_n1267), .A3(new_n1076), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1258), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1266), .A2(new_n1269), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1259), .A2(new_n1265), .A3(new_n1268), .A4(new_n1258), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1194), .A2(G378), .A3(new_n1224), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1192), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1191), .B1(new_n1183), .B2(new_n1181), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1226), .B(new_n1167), .C1(new_n1274), .C2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1196), .A2(new_n1223), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1185), .A2(new_n743), .A3(new_n1187), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1276), .A2(new_n1277), .A3(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1164), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1273), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1254), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1255), .A2(G2897), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1166), .A2(KEYINPUT60), .A3(new_n1158), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT60), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1227), .A2(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1285), .A2(new_n1035), .A3(new_n1162), .A4(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1288), .A2(G384), .A3(new_n1246), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(G384), .B1(new_n1288), .B2(new_n1246), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1284), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1291), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1293), .A2(new_n1289), .A3(new_n1283), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT61), .B1(new_n1282), .B2(new_n1295), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1281), .A2(new_n1254), .A3(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(KEYINPUT62), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1296), .A2(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1298), .A2(KEYINPUT62), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1272), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT63), .ZN(new_n1303));
  NOR3_X1   g1103(.A1(new_n1290), .A2(new_n1291), .A3(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1281), .A2(new_n1254), .A3(new_n1304), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1266), .A2(new_n1269), .ZN(new_n1306));
  AOI22_X1  g1106(.A1(new_n1259), .A2(new_n1265), .B1(new_n1268), .B2(new_n1258), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1305), .A2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1255), .B1(new_n1273), .B2(new_n1280), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT63), .B1(new_n1310), .B2(new_n1297), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1309), .A2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(KEYINPUT126), .B1(new_n1312), .B2(new_n1296), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1272), .B1(new_n1310), .B2(new_n1304), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1298), .A2(new_n1303), .ZN(new_n1315));
  AND4_X1   g1115(.A1(KEYINPUT126), .A2(new_n1296), .A3(new_n1314), .A4(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1302), .B1(new_n1313), .B2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT127), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  OAI211_X1 g1119(.A(KEYINPUT127), .B(new_n1302), .C1(new_n1313), .C2(new_n1316), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(G405));
  XNOR2_X1  g1121(.A(G375), .B(G378), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(new_n1322), .B(new_n1297), .ZN(new_n1323));
  XNOR2_X1  g1123(.A(new_n1323), .B(new_n1308), .ZN(G402));
endmodule


