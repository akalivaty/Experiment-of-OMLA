//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  INV_X1    g001(.A(G197gat), .ZN(new_n203));
  INV_X1    g002(.A(G204gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G197gat), .A2(G204gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G211gat), .A2(G218gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT22), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G211gat), .B(G218gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(KEYINPUT73), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n212), .ZN(new_n214));
  AOI22_X1  g013(.A1(new_n205), .A2(new_n206), .B1(new_n209), .B2(new_n208), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT73), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  AND2_X1   g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n219), .B1(new_n220), .B2(KEYINPUT24), .ZN(new_n221));
  NAND2_X1  g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223));
  AND3_X1   g022(.A1(new_n222), .A2(KEYINPUT66), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT66), .B1(new_n222), .B2(new_n223), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n221), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT67), .ZN(new_n227));
  NOR2_X1   g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n228), .B1(KEYINPUT23), .B2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n230), .B1(KEYINPUT23), .B2(new_n228), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT67), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n221), .B(new_n232), .C1(new_n224), .C2(new_n225), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n227), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT25), .ZN(new_n235));
  NAND3_X1  g034(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(G183gat), .B2(G190gat), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n238));
  AND2_X1   g037(.A1(new_n229), .A2(KEYINPUT23), .ZN(new_n239));
  OAI22_X1  g038(.A1(new_n237), .A2(new_n238), .B1(new_n239), .B2(new_n228), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT25), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT65), .B(G169gat), .ZN(new_n242));
  INV_X1    g041(.A(G176gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT23), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n241), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT28), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT27), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(new_n249), .A3(G183gat), .ZN(new_n250));
  INV_X1    g049(.A(G190gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n249), .B1(new_n248), .B2(G183gat), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n247), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT27), .B(G183gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(KEYINPUT28), .A3(new_n251), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n220), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT26), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n229), .A2(new_n258), .ZN(new_n259));
  NOR3_X1   g058(.A1(KEYINPUT69), .A2(G169gat), .A3(G176gat), .ZN(new_n260));
  MUX2_X1   g059(.A(new_n259), .B(new_n258), .S(new_n260), .Z(new_n261));
  AOI21_X1  g060(.A(new_n246), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G226gat), .A2(G233gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(KEYINPUT74), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n235), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT29), .ZN(new_n266));
  AOI22_X1  g065(.A1(new_n235), .A2(new_n262), .B1(new_n266), .B2(new_n264), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n218), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n235), .A2(new_n262), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n264), .A2(new_n266), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n218), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n235), .A2(new_n262), .A3(new_n264), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT75), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n268), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  OAI211_X1 g075(.A(KEYINPUT75), .B(new_n218), .C1(new_n265), .C2(new_n267), .ZN(new_n277));
  XNOR2_X1  g076(.A(G64gat), .B(G92gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT76), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(G8gat), .ZN(new_n280));
  INV_X1    g079(.A(G36gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  AND3_X1   g082(.A1(new_n276), .A2(new_n277), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n283), .B1(new_n276), .B2(new_n277), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n284), .B1(KEYINPUT30), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G22gat), .B(G50gat), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT2), .ZN(new_n289));
  INV_X1    g088(.A(G148gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G141gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n290), .A2(G141gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n289), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(G155gat), .A2(G162gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT78), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(new_n290), .B2(G141gat), .ZN(new_n299));
  INV_X1    g098(.A(G141gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n300), .A2(KEYINPUT78), .A3(G148gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n291), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303));
  INV_X1    g102(.A(G155gat), .ZN(new_n304));
  INV_X1    g103(.A(G162gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n303), .B1(new_n306), .B2(KEYINPUT2), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n294), .A2(new_n297), .B1(new_n302), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n213), .A2(new_n217), .A3(new_n266), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT3), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT86), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n302), .A2(new_n307), .ZN(new_n314));
  XNOR2_X1  g113(.A(G141gat), .B(G148gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n297), .B1(new_n315), .B2(KEYINPUT2), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(new_n316), .A3(new_n310), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(new_n266), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n218), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n314), .A2(new_n316), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT3), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n321), .B(KEYINPUT86), .C1(new_n309), .C2(new_n308), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n313), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  AND2_X1   g122(.A1(G228gat), .A2(G233gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G78gat), .B(G106gat), .ZN(new_n326));
  XOR2_X1   g125(.A(new_n326), .B(KEYINPUT31), .Z(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT29), .B1(new_n214), .B2(new_n215), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n211), .A2(new_n212), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(new_n310), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n324), .B1(new_n332), .B2(new_n320), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n319), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n325), .A2(new_n328), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n328), .B1(new_n325), .B2(new_n334), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n288), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n337), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n339), .A2(new_n287), .A3(new_n335), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT77), .B1(new_n285), .B2(KEYINPUT30), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n276), .A2(new_n277), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(new_n282), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT77), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT30), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AND4_X1   g146(.A1(new_n286), .A2(new_n341), .A3(new_n342), .A4(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(G134gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G127gat), .ZN(new_n350));
  INV_X1    g149(.A(G127gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G134gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G113gat), .B(G120gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n353), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(G120gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G113gat), .ZN(new_n359));
  INV_X1    g158(.A(G113gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(G120gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G127gat), .B(G134gat), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(new_n363), .A3(new_n355), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n357), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n269), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n365), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n235), .A2(new_n262), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G227gat), .ZN(new_n370));
  INV_X1    g169(.A(G233gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT34), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  XOR2_X1   g172(.A(new_n372), .B(KEYINPUT64), .Z(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n375), .A2(KEYINPUT34), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n366), .A2(new_n368), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G15gat), .B(G43gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(G71gat), .B(G99gat), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n379), .B(new_n380), .Z(new_n381));
  AOI21_X1  g180(.A(new_n374), .B1(new_n366), .B2(new_n368), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n381), .B1(new_n382), .B2(KEYINPUT33), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT32), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  AOI221_X4 g185(.A(new_n384), .B1(KEYINPUT33), .B2(new_n381), .C1(new_n369), .C2(new_n375), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n378), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n387), .ZN(new_n389));
  INV_X1    g188(.A(new_n378), .ZN(new_n390));
  INV_X1    g189(.A(new_n368), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n367), .B1(new_n235), .B2(new_n262), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n375), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT32), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n394), .B(new_n381), .C1(KEYINPUT33), .C2(new_n382), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n389), .A2(new_n390), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n388), .A2(new_n396), .A3(KEYINPUT72), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT72), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n398), .B(new_n378), .C1(new_n386), .C2(new_n387), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT89), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT4), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n367), .A2(new_n402), .A3(new_n308), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT83), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n320), .A2(new_n365), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n406), .A2(KEYINPUT83), .A3(new_n402), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT4), .B1(new_n320), .B2(new_n365), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n405), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n357), .A2(new_n364), .A3(KEYINPUT79), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT79), .B1(new_n357), .B2(new_n364), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n321), .B(new_n317), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G225gat), .A2(G233gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n414), .A2(KEYINPUT5), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n409), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n403), .A2(new_n408), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n417), .A2(new_n412), .A3(new_n413), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT79), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n365), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n357), .A2(new_n364), .A3(KEYINPUT79), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n308), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n414), .B1(new_n422), .B2(new_n406), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n418), .A2(KEYINPUT5), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT80), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT5), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n320), .B1(new_n410), .B2(new_n411), .ZN(new_n428));
  INV_X1    g227(.A(new_n406), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n427), .B1(new_n430), .B2(new_n414), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n431), .A2(KEYINPUT80), .A3(new_n418), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n416), .B1(new_n426), .B2(new_n432), .ZN(new_n433));
  XOR2_X1   g232(.A(G1gat), .B(G29gat), .Z(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(KEYINPUT82), .ZN(new_n435));
  XNOR2_X1  g234(.A(G57gat), .B(G85gat), .ZN(new_n436));
  XOR2_X1   g235(.A(new_n435), .B(new_n436), .Z(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n401), .B1(new_n433), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n409), .A2(new_n412), .A3(new_n415), .ZN(new_n441));
  AND4_X1   g240(.A1(KEYINPUT80), .A2(new_n418), .A3(KEYINPUT5), .A4(new_n423), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT80), .B1(new_n431), .B2(new_n418), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n439), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(KEYINPUT89), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n440), .A2(new_n446), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n439), .B(new_n441), .C1(new_n442), .C2(new_n443), .ZN(new_n448));
  XOR2_X1   g247(.A(KEYINPUT84), .B(KEYINPUT6), .Z(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n426), .A2(new_n432), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n439), .B1(new_n454), .B2(new_n441), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n449), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n348), .A2(new_n400), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT85), .B1(new_n451), .B2(new_n455), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n445), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT85), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n460), .A2(new_n461), .A3(new_n450), .A4(new_n448), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n459), .A2(new_n456), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n284), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n285), .A2(KEYINPUT30), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n347), .A2(new_n342), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n388), .A2(new_n396), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n468), .A2(KEYINPUT35), .A3(new_n341), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n202), .A2(new_n458), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n460), .A2(new_n450), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n471), .B1(new_n447), .B2(new_n452), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT37), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n343), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n276), .A2(KEYINPUT37), .A3(new_n277), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(new_n283), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n285), .B1(new_n476), .B2(KEYINPUT38), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT38), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT90), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n268), .A2(new_n274), .A3(new_n479), .ZN(new_n480));
  OAI211_X1 g279(.A(KEYINPUT90), .B(new_n218), .C1(new_n265), .C2(new_n267), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(KEYINPUT37), .A3(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n474), .A2(new_n478), .A3(new_n283), .A4(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n472), .A2(new_n477), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n409), .A2(new_n412), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n414), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n486), .B(KEYINPUT39), .C1(new_n414), .C2(new_n430), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n487), .B(new_n439), .C1(KEYINPUT39), .C2(new_n486), .ZN(new_n488));
  NOR2_X1   g287(.A1(KEYINPUT88), .A2(KEYINPUT40), .ZN(new_n489));
  OR2_X1    g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n489), .A2(new_n488), .B1(new_n440), .B2(new_n446), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n466), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n484), .A2(new_n492), .A3(new_n341), .ZN(new_n493));
  XNOR2_X1  g292(.A(KEYINPUT71), .B(KEYINPUT36), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n397), .A2(new_n399), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n468), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT36), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n338), .A2(new_n340), .A3(KEYINPUT87), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT87), .B1(new_n338), .B2(new_n340), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(new_n463), .B2(new_n466), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n493), .A2(new_n498), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n470), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n505));
  XNOR2_X1  g304(.A(G183gat), .B(G211gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  XOR2_X1   g307(.A(G15gat), .B(G22gat), .Z(new_n509));
  INV_X1    g308(.A(G1gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT95), .ZN(new_n512));
  AOI21_X1  g311(.A(G8gat), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n510), .A2(KEYINPUT16), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n511), .B1(new_n514), .B2(new_n509), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n513), .B(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT21), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT99), .ZN(new_n518));
  INV_X1    g317(.A(G57gat), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n518), .B1(new_n519), .B2(G64gat), .ZN(new_n520));
  INV_X1    g319(.A(G64gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n521), .A2(KEYINPUT99), .A3(G57gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n519), .A2(G64gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT100), .ZN(new_n526));
  XOR2_X1   g325(.A(G71gat), .B(G78gat), .Z(new_n527));
  AOI21_X1  g326(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n528));
  OR2_X1    g327(.A1(new_n528), .A2(KEYINPUT101), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(KEYINPUT101), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT100), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n523), .A2(new_n532), .A3(new_n524), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n526), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT9), .ZN(new_n535));
  XNOR2_X1  g334(.A(G57gat), .B(G64gat), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n527), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n516), .B1(new_n517), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT102), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G231gat), .A2(G233gat), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n542), .B(KEYINPUT103), .Z(new_n543));
  OR2_X1    g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n541), .A2(new_n543), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n538), .A2(new_n517), .ZN(new_n546));
  XOR2_X1   g345(.A(G127gat), .B(G155gat), .Z(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n544), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n548), .B1(new_n544), .B2(new_n545), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n508), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n551), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n553), .A2(new_n507), .A3(new_n549), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(G29gat), .A2(G36gat), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT14), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G29gat), .A2(G36gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT93), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(G43gat), .B(G50gat), .Z(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT92), .ZN(new_n564));
  XNOR2_X1  g363(.A(G43gat), .B(G50gat), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT92), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n564), .A2(KEYINPUT15), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT94), .B1(new_n562), .B2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n565), .B(KEYINPUT92), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT94), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n570), .A2(new_n571), .A3(KEYINPUT15), .A4(new_n561), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT17), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n562), .B(new_n568), .C1(KEYINPUT15), .C2(new_n565), .ZN(new_n575));
  AND3_X1   g374(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n574), .B1(new_n573), .B2(new_n575), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n516), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n573), .A2(new_n575), .ZN(new_n580));
  INV_X1    g379(.A(new_n516), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n578), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT96), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n584), .A2(KEYINPUT18), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT98), .B1(new_n580), .B2(new_n581), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n587), .B1(new_n581), .B2(new_n580), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n579), .B(KEYINPUT97), .Z(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT13), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n516), .A2(new_n573), .A3(KEYINPUT98), .A4(new_n575), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n585), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n578), .A2(new_n579), .A3(new_n582), .A4(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n586), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT11), .B(G169gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(G197gat), .ZN(new_n597));
  XOR2_X1   g396(.A(G113gat), .B(G141gat), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n599), .B(KEYINPUT91), .Z(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT12), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n595), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n586), .A2(new_n601), .A3(new_n592), .A4(new_n594), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT8), .ZN(new_n607));
  NAND2_X1  g406(.A1(G85gat), .A2(G92gat), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT7), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(G85gat), .ZN(new_n611));
  INV_X1    g410(.A(G92gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n607), .A2(new_n610), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G99gat), .B(G106gat), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  AOI22_X1  g417(.A1(KEYINPUT8), .A2(new_n606), .B1(new_n611), .B2(new_n612), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n619), .A2(new_n616), .A3(new_n610), .A4(new_n614), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n538), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT10), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n534), .A2(new_n621), .A3(new_n537), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n534), .A2(new_n621), .A3(new_n537), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT10), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G230gat), .A2(G233gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n630), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n621), .B1(new_n534), .B2(new_n537), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n632), .B1(new_n627), .B2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G120gat), .B(G148gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(new_n243), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(new_n204), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n631), .A2(new_n634), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n625), .A2(new_n624), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n627), .A2(new_n633), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n641), .B1(new_n642), .B2(new_n624), .ZN(new_n643));
  OAI21_X1  g442(.A(KEYINPUT104), .B1(new_n643), .B2(new_n632), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n632), .B1(new_n626), .B2(new_n628), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT104), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n644), .A2(new_n634), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n640), .B1(new_n648), .B2(new_n637), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n605), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g449(.A1(G232gat), .A2(G233gat), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n651), .A2(KEYINPUT41), .ZN(new_n652));
  XNOR2_X1  g451(.A(G190gat), .B(G218gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n622), .B1(new_n576), .B2(new_n577), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n651), .A2(KEYINPUT41), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n580), .A2(new_n621), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G134gat), .B(G162gat), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n659), .A2(new_n660), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n655), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n659), .A2(new_n660), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n665), .A2(new_n654), .A3(new_n661), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n555), .A2(new_n650), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n504), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n463), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(new_n510), .ZN(G1324gat));
  INV_X1    g471(.A(new_n669), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT16), .B(G8gat), .Z(new_n674));
  NAND3_X1  g473(.A1(new_n673), .A2(new_n466), .A3(new_n674), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n675), .A2(KEYINPUT42), .ZN(new_n676));
  INV_X1    g475(.A(new_n466), .ZN(new_n677));
  OAI21_X1  g476(.A(G8gat), .B1(new_n669), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n675), .A2(KEYINPUT42), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n676), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n680), .B1(new_n676), .B2(new_n679), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(G1325gat));
  INV_X1    g482(.A(new_n498), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n673), .A2(G15gat), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n400), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n669), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(G15gat), .B2(new_n687), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT106), .Z(G1326gat));
  INV_X1    g488(.A(new_n501), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n669), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT43), .B(G22gat), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  AND3_X1   g492(.A1(new_n493), .A2(new_n498), .A3(new_n502), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n458), .A2(new_n202), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n467), .A2(new_n469), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OAI211_X1 g496(.A(KEYINPUT107), .B(new_n667), .C1(new_n694), .C2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n667), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n701), .B1(new_n470), .B2(new_n503), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n702), .A2(KEYINPUT107), .A3(KEYINPUT44), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n555), .A2(new_n649), .A3(new_n605), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n700), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G29gat), .B1(new_n706), .B2(new_n670), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n702), .A2(new_n705), .ZN(new_n708));
  OR3_X1    g507(.A1(new_n708), .A2(G29gat), .A3(new_n670), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n709), .A2(KEYINPUT45), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n709), .A2(KEYINPUT45), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n707), .B1(new_n710), .B2(new_n711), .ZN(G1328gat));
  OAI21_X1  g511(.A(G36gat), .B1(new_n706), .B2(new_n677), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n504), .A2(new_n281), .A3(new_n667), .A4(new_n705), .ZN(new_n714));
  OAI21_X1  g513(.A(KEYINPUT46), .B1(new_n714), .B2(new_n677), .ZN(new_n715));
  AOI211_X1 g514(.A(new_n701), .B(new_n704), .C1(new_n470), .C2(new_n503), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT46), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n716), .A2(new_n717), .A3(new_n281), .A4(new_n466), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n713), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n713), .A2(new_n719), .A3(KEYINPUT108), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(G1329gat));
  OAI21_X1  g523(.A(G43gat), .B1(new_n706), .B2(new_n498), .ZN(new_n725));
  OR3_X1    g524(.A1(new_n708), .A2(G43gat), .A3(new_n686), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT47), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n725), .B(new_n726), .C1(new_n728), .C2(KEYINPUT47), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(G1330gat));
  OAI21_X1  g531(.A(G50gat), .B1(new_n706), .B2(new_n341), .ZN(new_n733));
  OR3_X1    g532(.A1(new_n708), .A2(G50gat), .A3(new_n690), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n733), .A2(KEYINPUT48), .A3(new_n734), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n700), .A2(new_n501), .A3(new_n703), .A4(new_n705), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G50gat), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n737), .A2(new_n734), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n735), .B1(new_n738), .B2(KEYINPUT48), .ZN(G1331gat));
  AOI21_X1  g538(.A(new_n649), .B1(new_n470), .B2(new_n503), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n555), .A2(new_n667), .A3(new_n605), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n670), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(new_n519), .ZN(G1332gat));
  XNOR2_X1  g543(.A(new_n466), .B(KEYINPUT110), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  AND2_X1   g547(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(new_n747), .B2(new_n748), .ZN(G1333gat));
  INV_X1    g550(.A(new_n742), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n752), .A2(G71gat), .A3(new_n684), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n742), .A2(new_n686), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n753), .B1(G71gat), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g555(.A1(new_n752), .A2(new_n501), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G78gat), .ZN(G1335gat));
  INV_X1    g557(.A(new_n555), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n605), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n504), .A2(new_n667), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT51), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n702), .A2(new_n763), .A3(new_n760), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT111), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n762), .A2(KEYINPUT111), .A3(new_n764), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n649), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n769), .A2(new_n611), .A3(new_n463), .A4(new_n770), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n759), .A2(new_n649), .A3(new_n605), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n700), .A2(new_n703), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(G85gat), .B1(new_n773), .B2(new_n670), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n771), .A2(new_n774), .ZN(G1336gat));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n776), .B1(new_n702), .B2(new_n760), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n777), .B1(new_n762), .B2(new_n764), .ZN(new_n778));
  AOI211_X1 g577(.A(new_n776), .B(KEYINPUT51), .C1(new_n702), .C2(new_n760), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n745), .A2(new_n612), .A3(new_n770), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n700), .A2(new_n466), .A3(new_n703), .A4(new_n772), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n782), .A2(G92gat), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT52), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(G92gat), .B1(new_n773), .B2(new_n746), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n785), .B(new_n786), .C1(new_n765), .C2(new_n780), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n784), .A2(new_n787), .ZN(G1337gat));
  NOR3_X1   g587(.A1(new_n686), .A2(G99gat), .A3(new_n649), .ZN(new_n789));
  XOR2_X1   g588(.A(new_n789), .B(KEYINPUT113), .Z(new_n790));
  NAND2_X1  g589(.A1(new_n769), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(G99gat), .B1(new_n773), .B2(new_n498), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(G1338gat));
  OR3_X1    g592(.A1(new_n341), .A2(new_n649), .A3(G106gat), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n778), .A2(new_n779), .A3(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n700), .A2(new_n501), .A3(new_n703), .A4(new_n772), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n796), .A2(G106gat), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT53), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(G106gat), .B1(new_n773), .B2(new_n341), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n799), .B(new_n800), .C1(new_n765), .C2(new_n794), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n801), .ZN(G1339gat));
  NAND2_X1  g601(.A1(new_n746), .A2(new_n463), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT54), .B1(new_n644), .B2(new_n647), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n626), .A2(new_n632), .A3(new_n628), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT54), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n637), .B1(new_n808), .B2(new_n645), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n805), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n804), .B1(new_n810), .B2(new_n640), .ZN(new_n811));
  INV_X1    g610(.A(new_n809), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n645), .A2(new_n646), .ZN(new_n814));
  AOI211_X1 g613(.A(KEYINPUT104), .B(new_n632), .C1(new_n626), .C2(new_n628), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n812), .A2(KEYINPUT55), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(KEYINPUT114), .A3(new_n639), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT55), .B1(new_n812), .B2(new_n816), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n811), .A2(new_n605), .A3(new_n818), .A4(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n590), .B1(new_n588), .B2(new_n591), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n579), .B1(new_n578), .B2(new_n582), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n599), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n604), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n770), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n667), .B1(new_n821), .B2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n811), .A2(new_n667), .A3(new_n818), .A4(new_n820), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n829), .A2(new_n825), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n555), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  NOR4_X1   g630(.A1(new_n555), .A2(new_n667), .A3(new_n770), .A4(new_n605), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n803), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n341), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n496), .A2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n837), .A2(new_n360), .A3(new_n605), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n834), .A2(new_n400), .A3(new_n690), .ZN(new_n839));
  INV_X1    g638(.A(new_n605), .ZN(new_n840));
  OAI21_X1  g639(.A(G113gat), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n838), .A2(new_n841), .ZN(G1340gat));
  OAI21_X1  g641(.A(G120gat), .B1(new_n839), .B2(new_n649), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n649), .A2(G120gat), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(KEYINPUT115), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n837), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n843), .A2(new_n846), .ZN(G1341gat));
  AOI21_X1  g646(.A(G127gat), .B1(new_n837), .B2(new_n759), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n839), .A2(new_n351), .A3(new_n555), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(G1342gat));
  AOI21_X1  g649(.A(new_n670), .B1(new_n831), .B2(new_n833), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n701), .A2(new_n466), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n851), .A2(new_n349), .A3(new_n836), .A4(new_n852), .ZN(new_n853));
  XOR2_X1   g652(.A(new_n853), .B(KEYINPUT56), .Z(new_n854));
  OR2_X1    g653(.A1(new_n839), .A2(new_n701), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n855), .A2(new_n856), .A3(G134gat), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n855), .B2(G134gat), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n854), .B1(new_n857), .B2(new_n858), .ZN(G1343gat));
  AOI21_X1  g658(.A(new_n341), .B1(new_n831), .B2(new_n833), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n819), .B1(new_n603), .B2(new_n604), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n817), .A2(new_n639), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  AOI22_X1  g664(.A1(new_n863), .A2(new_n865), .B1(new_n826), .B2(new_n770), .ZN(new_n866));
  OAI22_X1  g665(.A1(new_n866), .A2(new_n667), .B1(new_n829), .B2(new_n825), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n832), .B1(new_n867), .B2(new_n555), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT57), .B1(new_n868), .B2(new_n690), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n803), .A2(new_n684), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n862), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(G141gat), .B1(new_n871), .B2(new_n840), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n498), .A2(new_n835), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n873), .A2(KEYINPUT117), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(KEYINPUT117), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n851), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(new_n745), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n300), .A3(new_n605), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n872), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(KEYINPUT58), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT58), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n872), .A2(new_n878), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(G1344gat));
  NOR2_X1   g682(.A1(new_n690), .A2(KEYINPUT57), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n829), .A2(KEYINPUT119), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n819), .B1(new_n864), .B2(new_n804), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n886), .A2(new_n887), .A3(new_n667), .A4(new_n818), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n885), .A2(new_n826), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n863), .A2(new_n865), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n827), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n701), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n759), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n884), .B1(new_n893), .B2(new_n832), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n894), .B1(new_n861), .B2(new_n860), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n870), .A2(new_n770), .ZN(new_n896));
  OAI21_X1  g695(.A(G148gat), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT59), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n862), .A2(new_n869), .A3(new_n770), .A4(new_n870), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n290), .A2(KEYINPUT59), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n899), .A2(KEYINPUT118), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT118), .B1(new_n899), .B2(new_n900), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n898), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n877), .A2(new_n290), .A3(new_n770), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1345gat));
  AOI21_X1  g704(.A(G155gat), .B1(new_n877), .B2(new_n759), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n871), .A2(new_n304), .A3(new_n555), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(G1346gat));
  OAI21_X1  g707(.A(G162gat), .B1(new_n871), .B2(new_n701), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n852), .A2(new_n305), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n876), .B2(new_n910), .ZN(G1347gat));
  NAND2_X1  g710(.A1(new_n670), .A2(new_n466), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n912), .A2(new_n686), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n913), .A2(KEYINPUT120), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n914), .A2(new_n501), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n831), .A2(new_n833), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n913), .A2(KEYINPUT120), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(G169gat), .B1(new_n918), .B2(new_n840), .ZN(new_n919));
  AOI211_X1 g718(.A(new_n463), .B(new_n746), .C1(new_n831), .C2(new_n833), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n836), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n840), .A2(new_n242), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n919), .B1(new_n921), .B2(new_n922), .ZN(G1348gat));
  NOR3_X1   g722(.A1(new_n918), .A2(new_n243), .A3(new_n649), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n920), .A2(new_n836), .A3(new_n770), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n243), .B2(new_n925), .ZN(G1349gat));
  NAND4_X1  g725(.A1(new_n915), .A2(new_n759), .A3(new_n916), .A4(new_n917), .ZN(new_n927));
  AOI22_X1  g726(.A1(new_n927), .A2(G183gat), .B1(KEYINPUT122), .B2(KEYINPUT60), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n920), .A2(new_n255), .A3(new_n836), .A4(new_n759), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT122), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT60), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n932), .B2(KEYINPUT121), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n930), .B(new_n933), .ZN(G1350gat));
  OR2_X1    g733(.A1(new_n918), .A2(new_n701), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n935), .A2(new_n936), .A3(G190gat), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n936), .B1(new_n935), .B2(G190gat), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n667), .A2(new_n251), .ZN(new_n939));
  OAI22_X1  g738(.A1(new_n937), .A2(new_n938), .B1(new_n921), .B2(new_n939), .ZN(G1351gat));
  NOR2_X1   g739(.A1(new_n684), .A2(new_n912), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n894), .B(new_n941), .C1(new_n861), .C2(new_n860), .ZN(new_n942));
  OAI21_X1  g741(.A(G197gat), .B1(new_n942), .B2(new_n840), .ZN(new_n943));
  INV_X1    g742(.A(new_n873), .ZN(new_n944));
  AND4_X1   g743(.A1(new_n670), .A2(new_n916), .A3(new_n745), .A4(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(new_n203), .A3(new_n605), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT123), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT123), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n943), .A2(new_n949), .A3(new_n946), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(G1352gat));
  OR3_X1    g750(.A1(new_n942), .A2(KEYINPUT124), .A3(new_n649), .ZN(new_n952));
  OAI21_X1  g751(.A(KEYINPUT124), .B1(new_n942), .B2(new_n649), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n952), .A2(G204gat), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n945), .A2(new_n204), .A3(new_n770), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT62), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n955), .B(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n954), .A2(new_n957), .ZN(G1353gat));
  INV_X1    g757(.A(G211gat), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n945), .A2(new_n959), .A3(new_n759), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT125), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT63), .ZN(new_n962));
  OAI211_X1 g761(.A(new_n962), .B(G211gat), .C1(new_n942), .C2(new_n555), .ZN(new_n963));
  OAI21_X1  g762(.A(G211gat), .B1(new_n942), .B2(new_n555), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(KEYINPUT63), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n961), .A2(new_n963), .A3(new_n965), .ZN(G1354gat));
  AOI21_X1  g765(.A(G218gat), .B1(new_n945), .B2(new_n667), .ZN(new_n967));
  INV_X1    g766(.A(new_n942), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n667), .A2(G218gat), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(KEYINPUT126), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n967), .B1(new_n968), .B2(new_n970), .ZN(G1355gat));
endmodule


