//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 0 0 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  XNOR2_X1  g0008(.A(KEYINPUT65), .B(G68), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G107), .A2(G264), .ZN(new_n215));
  NAND4_X1  g0015(.A1(new_n212), .A2(new_n213), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n205), .B1(new_n211), .B2(new_n216), .ZN(new_n217));
  NOR2_X1   g0017(.A1(G58), .A2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT64), .Z(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n208), .B1(KEYINPUT1), .B2(new_n217), .C1(new_n221), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n217), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT67), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G226), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n231), .B(new_n232), .Z(new_n233));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT68), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n233), .B(new_n237), .Z(G358));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT69), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G41), .ZN(new_n248));
  OAI211_X1 g0048(.A(G1), .B(G13), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G33), .ZN(new_n252));
  AND2_X1   g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(G222), .A3(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n253), .A2(G223), .A3(G1698), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n255), .B(new_n256), .C1(new_n202), .C2(new_n253), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n249), .B1(new_n257), .B2(KEYINPUT71), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(KEYINPUT71), .B2(new_n257), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n261));
  INV_X1    g0061(.A(G274), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n249), .A2(new_n261), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT70), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT70), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n249), .A2(new_n266), .A3(new_n261), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n263), .B1(new_n268), .B2(G226), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n259), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(G179), .ZN(new_n271));
  NAND3_X1  g0071(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n222), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT8), .ZN(new_n274));
  INV_X1    g0074(.A(G58), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n274), .B1(new_n275), .B2(KEYINPUT72), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT72), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(KEYINPUT8), .A3(G58), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n223), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G150), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G20), .A2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  OAI22_X1  g0084(.A1(new_n282), .A2(new_n284), .B1(new_n201), .B2(new_n223), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n273), .B1(new_n281), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT73), .ZN(new_n287));
  INV_X1    g0087(.A(G13), .ZN(new_n288));
  NOR3_X1   g0088(.A1(new_n288), .A2(new_n223), .A3(G1), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(new_n273), .ZN(new_n290));
  INV_X1    g0090(.A(G50), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n291), .B1(new_n260), .B2(G20), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n290), .A2(new_n292), .B1(new_n291), .B2(new_n289), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n287), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n286), .A2(KEYINPUT73), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(G169), .B1(new_n259), .B2(new_n269), .ZN(new_n297));
  NOR3_X1   g0097(.A1(new_n271), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(KEYINPUT9), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT9), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(new_n294), .B2(new_n295), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n270), .A2(G200), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n259), .A2(G190), .A3(new_n269), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT10), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT10), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n302), .A2(new_n303), .A3(new_n307), .A4(new_n304), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n298), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n273), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n288), .A2(G1), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G20), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n310), .A2(new_n312), .A3(KEYINPUT78), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT78), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n314), .B1(new_n289), .B2(new_n273), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n260), .A2(G20), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(G68), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n209), .A2(G20), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT12), .ZN(new_n320));
  INV_X1    g0120(.A(new_n311), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G68), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT12), .B1(new_n289), .B2(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n280), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n326), .A2(G77), .B1(new_n283), .B2(G50), .ZN(new_n327));
  AOI211_X1 g0127(.A(KEYINPUT11), .B(new_n310), .C1(new_n327), .C2(new_n319), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT11), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n319), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n329), .B1(new_n330), .B2(new_n273), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n318), .B(new_n325), .C1(new_n328), .C2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n267), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n266), .B1(new_n249), .B2(new_n261), .ZN(new_n335));
  OAI21_X1  g0135(.A(G238), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G232), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G1698), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(G226), .B2(G1698), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n250), .A2(new_n252), .ZN(new_n340));
  INV_X1    g0140(.A(G97), .ZN(new_n341));
  OAI22_X1  g0141(.A1(new_n339), .A2(new_n340), .B1(new_n247), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n263), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n336), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT13), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT13), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n336), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n346), .A2(G190), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n333), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G200), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n351), .B1(new_n346), .B2(new_n348), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n348), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n347), .B1(new_n336), .B2(new_n344), .ZN(new_n355));
  OAI21_X1  g0155(.A(G169), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT14), .ZN(new_n357));
  INV_X1    g0157(.A(G169), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n358), .B1(new_n346), .B2(new_n348), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT14), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n346), .A2(G179), .A3(new_n348), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n357), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n353), .B1(new_n363), .B2(new_n332), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n316), .A2(G77), .A3(new_n317), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n365), .B(KEYINPUT79), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT76), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n283), .B(new_n367), .ZN(new_n368));
  XNOR2_X1  g0168(.A(KEYINPUT8), .B(G58), .ZN(new_n369));
  OAI22_X1  g0169(.A1(new_n368), .A2(new_n369), .B1(new_n223), .B2(new_n202), .ZN(new_n370));
  XNOR2_X1  g0170(.A(KEYINPUT15), .B(G87), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n370), .A2(KEYINPUT77), .B1(new_n326), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT77), .ZN(new_n374));
  OAI221_X1 g0174(.A(new_n374), .B1(new_n223), .B2(new_n202), .C1(new_n368), .C2(new_n369), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n376), .A2(new_n273), .B1(new_n202), .B2(new_n289), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n366), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n340), .A2(G107), .ZN(new_n379));
  MUX2_X1   g0179(.A(new_n337), .B(new_n210), .S(G1698), .Z(new_n380));
  OAI21_X1  g0180(.A(new_n379), .B1(new_n340), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n249), .B1(new_n381), .B2(KEYINPUT74), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(KEYINPUT74), .B2(new_n381), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n263), .B1(new_n268), .B2(G244), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT75), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n383), .A2(KEYINPUT75), .A3(new_n384), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n378), .B1(new_n388), .B2(G190), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n386), .A2(G200), .A3(new_n387), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(G179), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n386), .A2(new_n358), .A3(new_n387), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n393), .A2(new_n378), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n309), .A2(new_n364), .A3(new_n391), .A4(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n279), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n317), .ZN(new_n399));
  OAI22_X1  g0199(.A1(new_n399), .A2(new_n273), .B1(new_n312), .B2(new_n398), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n263), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n264), .B2(new_n337), .ZN(new_n403));
  XNOR2_X1  g0203(.A(new_n403), .B(KEYINPUT85), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G87), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n405), .B(KEYINPUT84), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT80), .B1(new_n251), .B2(G33), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT80), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n408), .A2(new_n247), .A3(KEYINPUT3), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n407), .A2(new_n409), .A3(new_n252), .ZN(new_n410));
  OR2_X1    g0210(.A1(G223), .A2(G1698), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(G226), .B2(new_n254), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n406), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n343), .ZN(new_n414));
  INV_X1    g0214(.A(G190), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n403), .B1(new_n343), .B2(new_n413), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n404), .A2(new_n416), .B1(new_n417), .B2(G200), .ZN(new_n418));
  INV_X1    g0218(.A(new_n209), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT7), .B1(new_n340), .B2(new_n223), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT7), .ZN(new_n421));
  AOI211_X1 g0221(.A(new_n421), .B(G20), .C1(new_n250), .C2(new_n252), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n419), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(G159), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n284), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n219), .B1(new_n209), .B2(new_n275), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n425), .B1(new_n426), .B2(G20), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n423), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT16), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n310), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT81), .ZN(new_n431));
  AOI21_X1  g0231(.A(G20), .B1(new_n431), .B2(new_n421), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n410), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n431), .A2(new_n421), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n410), .B(new_n432), .C1(new_n431), .C2(new_n421), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(G68), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT82), .ZN(new_n438));
  AOI211_X1 g0238(.A(new_n438), .B(new_n425), .C1(new_n426), .C2(G20), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n323), .A2(KEYINPUT65), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT65), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(G68), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n275), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(G20), .B1(new_n443), .B2(new_n218), .ZN(new_n444));
  INV_X1    g0244(.A(new_n425), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT82), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n437), .B(KEYINPUT16), .C1(new_n439), .C2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT83), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n430), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n448), .B1(new_n430), .B2(new_n447), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n401), .B(new_n418), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n451), .B(KEYINPUT17), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT18), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n430), .A2(new_n447), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT83), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n430), .A2(new_n447), .A3(new_n448), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n400), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(G179), .B1(new_n413), .B2(new_n343), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n404), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n417), .A2(G169), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n453), .B1(new_n457), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n401), .B1(new_n449), .B2(new_n450), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n465), .A2(KEYINPUT18), .A3(new_n462), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n452), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n397), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n250), .A2(new_n252), .A3(G250), .A4(G1698), .ZN(new_n471));
  AND2_X1   g0271(.A1(KEYINPUT4), .A2(G244), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n250), .A2(new_n252), .A3(new_n472), .A4(new_n254), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G283), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n471), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT4), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n407), .A2(new_n409), .A3(G244), .A4(new_n252), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n476), .B1(new_n477), .B2(G1698), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n343), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT5), .B(G41), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n260), .A2(G45), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n481), .A2(new_n249), .A3(G274), .A4(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n482), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(G257), .A3(new_n249), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n480), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n358), .ZN(new_n487));
  INV_X1    g0287(.A(G107), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n421), .B1(new_n253), .B2(G20), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n340), .A2(KEYINPUT7), .A3(new_n223), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT6), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n492), .A2(new_n341), .A3(G107), .ZN(new_n493));
  XNOR2_X1  g0293(.A(G97), .B(G107), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n493), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  OAI22_X1  g0295(.A1(new_n495), .A2(new_n223), .B1(new_n202), .B2(new_n284), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n273), .B1(new_n491), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n312), .A2(G97), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n260), .A2(G33), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n290), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n499), .B1(new_n501), .B2(new_n341), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n497), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT86), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n485), .A2(new_n483), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT87), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n485), .A2(KEYINPUT87), .A3(new_n483), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n480), .A2(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n249), .B1(new_n475), .B2(new_n478), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT86), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n487), .B(new_n504), .C1(new_n513), .C2(G179), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n351), .B1(new_n510), .B2(new_n512), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n494), .A2(new_n492), .ZN(new_n516));
  INV_X1    g0316(.A(new_n493), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n518), .A2(G20), .B1(G77), .B2(new_n283), .ZN(new_n519));
  OAI21_X1  g0319(.A(G107), .B1(new_n420), .B2(new_n422), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n502), .B1(new_n521), .B2(new_n273), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(new_n486), .B2(new_n415), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n515), .A2(new_n523), .A3(KEYINPUT88), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT88), .ZN(new_n525));
  INV_X1    g0325(.A(new_n509), .ZN(new_n526));
  AOI21_X1  g0326(.A(KEYINPUT87), .B1(new_n485), .B2(new_n483), .ZN(new_n527));
  OAI22_X1  g0327(.A1(new_n526), .A2(new_n527), .B1(new_n511), .B2(KEYINPUT86), .ZN(new_n528));
  INV_X1    g0328(.A(new_n512), .ZN(new_n529));
  OAI21_X1  g0329(.A(G200), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n511), .A2(new_n415), .A3(new_n506), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n504), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n525), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n514), .B1(new_n524), .B2(new_n533), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n407), .A2(new_n409), .A3(new_n252), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT89), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n535), .A2(new_n536), .A3(G264), .A4(G1698), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(G257), .A3(new_n254), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n340), .A2(G303), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G264), .A2(G1698), .ZN(new_n540));
  OAI21_X1  g0340(.A(KEYINPUT89), .B1(new_n410), .B2(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n537), .A2(new_n538), .A3(new_n539), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n343), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n343), .B1(new_n482), .B2(new_n481), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G270), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n483), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(G116), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G20), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n321), .A2(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n474), .B(new_n223), .C1(G33), .C2(new_n341), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n551), .A2(new_n273), .A3(new_n549), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT20), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n551), .A2(KEYINPUT20), .A3(new_n273), .A4(new_n549), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n550), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n313), .A2(new_n315), .A3(G116), .A4(new_n500), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n543), .A2(G179), .A3(new_n547), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT90), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n546), .B1(new_n542), .B2(new_n343), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT90), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n561), .A2(new_n562), .A3(G179), .A4(new_n558), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n543), .A2(new_n547), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT21), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n358), .B1(new_n556), .B2(new_n557), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n566), .ZN(new_n568));
  OAI21_X1  g0368(.A(KEYINPUT21), .B1(new_n568), .B2(new_n561), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n560), .A2(new_n563), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n561), .A2(G190), .ZN(new_n571));
  INV_X1    g0371(.A(new_n558), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n571), .B(new_n572), .C1(new_n351), .C2(new_n561), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT91), .ZN(new_n574));
  NAND2_X1  g0374(.A1(G33), .A2(G116), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n574), .B1(new_n575), .B2(G20), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n223), .A2(KEYINPUT91), .A3(G33), .A4(G116), .ZN(new_n577));
  OAI21_X1  g0377(.A(KEYINPUT23), .B1(new_n223), .B2(G107), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n250), .A2(new_n252), .A3(new_n223), .A4(G87), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT22), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(G87), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n581), .A2(new_n583), .A3(G20), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n584), .A2(new_n407), .A3(new_n409), .A4(new_n252), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT23), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n586), .A2(new_n488), .A3(G20), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(KEYINPUT92), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT92), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n589), .A2(new_n586), .A3(new_n488), .A4(G20), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n579), .A2(new_n582), .A3(new_n585), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT24), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n580), .A2(new_n581), .B1(new_n588), .B2(new_n590), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT24), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n594), .A2(new_n595), .A3(new_n585), .A4(new_n579), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n273), .ZN(new_n598));
  INV_X1    g0398(.A(G250), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n254), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(G257), .B2(new_n254), .ZN(new_n601));
  INV_X1    g0401(.A(G294), .ZN(new_n602));
  OAI22_X1  g0402(.A1(new_n410), .A2(new_n601), .B1(new_n247), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n603), .A2(new_n343), .B1(new_n544), .B2(G264), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n483), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(G200), .ZN(new_n606));
  INV_X1    g0406(.A(new_n501), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT25), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n312), .B2(G107), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n289), .A2(KEYINPUT25), .A3(new_n488), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n607), .A2(G107), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n604), .A2(G190), .A3(new_n483), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n598), .A2(new_n606), .A3(new_n611), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n605), .A2(new_n358), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n604), .A2(new_n392), .A3(new_n483), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n310), .B1(new_n593), .B2(new_n596), .ZN(new_n616));
  INV_X1    g0416(.A(new_n611), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n614), .B(new_n615), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT19), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n223), .B1(new_n247), .B2(new_n341), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n583), .A2(new_n341), .A3(new_n488), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NOR3_X1   g0423(.A1(new_n280), .A2(KEYINPUT19), .A3(new_n341), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n223), .A2(G68), .ZN(new_n625));
  OAI22_X1  g0425(.A1(new_n623), .A2(new_n624), .B1(new_n410), .B2(new_n625), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n626), .A2(new_n273), .B1(new_n289), .B2(new_n371), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n607), .A2(G87), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n407), .A2(new_n409), .A3(new_n254), .A4(new_n252), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n575), .B1(new_n630), .B2(new_n210), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n477), .A2(new_n254), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n343), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n343), .A2(new_n599), .A3(new_n482), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n634), .B1(G274), .B2(new_n482), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n629), .B1(G200), .B2(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n633), .A2(new_n635), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(G190), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n607), .A2(new_n372), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n636), .A2(new_n358), .B1(new_n627), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n638), .A2(new_n392), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n637), .A2(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n570), .A2(new_n573), .A3(new_n619), .A4(new_n643), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n470), .A2(new_n534), .A3(new_n644), .ZN(G372));
  INV_X1    g0445(.A(KEYINPUT93), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n465), .A2(KEYINPUT18), .A3(new_n462), .ZN(new_n647));
  AOI21_X1  g0447(.A(KEYINPUT18), .B1(new_n465), .B2(new_n462), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n464), .A2(KEYINPUT93), .A3(new_n466), .ZN(new_n650));
  INV_X1    g0450(.A(new_n353), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n395), .A2(new_n651), .B1(new_n332), .B2(new_n363), .ZN(new_n652));
  INV_X1    g0452(.A(new_n452), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n649), .B(new_n650), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n306), .A2(new_n308), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n298), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n636), .A2(G200), .ZN(new_n658));
  INV_X1    g0458(.A(new_n629), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n639), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n641), .A2(new_n642), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n657), .B1(new_n514), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n511), .A2(new_n506), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n504), .B1(G169), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n528), .A2(new_n529), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n665), .B1(new_n392), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n667), .A2(KEYINPUT26), .A3(new_n643), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n660), .A2(new_n613), .A3(new_n661), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n560), .A2(new_n563), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n567), .A2(new_n569), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n618), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n670), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n669), .B(new_n661), .C1(new_n534), .C2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n656), .B1(new_n470), .B2(new_n677), .ZN(G369));
  INV_X1    g0478(.A(KEYINPUT95), .ZN(new_n679));
  OR3_X1    g0479(.A1(new_n321), .A2(KEYINPUT27), .A3(G20), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT27), .B1(new_n321), .B2(G20), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G213), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G343), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n679), .B1(new_n618), .B2(new_n685), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n614), .A2(new_n615), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n598), .A2(new_n611), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n687), .A2(new_n688), .A3(KEYINPUT95), .A4(new_n684), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n684), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n691), .A2(new_n618), .A3(new_n613), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n558), .A2(new_n684), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n671), .A2(new_n672), .A3(new_n573), .A4(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n570), .B2(new_n694), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT94), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n696), .A2(new_n697), .A3(G330), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n697), .B1(new_n696), .B2(G330), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n693), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n618), .A2(new_n684), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n570), .A2(new_n684), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n701), .B1(new_n693), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n700), .A2(new_n703), .ZN(G399));
  INV_X1    g0504(.A(new_n206), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n622), .A2(G116), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(G1), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n220), .B2(new_n707), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n513), .A2(new_n605), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n564), .A2(new_n392), .A3(new_n636), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT97), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT97), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n564), .A2(new_n715), .A3(new_n392), .A4(new_n636), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n712), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n561), .A2(G179), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n664), .A2(new_n604), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n719), .A2(new_n720), .A3(KEYINPUT30), .A4(new_n638), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n638), .A2(new_n664), .A3(new_n604), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(new_n718), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n684), .B1(new_n717), .B2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT31), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XOR2_X1   g0528(.A(KEYINPUT96), .B(KEYINPUT31), .Z(new_n729));
  OAI21_X1  g0529(.A(new_n728), .B1(new_n726), .B2(new_n729), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n644), .A2(new_n534), .A3(new_n684), .ZN(new_n731));
  OAI21_X1  g0531(.A(G330), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n676), .A2(new_n685), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(KEYINPUT29), .ZN(new_n734));
  OAI21_X1  g0534(.A(KEYINPUT88), .B1(new_n515), .B2(new_n523), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n530), .A2(new_n525), .A3(new_n532), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n667), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n737), .B(new_n670), .C1(new_n673), .C2(new_n674), .ZN(new_n738));
  AOI22_X1  g0538(.A1(new_n663), .A2(new_n668), .B1(new_n642), .B2(new_n641), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n684), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT29), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n732), .A2(new_n734), .A3(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n711), .B1(new_n744), .B2(G1), .ZN(G364));
  NAND2_X1  g0545(.A1(new_n696), .A2(G330), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(KEYINPUT94), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n696), .A2(new_n697), .A3(G330), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n288), .A2(G20), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n260), .B1(new_n751), .B2(G45), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n706), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n750), .B(new_n755), .C1(G330), .C2(new_n696), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n223), .A2(G190), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n392), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G179), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n424), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT32), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n253), .B1(new_n202), .B2(new_n759), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n351), .A2(G179), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n757), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n488), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n223), .A2(new_n415), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n765), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n767), .B1(G87), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n392), .A2(new_n351), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n768), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n768), .A2(new_n758), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n771), .B1(new_n291), .B2(new_n773), .C1(new_n275), .C2(new_n774), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n764), .B(new_n775), .C1(new_n763), .C2(new_n762), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n760), .A2(G190), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G20), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G97), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT100), .ZN(new_n780));
  AND3_X1   g0580(.A1(new_n772), .A2(new_n780), .A3(new_n757), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n780), .B1(new_n772), .B2(new_n757), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n779), .B1(new_n784), .B2(new_n323), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT101), .Z(new_n786));
  INV_X1    g0586(.A(G303), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n340), .B1(new_n769), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT102), .ZN(new_n789));
  INV_X1    g0589(.A(new_n761), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G329), .ZN(new_n791));
  INV_X1    g0591(.A(G283), .ZN(new_n792));
  INV_X1    g0592(.A(G322), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n791), .B1(new_n792), .B2(new_n766), .C1(new_n793), .C2(new_n774), .ZN(new_n794));
  INV_X1    g0594(.A(new_n773), .ZN(new_n795));
  INV_X1    g0595(.A(new_n759), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G326), .A2(new_n795), .B1(new_n796), .B2(G311), .ZN(new_n797));
  INV_X1    g0597(.A(new_n778), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n602), .B2(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(KEYINPUT33), .B(G317), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n794), .B(new_n799), .C1(new_n783), .C2(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n776), .A2(new_n786), .B1(new_n789), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n222), .B1(G20), .B2(new_n358), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n754), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n705), .A2(new_n340), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n806), .A2(G355), .B1(new_n548), .B2(new_n705), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n242), .A2(G45), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT98), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n535), .A2(new_n705), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n221), .B2(G45), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n807), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(G13), .A2(G33), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(G20), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n803), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT99), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n805), .B1(new_n812), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n815), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n819), .B1(new_n696), .B2(new_n820), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n756), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(G396));
  NAND4_X1  g0623(.A1(new_n393), .A2(new_n378), .A3(new_n394), .A4(new_n685), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n389), .A2(new_n390), .B1(new_n378), .B2(new_n684), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n825), .B2(new_n395), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(new_n814), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n803), .A2(new_n813), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n774), .ZN(new_n831));
  AOI22_X1  g0631(.A1(G137), .A2(new_n795), .B1(new_n831), .B2(G143), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n832), .B1(new_n424), .B2(new_n759), .C1(new_n784), .C2(new_n282), .ZN(new_n833));
  XOR2_X1   g0633(.A(KEYINPUT104), .B(KEYINPUT34), .Z(new_n834));
  XNOR2_X1  g0634(.A(new_n833), .B(new_n834), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n769), .A2(new_n291), .B1(new_n766), .B2(new_n323), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n535), .B1(new_n798), .B2(new_n275), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n836), .B(new_n837), .C1(G132), .C2(new_n790), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n340), .B1(new_n769), .B2(new_n488), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT103), .ZN(new_n840));
  INV_X1    g0640(.A(G311), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n779), .B1(new_n787), .B2(new_n773), .C1(new_n841), .C2(new_n761), .ZN(new_n842));
  INV_X1    g0642(.A(new_n766), .ZN(new_n843));
  AOI22_X1  g0643(.A1(G87), .A2(new_n843), .B1(new_n796), .B2(G116), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n602), .B2(new_n774), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n842), .B(new_n845), .C1(G283), .C2(new_n783), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n835), .A2(new_n838), .B1(new_n840), .B2(new_n846), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n754), .B1(G77), .B2(new_n830), .C1(new_n847), .C2(new_n804), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n828), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n740), .B(new_n826), .ZN(new_n850));
  INV_X1    g0650(.A(new_n732), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n852), .A2(KEYINPUT105), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n850), .A2(new_n851), .ZN(new_n854));
  NOR3_X1   g0654(.A1(new_n853), .A2(new_n754), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n852), .A2(KEYINPUT105), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n849), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G384));
  NOR2_X1   g0658(.A1(new_n751), .A2(new_n260), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n362), .B1(new_n359), .B2(new_n360), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n356), .A2(KEYINPUT14), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n332), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n332), .A2(new_n684), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n862), .A2(new_n651), .A3(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT106), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n364), .A2(KEYINPUT106), .A3(new_n863), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n363), .A2(new_n332), .A3(new_n684), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n826), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n727), .B(new_n684), .C1(new_n717), .C2(new_n725), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n721), .A2(new_n724), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n714), .A2(new_n716), .ZN(new_n874));
  INV_X1    g0674(.A(new_n712), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n729), .B1(new_n877), .B2(new_n684), .ZN(new_n878));
  AND4_X1   g0678(.A1(new_n570), .A2(new_n573), .A3(new_n619), .A4(new_n643), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(new_n737), .A3(new_n685), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n872), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n870), .A2(KEYINPUT40), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g0682(.A(KEYINPUT108), .B(KEYINPUT38), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n649), .A2(new_n452), .A3(new_n650), .ZN(new_n885));
  INV_X1    g0685(.A(new_n682), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n465), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n646), .B1(new_n457), .B2(new_n463), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n465), .A2(KEYINPUT93), .A3(new_n462), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n890), .A2(new_n451), .A3(new_n887), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(KEYINPUT37), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT109), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n887), .A2(new_n451), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT37), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n457), .B2(new_n463), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n894), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n897), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n899), .A2(KEYINPUT109), .A3(new_n451), .A4(new_n887), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n893), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n884), .B1(new_n889), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n895), .A2(new_n897), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n439), .A2(new_n446), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT16), .B1(new_n904), .B2(new_n437), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n447), .A2(new_n273), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n401), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n462), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n451), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT107), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n907), .A2(new_n886), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n908), .A2(new_n451), .A3(KEYINPUT107), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n903), .B1(new_n914), .B2(KEYINPUT37), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT38), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n912), .B1(new_n452), .B2(new_n467), .ZN(new_n917));
  NOR3_X1   g0717(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n882), .B1(new_n902), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT110), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n870), .A2(new_n881), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n913), .A2(new_n912), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT107), .B1(new_n908), .B2(new_n451), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT37), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n895), .B2(new_n897), .ZN(new_n926));
  INV_X1    g0726(.A(new_n917), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT38), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n922), .B1(new_n928), .B2(new_n918), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT40), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n882), .B(KEYINPUT110), .C1(new_n902), .C2(new_n918), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n921), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n933), .A2(new_n469), .A3(new_n881), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(G330), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n933), .B1(new_n469), .B2(new_n881), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT39), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n902), .B2(new_n918), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n363), .A2(new_n332), .A3(new_n685), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n926), .A2(KEYINPUT38), .A3(new_n927), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n916), .B1(new_n915), .B2(new_n917), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n942), .A2(new_n943), .A3(KEYINPUT39), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n939), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n886), .B1(new_n649), .B2(new_n650), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n740), .A2(new_n827), .B1(new_n395), .B2(new_n685), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n864), .A2(new_n865), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT106), .B1(new_n364), .B2(new_n863), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n869), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n942), .A2(new_n943), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n946), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n945), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n734), .A2(new_n742), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n469), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n656), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n955), .B(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n859), .B1(new_n937), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n959), .B2(new_n937), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n548), .B(new_n225), .C1(new_n518), .C2(KEYINPUT35), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(KEYINPUT35), .B2(new_n518), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT36), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n443), .A2(new_n220), .A3(new_n202), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n323), .A2(G50), .ZN(new_n966));
  OAI211_X1 g0766(.A(G1), .B(new_n288), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n961), .A2(new_n964), .A3(new_n967), .ZN(G367));
  INV_X1    g0768(.A(new_n810), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n818), .B1(new_n206), .B2(new_n371), .C1(new_n237), .C2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n755), .B1(new_n970), .B2(KEYINPUT115), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(KEYINPUT115), .B2(new_n970), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n798), .A2(new_n323), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n769), .A2(new_n275), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(G143), .B2(new_n795), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n975), .B(new_n253), .C1(new_n282), .C2(new_n774), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n784), .A2(new_n424), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n766), .A2(new_n202), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(G50), .B2(new_n796), .ZN(new_n979));
  INV_X1    g0779(.A(G137), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n979), .B1(new_n980), .B2(new_n761), .ZN(new_n981));
  OR4_X1    g0781(.A1(new_n973), .A2(new_n976), .A3(new_n977), .A4(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n769), .A2(new_n548), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT46), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(G107), .B2(new_n778), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n783), .A2(G294), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n766), .A2(new_n341), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n774), .A2(new_n787), .ZN(new_n988));
  XOR2_X1   g0788(.A(KEYINPUT116), .B(G311), .Z(new_n989));
  AOI211_X1 g0789(.A(new_n987), .B(new_n988), .C1(new_n795), .C2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(G317), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n759), .A2(new_n792), .B1(new_n761), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n992), .A2(new_n535), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n985), .A2(new_n986), .A3(new_n990), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n982), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT47), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n972), .B1(new_n996), .B2(new_n803), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n659), .A2(new_n685), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n643), .A2(KEYINPUT111), .A3(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n661), .B2(new_n999), .ZN(new_n1001));
  AOI21_X1  g0801(.A(KEYINPUT111), .B1(new_n643), .B2(new_n999), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n997), .B1(new_n1004), .B2(new_n820), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT44), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n667), .A2(new_n684), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n522), .A2(new_n685), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1008), .B1(new_n534), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1007), .B1(new_n703), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n701), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n619), .A2(new_n691), .B1(new_n686), .B2(new_n689), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n673), .A2(new_n685), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1009), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n737), .A2(new_n1016), .B1(new_n667), .B2(new_n684), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1015), .A2(new_n1017), .A3(KEYINPUT44), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1011), .A2(new_n1018), .A3(KEYINPUT113), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT45), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n703), .A2(new_n1010), .A3(KEYINPUT45), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g0823(.A(KEYINPUT114), .B(new_n693), .C1(new_n698), .C2(new_n699), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT113), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1025), .B(new_n1007), .C1(new_n703), .C2(new_n1010), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1019), .A2(new_n1023), .A3(new_n1024), .A4(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT114), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n700), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(KEYINPUT44), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n1021), .A2(new_n1022), .B1(new_n1032), .B2(new_n1025), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1033), .A2(new_n1029), .A3(new_n1024), .A4(new_n1019), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n693), .B(new_n1014), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n749), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n749), .A2(new_n1036), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1039), .A2(new_n743), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n743), .B1(new_n1035), .B2(new_n1040), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n706), .B(KEYINPUT41), .Z(new_n1042));
  OAI21_X1  g0842(.A(new_n752), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n1010), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(KEYINPUT42), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT42), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1044), .A2(new_n1010), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n674), .B1(new_n524), .B2(new_n533), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n514), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n685), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1046), .A2(new_n1048), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT43), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1003), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(KEYINPUT43), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1052), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1045), .A2(KEYINPUT42), .B1(new_n685), .B2(new_n1050), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1057), .A2(new_n1003), .A3(new_n1053), .A4(new_n1048), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n700), .A2(new_n1017), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT112), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  AOI211_X1 g0865(.A(KEYINPUT112), .B(new_n1060), .C1(new_n1056), .C2(new_n1058), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1062), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1006), .B1(new_n1043), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(G387));
  INV_X1    g0870(.A(new_n1039), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1013), .A2(new_n815), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n708), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n806), .A2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(G107), .B2(new_n206), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n233), .A2(G45), .ZN(new_n1076));
  AOI211_X1 g0876(.A(G45), .B(new_n1073), .C1(G68), .C2(G77), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n369), .A2(G50), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT50), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n969), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1075), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n754), .B1(new_n1081), .B2(new_n817), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n410), .B(new_n987), .C1(G77), .C2(new_n770), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n783), .A2(new_n398), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n798), .A2(new_n371), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n773), .A2(new_n424), .B1(new_n759), .B2(new_n323), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n774), .A2(new_n291), .B1(new_n761), .B2(new_n282), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .A4(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n774), .A2(new_n991), .B1(new_n759), .B2(new_n787), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT117), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n783), .A2(new_n989), .B1(G322), .B2(new_n795), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n1094), .A2(KEYINPUT48), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1094), .A2(KEYINPUT48), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n798), .A2(new_n792), .B1(new_n769), .B2(new_n602), .ZN(new_n1097));
  NOR3_X1   g0897(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  XOR2_X1   g0899(.A(KEYINPUT118), .B(KEYINPUT49), .Z(new_n1100));
  NOR2_X1   g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G116), .A2(new_n843), .B1(new_n790), .B2(G326), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1100), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n410), .B(new_n1102), .C1(new_n1098), .C2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1090), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1082), .B1(new_n1105), .B2(new_n803), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1071), .A2(new_n753), .B1(new_n1072), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1039), .A2(new_n743), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n734), .A2(new_n742), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1109), .A2(new_n1037), .A3(new_n732), .A4(new_n1038), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1108), .A2(new_n1110), .A3(new_n706), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1107), .A2(new_n1111), .ZN(G393));
  NAND2_X1  g0912(.A1(new_n1017), .A2(new_n815), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n818), .B1(new_n341), .B2(new_n206), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n245), .A2(new_n810), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n754), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n369), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1117), .A2(new_n796), .B1(new_n843), .B2(G87), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n419), .A2(new_n770), .B1(new_n790), .B2(G143), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n778), .A2(G77), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1118), .A2(new_n1119), .A3(new_n535), .A4(new_n1120), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n773), .A2(new_n282), .B1(new_n774), .B2(new_n424), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT51), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n291), .B2(new_n784), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n253), .B(new_n767), .C1(G116), .C2(new_n778), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n769), .A2(new_n792), .B1(new_n761), .B2(new_n793), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(G294), .B2(new_n796), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1125), .B(new_n1127), .C1(new_n787), .C2(new_n784), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n773), .A2(new_n991), .B1(new_n774), .B2(new_n841), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(KEYINPUT119), .B(KEYINPUT52), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1129), .B(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n1121), .A2(new_n1124), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1116), .B1(new_n1132), .B2(new_n803), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1035), .A2(new_n753), .B1(new_n1113), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1035), .A2(new_n1040), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1110), .A2(new_n1031), .A3(new_n1034), .ZN(new_n1136));
  AND4_X1   g0936(.A1(KEYINPUT120), .A2(new_n1135), .A3(new_n706), .A4(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n707), .B1(new_n1035), .B2(new_n1040), .ZN(new_n1138));
  AOI21_X1  g0938(.A(KEYINPUT120), .B1(new_n1138), .B2(new_n1136), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1134), .B1(new_n1137), .B2(new_n1139), .ZN(G390));
  NAND2_X1  g0940(.A1(new_n889), .A2(new_n901), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n883), .ZN(new_n1142));
  AOI21_X1  g0942(.A(KEYINPUT39), .B1(new_n1142), .B2(new_n942), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n942), .A2(new_n943), .A3(KEYINPUT39), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n813), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(G125), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n253), .B1(new_n761), .B2(new_n1146), .C1(new_n798), .C2(new_n424), .ZN(new_n1147));
  INV_X1    g0947(.A(G128), .ZN(new_n1148));
  INV_X1    g0948(.A(G132), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n773), .A2(new_n1148), .B1(new_n774), .B2(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT54), .B(G143), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n291), .A2(new_n766), .B1(new_n759), .B2(new_n1151), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1147), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n769), .A2(new_n282), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT53), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1153), .B(new_n1155), .C1(new_n980), .C2(new_n784), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n773), .A2(new_n792), .B1(new_n766), .B2(new_n323), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n253), .B(new_n1157), .C1(G87), .C2(new_n770), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n783), .A2(G107), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n759), .A2(new_n341), .B1(new_n761), .B2(new_n602), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(G116), .B2(new_n831), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1158), .A2(new_n1120), .A3(new_n1159), .A4(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n804), .B1(new_n1156), .B2(new_n1162), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n755), .B(new_n1163), .C1(new_n279), .C2(new_n829), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1145), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n940), .B1(new_n947), .B2(new_n951), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n824), .B1(new_n733), .B2(new_n826), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n941), .B1(new_n1168), .B2(new_n950), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n918), .B2(new_n902), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n851), .A2(new_n870), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1167), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT121), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n950), .A2(new_n827), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n729), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n726), .A2(new_n1175), .ZN(new_n1176));
  OAI211_X1 g0976(.A(G330), .B(new_n871), .C1(new_n731), .C2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1173), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n870), .A2(new_n881), .A3(KEYINPUT121), .A4(G330), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1169), .B1(new_n939), .B2(new_n944), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1166), .B1(new_n942), .B2(new_n1142), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1180), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1172), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1165), .B1(new_n1184), .B2(new_n752), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n957), .B(new_n656), .C1(new_n470), .C2(new_n1177), .ZN(new_n1186));
  OAI211_X1 g0986(.A(G330), .B(new_n827), .C1(new_n730), .C2(new_n731), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n1187), .A2(new_n951), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1168), .B1(new_n1180), .B2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n951), .B1(new_n1177), .B2(new_n826), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1171), .A2(new_n947), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1186), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1172), .A2(new_n1183), .A3(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1192), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n707), .B1(new_n1184), .B2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1185), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(G378));
  NOR2_X1   g0997(.A1(new_n296), .A2(new_n682), .ZN(new_n1198));
  XOR2_X1   g0998(.A(KEYINPUT123), .B(KEYINPUT56), .Z(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  AND2_X1   g1000(.A1(new_n309), .A2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n309), .A2(new_n1200), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1198), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n309), .A2(new_n1200), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n309), .A2(new_n1200), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1198), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1203), .A2(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(KEYINPUT124), .B(KEYINPUT55), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1203), .A2(new_n1207), .A3(new_n1209), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n813), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n754), .B1(new_n830), .B2(G50), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT122), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n535), .A2(G41), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G97), .B2(new_n783), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(G107), .A2(new_n831), .B1(new_n790), .B2(G283), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G116), .A2(new_n795), .B1(new_n796), .B2(new_n372), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n769), .A2(new_n202), .B1(new_n766), .B2(new_n275), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n973), .A2(new_n1223), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .A4(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT58), .ZN(new_n1226));
  AOI21_X1  g1026(.A(G50), .B1(new_n247), .B2(new_n248), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1225), .A2(new_n1226), .B1(new_n1219), .B2(new_n1227), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n769), .A2(new_n1151), .B1(new_n759), .B2(new_n980), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n773), .A2(new_n1146), .B1(new_n774), .B2(new_n1148), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1229), .B(new_n1230), .C1(G150), .C2(new_n778), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n1149), .B2(new_n784), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n843), .A2(G159), .ZN(new_n1234));
  AOI211_X1 g1034(.A(G33), .B(G41), .C1(new_n790), .C2(G124), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n1228), .B1(new_n1226), .B2(new_n1225), .C1(new_n1236), .C2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1217), .B1(new_n1238), .B2(new_n803), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1215), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n955), .A2(new_n1214), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n945), .A2(new_n1213), .A3(new_n954), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1242), .A2(new_n933), .A3(G330), .A4(new_n1243), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n921), .A2(new_n931), .A3(G330), .A4(new_n932), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n945), .A2(new_n1213), .A3(new_n954), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1213), .B1(new_n945), .B2(new_n954), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1245), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1244), .A2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1241), .B1(new_n1249), .B2(new_n753), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1186), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1193), .A2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1249), .A2(KEYINPUT57), .A3(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n706), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1244), .A2(new_n1248), .B1(new_n1193), .B2(new_n1251), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1255), .A2(KEYINPUT57), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1250), .B1(new_n1254), .B2(new_n1256), .ZN(G375));
  AOI21_X1  g1057(.A(new_n755), .B1(new_n323), .B2(new_n829), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(G107), .A2(new_n796), .B1(new_n790), .B2(G303), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1259), .B1(new_n341), .B2(new_n769), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(G116), .B2(new_n783), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n773), .A2(new_n602), .B1(new_n774), .B2(new_n792), .ZN(new_n1262));
  NOR4_X1   g1062(.A1(new_n1085), .A2(new_n1262), .A3(new_n253), .A4(new_n978), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n769), .A2(new_n424), .B1(new_n766), .B2(new_n275), .ZN(new_n1264));
  AOI211_X1 g1064(.A(new_n410), .B(new_n1264), .C1(G50), .C2(new_n778), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n759), .A2(new_n282), .B1(new_n761), .B2(new_n1148), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n773), .A2(new_n1149), .B1(new_n774), .B2(new_n980), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1151), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n1266), .B(new_n1267), .C1(new_n783), .C2(new_n1268), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n1261), .A2(new_n1263), .B1(new_n1265), .B2(new_n1269), .ZN(new_n1270));
  OAI221_X1 g1070(.A(new_n1258), .B1(new_n804), .B2(new_n1270), .C1(new_n950), .C2(new_n814), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1272), .B1(new_n1273), .B2(new_n753), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1042), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1194), .A2(new_n1275), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1273), .A2(new_n1251), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1274), .B1(new_n1276), .B2(new_n1277), .ZN(G381));
  AOI22_X1  g1078(.A1(new_n1242), .A2(new_n1243), .B1(new_n933), .B2(G330), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1246), .A2(new_n1247), .A3(new_n1245), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n753), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1240), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n707), .B1(new_n1255), .B2(KEYINPUT57), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1249), .A2(new_n1252), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT57), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1282), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1196), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1107), .A2(new_n1111), .A3(new_n822), .ZN(new_n1289));
  OR3_X1    g1089(.A1(G381), .A2(G384), .A3(new_n1289), .ZN(new_n1290));
  OR4_X1    g1090(.A1(G387), .A2(new_n1288), .A3(G390), .A4(new_n1290), .ZN(G407));
  OAI211_X1 g1091(.A(G407), .B(G213), .C1(G343), .C2(new_n1288), .ZN(G409));
  NAND2_X1  g1092(.A1(G375), .A2(G378), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1249), .A2(new_n1275), .A3(new_n1252), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1196), .A2(new_n1250), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n683), .A2(G213), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1277), .B1(KEYINPUT60), .B2(new_n1194), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1189), .A2(new_n1186), .A3(KEYINPUT60), .A4(new_n1191), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n706), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1274), .B1(new_n1298), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n857), .ZN(new_n1302));
  OAI211_X1 g1102(.A(G384), .B(new_n1274), .C1(new_n1298), .C2(new_n1300), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1293), .A2(new_n1297), .A3(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(KEYINPUT62), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1296), .B(new_n1295), .C1(new_n1287), .C2(new_n1196), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n683), .A2(G213), .A3(G2897), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1302), .A2(new_n1303), .A3(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1309), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(KEYINPUT61), .B1(new_n1308), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT62), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1293), .A2(new_n1297), .A3(new_n1314), .A4(new_n1305), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1307), .A2(new_n1313), .A3(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT126), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1135), .A2(new_n706), .A3(new_n1136), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT120), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1138), .A2(KEYINPUT120), .A3(new_n1136), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  OAI22_X1  g1122(.A1(new_n1064), .A2(new_n1066), .B1(new_n1061), .B2(new_n1059), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1110), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1275), .B1(new_n1324), .B2(new_n743), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1323), .B1(new_n1325), .B2(new_n752), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1322), .B(new_n1134), .C1(new_n1326), .C2(new_n1006), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(G390), .A2(new_n1069), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n822), .B1(new_n1107), .B2(new_n1111), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1330), .A2(KEYINPUT125), .A3(new_n1289), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT125), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1289), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1332), .B1(new_n1333), .B2(new_n1329), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1331), .A2(new_n1334), .ZN(new_n1335));
  AND4_X1   g1135(.A1(new_n1317), .A2(new_n1327), .A3(new_n1328), .A4(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(KEYINPUT126), .B1(G390), .B2(new_n1069), .ZN(new_n1337));
  AOI22_X1  g1137(.A1(new_n1337), .A2(new_n1335), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1336), .A2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1316), .A2(new_n1339), .ZN(new_n1340));
  AOI211_X1 g1140(.A(KEYINPUT61), .B(new_n1339), .C1(new_n1308), .C2(new_n1312), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT63), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1306), .A2(new_n1342), .ZN(new_n1343));
  OAI21_X1  g1143(.A(KEYINPUT127), .B1(new_n1306), .B2(new_n1342), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1345), .B1(G378), .B2(G375), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT127), .ZN(new_n1347));
  NAND4_X1  g1147(.A1(new_n1346), .A2(new_n1347), .A3(KEYINPUT63), .A4(new_n1305), .ZN(new_n1348));
  NAND4_X1  g1148(.A1(new_n1341), .A2(new_n1343), .A3(new_n1344), .A4(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1340), .A2(new_n1349), .ZN(G405));
  NAND2_X1  g1150(.A1(new_n1293), .A2(new_n1288), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(new_n1305), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1293), .A2(new_n1288), .A3(new_n1304), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1354));
  INV_X1    g1154(.A(new_n1339), .ZN(new_n1355));
  XNOR2_X1  g1155(.A(new_n1354), .B(new_n1355), .ZN(G402));
endmodule


