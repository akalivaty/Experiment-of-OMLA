

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U554 ( .A1(G8), .A2(n713), .ZN(n773) );
  XNOR2_X1 U555 ( .A(n524), .B(n523), .ZN(n525) );
  INV_X1 U556 ( .A(KEYINPUT23), .ZN(n523) );
  NOR2_X1 U557 ( .A1(n768), .A2(n767), .ZN(n521) );
  OR2_X1 U558 ( .A1(n773), .A2(n763), .ZN(n522) );
  XNOR2_X1 U559 ( .A(KEYINPUT98), .B(KEYINPUT30), .ZN(n732) );
  XNOR2_X1 U560 ( .A(n733), .B(n732), .ZN(n734) );
  XNOR2_X1 U561 ( .A(KEYINPUT97), .B(KEYINPUT29), .ZN(n723) );
  XNOR2_X1 U562 ( .A(n724), .B(n723), .ZN(n730) );
  INV_X1 U563 ( .A(KEYINPUT99), .ZN(n743) );
  INV_X1 U564 ( .A(KEYINPUT33), .ZN(n764) );
  INV_X1 U565 ( .A(G2105), .ZN(n529) );
  XOR2_X1 U566 ( .A(KEYINPUT0), .B(G543), .Z(n635) );
  AND2_X2 U567 ( .A1(n529), .A2(G2104), .ZN(n897) );
  NOR2_X1 U568 ( .A1(G651), .A2(n635), .ZN(n663) );
  NOR2_X1 U569 ( .A1(n534), .A2(n533), .ZN(n695) );
  BUF_X1 U570 ( .A(n695), .Z(G160) );
  AND2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n893) );
  NAND2_X1 U572 ( .A1(n893), .A2(G113), .ZN(n526) );
  NAND2_X1 U573 ( .A1(G101), .A2(n897), .ZN(n524) );
  NAND2_X1 U574 ( .A1(n526), .A2(n525), .ZN(n534) );
  XNOR2_X1 U575 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n528) );
  NOR2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n527) );
  XNOR2_X1 U577 ( .A(n528), .B(n527), .ZN(n618) );
  NAND2_X1 U578 ( .A1(G137), .A2(n618), .ZN(n532) );
  NOR2_X1 U579 ( .A1(n529), .A2(G2104), .ZN(n530) );
  XNOR2_X1 U580 ( .A(n530), .B(KEYINPUT64), .ZN(n616) );
  NAND2_X1 U581 ( .A1(G125), .A2(n616), .ZN(n531) );
  NAND2_X1 U582 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U583 ( .A(G2443), .B(G2446), .Z(n536) );
  XNOR2_X1 U584 ( .A(G2427), .B(G2451), .ZN(n535) );
  XNOR2_X1 U585 ( .A(n536), .B(n535), .ZN(n542) );
  XOR2_X1 U586 ( .A(G2430), .B(G2454), .Z(n538) );
  XNOR2_X1 U587 ( .A(G1341), .B(G1348), .ZN(n537) );
  XNOR2_X1 U588 ( .A(n538), .B(n537), .ZN(n540) );
  XOR2_X1 U589 ( .A(G2435), .B(G2438), .Z(n539) );
  XNOR2_X1 U590 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U591 ( .A(n542), .B(n541), .Z(n543) );
  AND2_X1 U592 ( .A1(G14), .A2(n543), .ZN(G401) );
  AND2_X1 U593 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U594 ( .A(G120), .ZN(G236) );
  INV_X1 U595 ( .A(G69), .ZN(G235) );
  INV_X1 U596 ( .A(G108), .ZN(G238) );
  INV_X1 U597 ( .A(G82), .ZN(G220) );
  NOR2_X1 U598 ( .A1(G651), .A2(G543), .ZN(n658) );
  NAND2_X1 U599 ( .A1(G90), .A2(n658), .ZN(n546) );
  INV_X1 U600 ( .A(G651), .ZN(n550) );
  OR2_X1 U601 ( .A1(n550), .A2(n635), .ZN(n544) );
  XOR2_X2 U602 ( .A(n544), .B(KEYINPUT66), .Z(n657) );
  NAND2_X1 U603 ( .A1(G77), .A2(n657), .ZN(n545) );
  NAND2_X1 U604 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U605 ( .A(n547), .B(KEYINPUT9), .ZN(n549) );
  NAND2_X1 U606 ( .A1(G52), .A2(n663), .ZN(n548) );
  NAND2_X1 U607 ( .A1(n549), .A2(n548), .ZN(n554) );
  NOR2_X1 U608 ( .A1(G543), .A2(n550), .ZN(n551) );
  XOR2_X1 U609 ( .A(KEYINPUT1), .B(n551), .Z(n574) );
  BUF_X1 U610 ( .A(n574), .Z(n662) );
  NAND2_X1 U611 ( .A1(G64), .A2(n662), .ZN(n552) );
  XNOR2_X1 U612 ( .A(KEYINPUT69), .B(n552), .ZN(n553) );
  NOR2_X1 U613 ( .A1(n554), .A2(n553), .ZN(G171) );
  NAND2_X1 U614 ( .A1(G91), .A2(n658), .ZN(n556) );
  NAND2_X1 U615 ( .A1(G53), .A2(n663), .ZN(n555) );
  NAND2_X1 U616 ( .A1(n556), .A2(n555), .ZN(n559) );
  NAND2_X1 U617 ( .A1(n662), .A2(G65), .ZN(n557) );
  XOR2_X1 U618 ( .A(KEYINPUT70), .B(n557), .Z(n558) );
  NOR2_X1 U619 ( .A1(n559), .A2(n558), .ZN(n561) );
  NAND2_X1 U620 ( .A1(G78), .A2(n657), .ZN(n560) );
  NAND2_X1 U621 ( .A1(n561), .A2(n560), .ZN(G299) );
  NAND2_X1 U622 ( .A1(G138), .A2(n618), .ZN(n563) );
  NAND2_X1 U623 ( .A1(G102), .A2(n897), .ZN(n562) );
  NAND2_X1 U624 ( .A1(n563), .A2(n562), .ZN(n567) );
  NAND2_X1 U625 ( .A1(G114), .A2(n893), .ZN(n565) );
  NAND2_X1 U626 ( .A1(G126), .A2(n616), .ZN(n564) );
  NAND2_X1 U627 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U628 ( .A1(n567), .A2(n566), .ZN(G164) );
  NAND2_X1 U629 ( .A1(G7), .A2(G661), .ZN(n568) );
  XOR2_X1 U630 ( .A(n568), .B(KEYINPUT10), .Z(n832) );
  NAND2_X1 U631 ( .A1(n832), .A2(G567), .ZN(n569) );
  XOR2_X1 U632 ( .A(KEYINPUT11), .B(n569), .Z(G234) );
  NAND2_X1 U633 ( .A1(n658), .A2(G81), .ZN(n570) );
  XNOR2_X1 U634 ( .A(n570), .B(KEYINPUT12), .ZN(n572) );
  NAND2_X1 U635 ( .A1(G68), .A2(n657), .ZN(n571) );
  NAND2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U637 ( .A(n573), .B(KEYINPUT13), .ZN(n578) );
  NAND2_X1 U638 ( .A1(G56), .A2(n574), .ZN(n575) );
  XNOR2_X1 U639 ( .A(n575), .B(KEYINPUT72), .ZN(n576) );
  XNOR2_X1 U640 ( .A(KEYINPUT14), .B(n576), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U642 ( .A(n579), .B(KEYINPUT73), .ZN(n581) );
  NAND2_X1 U643 ( .A1(G43), .A2(n663), .ZN(n580) );
  NAND2_X1 U644 ( .A1(n581), .A2(n580), .ZN(n946) );
  INV_X1 U645 ( .A(G860), .ZN(n608) );
  OR2_X1 U646 ( .A1(n946), .A2(n608), .ZN(n582) );
  XNOR2_X1 U647 ( .A(KEYINPUT74), .B(n582), .ZN(G153) );
  INV_X1 U648 ( .A(G171), .ZN(G301) );
  NAND2_X1 U649 ( .A1(G868), .A2(G301), .ZN(n591) );
  NAND2_X1 U650 ( .A1(G92), .A2(n658), .ZN(n584) );
  NAND2_X1 U651 ( .A1(G79), .A2(n657), .ZN(n583) );
  NAND2_X1 U652 ( .A1(n584), .A2(n583), .ZN(n588) );
  NAND2_X1 U653 ( .A1(G66), .A2(n662), .ZN(n586) );
  NAND2_X1 U654 ( .A1(G54), .A2(n663), .ZN(n585) );
  NAND2_X1 U655 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U656 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U657 ( .A(KEYINPUT15), .B(n589), .ZN(n838) );
  INV_X1 U658 ( .A(G868), .ZN(n678) );
  NAND2_X1 U659 ( .A1(n838), .A2(n678), .ZN(n590) );
  NAND2_X1 U660 ( .A1(n591), .A2(n590), .ZN(G284) );
  XNOR2_X1 U661 ( .A(KEYINPUT7), .B(KEYINPUT76), .ZN(n603) );
  NAND2_X1 U662 ( .A1(n658), .A2(G89), .ZN(n592) );
  XNOR2_X1 U663 ( .A(n592), .B(KEYINPUT4), .ZN(n594) );
  NAND2_X1 U664 ( .A1(G76), .A2(n657), .ZN(n593) );
  NAND2_X1 U665 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U666 ( .A(KEYINPUT5), .B(n595), .ZN(n601) );
  NAND2_X1 U667 ( .A1(n662), .A2(G63), .ZN(n596) );
  XOR2_X1 U668 ( .A(KEYINPUT75), .B(n596), .Z(n598) );
  NAND2_X1 U669 ( .A1(n663), .A2(G51), .ZN(n597) );
  NAND2_X1 U670 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U671 ( .A(KEYINPUT6), .B(n599), .Z(n600) );
  NAND2_X1 U672 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U673 ( .A(n603), .B(n602), .ZN(G168) );
  XOR2_X1 U674 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  XOR2_X1 U675 ( .A(KEYINPUT77), .B(n678), .Z(n604) );
  NOR2_X1 U676 ( .A1(G286), .A2(n604), .ZN(n606) );
  NOR2_X1 U677 ( .A1(G868), .A2(G299), .ZN(n605) );
  NOR2_X1 U678 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U679 ( .A(KEYINPUT78), .B(n607), .ZN(G297) );
  NAND2_X1 U680 ( .A1(n608), .A2(G559), .ZN(n609) );
  INV_X1 U681 ( .A(n838), .ZN(n940) );
  NAND2_X1 U682 ( .A1(n609), .A2(n940), .ZN(n610) );
  XNOR2_X1 U683 ( .A(n610), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U684 ( .A1(G868), .A2(n946), .ZN(n613) );
  NAND2_X1 U685 ( .A1(G868), .A2(n940), .ZN(n611) );
  NOR2_X1 U686 ( .A1(G559), .A2(n611), .ZN(n612) );
  NOR2_X1 U687 ( .A1(n613), .A2(n612), .ZN(G282) );
  NAND2_X1 U688 ( .A1(G99), .A2(n897), .ZN(n615) );
  NAND2_X1 U689 ( .A1(G111), .A2(n893), .ZN(n614) );
  NAND2_X1 U690 ( .A1(n615), .A2(n614), .ZN(n623) );
  BUF_X1 U691 ( .A(n616), .Z(n894) );
  NAND2_X1 U692 ( .A1(n894), .A2(G123), .ZN(n617) );
  XNOR2_X1 U693 ( .A(n617), .B(KEYINPUT18), .ZN(n621) );
  INV_X1 U694 ( .A(n618), .ZN(n619) );
  INV_X1 U695 ( .A(n619), .ZN(n898) );
  NAND2_X1 U696 ( .A1(n898), .A2(G135), .ZN(n620) );
  NAND2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U698 ( .A1(n623), .A2(n622), .ZN(n999) );
  XNOR2_X1 U699 ( .A(n999), .B(G2096), .ZN(n624) );
  INV_X1 U700 ( .A(G2100), .ZN(n863) );
  NAND2_X1 U701 ( .A1(n624), .A2(n863), .ZN(G156) );
  NAND2_X1 U702 ( .A1(G93), .A2(n658), .ZN(n626) );
  NAND2_X1 U703 ( .A1(G80), .A2(n657), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U705 ( .A1(G67), .A2(n662), .ZN(n628) );
  NAND2_X1 U706 ( .A1(G55), .A2(n663), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n628), .A2(n627), .ZN(n629) );
  OR2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n677) );
  NAND2_X1 U709 ( .A1(G559), .A2(n940), .ZN(n631) );
  XNOR2_X1 U710 ( .A(n631), .B(n946), .ZN(n675) );
  NOR2_X1 U711 ( .A1(G860), .A2(n675), .ZN(n632) );
  XOR2_X1 U712 ( .A(KEYINPUT79), .B(n632), .Z(n633) );
  XOR2_X1 U713 ( .A(n677), .B(n633), .Z(G145) );
  NAND2_X1 U714 ( .A1(G49), .A2(n663), .ZN(n634) );
  XNOR2_X1 U715 ( .A(n634), .B(KEYINPUT80), .ZN(n640) );
  NAND2_X1 U716 ( .A1(G87), .A2(n635), .ZN(n637) );
  NAND2_X1 U717 ( .A1(G74), .A2(G651), .ZN(n636) );
  NAND2_X1 U718 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U719 ( .A1(n662), .A2(n638), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U721 ( .A(KEYINPUT81), .B(n641), .Z(G288) );
  NAND2_X1 U722 ( .A1(G88), .A2(n658), .ZN(n643) );
  NAND2_X1 U723 ( .A1(G75), .A2(n657), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U725 ( .A1(G62), .A2(n662), .ZN(n645) );
  NAND2_X1 U726 ( .A1(G50), .A2(n663), .ZN(n644) );
  NAND2_X1 U727 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U728 ( .A1(n647), .A2(n646), .ZN(G166) );
  INV_X1 U729 ( .A(G166), .ZN(G303) );
  NAND2_X1 U730 ( .A1(G86), .A2(n658), .ZN(n649) );
  NAND2_X1 U731 ( .A1(G61), .A2(n662), .ZN(n648) );
  NAND2_X1 U732 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U733 ( .A(KEYINPUT82), .B(n650), .ZN(n654) );
  NAND2_X1 U734 ( .A1(n657), .A2(G73), .ZN(n651) );
  XNOR2_X1 U735 ( .A(n651), .B(KEYINPUT2), .ZN(n652) );
  XNOR2_X1 U736 ( .A(n652), .B(KEYINPUT83), .ZN(n653) );
  NOR2_X1 U737 ( .A1(n654), .A2(n653), .ZN(n656) );
  NAND2_X1 U738 ( .A1(n663), .A2(G48), .ZN(n655) );
  NAND2_X1 U739 ( .A1(n656), .A2(n655), .ZN(G305) );
  NAND2_X1 U740 ( .A1(G72), .A2(n657), .ZN(n660) );
  NAND2_X1 U741 ( .A1(n658), .A2(G85), .ZN(n659) );
  NAND2_X1 U742 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U743 ( .A(KEYINPUT67), .B(n661), .ZN(n668) );
  NAND2_X1 U744 ( .A1(G60), .A2(n662), .ZN(n665) );
  NAND2_X1 U745 ( .A1(G47), .A2(n663), .ZN(n664) );
  NAND2_X1 U746 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U747 ( .A(KEYINPUT68), .B(n666), .Z(n667) );
  NAND2_X1 U748 ( .A1(n668), .A2(n667), .ZN(G290) );
  XNOR2_X1 U749 ( .A(KEYINPUT19), .B(KEYINPUT84), .ZN(n670) );
  XOR2_X1 U750 ( .A(G288), .B(G303), .Z(n669) );
  XNOR2_X1 U751 ( .A(n670), .B(n669), .ZN(n671) );
  XOR2_X1 U752 ( .A(n677), .B(n671), .Z(n673) );
  XOR2_X1 U753 ( .A(G305), .B(G299), .Z(n672) );
  XNOR2_X1 U754 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U755 ( .A(n674), .B(G290), .ZN(n840) );
  XNOR2_X1 U756 ( .A(n675), .B(n840), .ZN(n676) );
  NAND2_X1 U757 ( .A1(n676), .A2(G868), .ZN(n680) );
  NAND2_X1 U758 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U759 ( .A1(n680), .A2(n679), .ZN(G295) );
  NAND2_X1 U760 ( .A1(G2084), .A2(G2078), .ZN(n681) );
  XOR2_X1 U761 ( .A(KEYINPUT20), .B(n681), .Z(n682) );
  NAND2_X1 U762 ( .A1(G2090), .A2(n682), .ZN(n683) );
  XNOR2_X1 U763 ( .A(KEYINPUT21), .B(n683), .ZN(n684) );
  NAND2_X1 U764 ( .A1(n684), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U765 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U766 ( .A(KEYINPUT71), .B(G132), .ZN(G219) );
  NOR2_X1 U767 ( .A1(G220), .A2(G219), .ZN(n685) );
  XOR2_X1 U768 ( .A(KEYINPUT22), .B(n685), .Z(n686) );
  NOR2_X1 U769 ( .A1(G218), .A2(n686), .ZN(n687) );
  NAND2_X1 U770 ( .A1(G96), .A2(n687), .ZN(n837) );
  NAND2_X1 U771 ( .A1(n837), .A2(G2106), .ZN(n693) );
  NOR2_X1 U772 ( .A1(G235), .A2(G236), .ZN(n688) );
  XNOR2_X1 U773 ( .A(n688), .B(KEYINPUT85), .ZN(n689) );
  NOR2_X1 U774 ( .A1(G238), .A2(n689), .ZN(n690) );
  NAND2_X1 U775 ( .A1(G57), .A2(n690), .ZN(n836) );
  NAND2_X1 U776 ( .A1(G567), .A2(n836), .ZN(n691) );
  XNOR2_X1 U777 ( .A(KEYINPUT86), .B(n691), .ZN(n692) );
  NAND2_X1 U778 ( .A1(n693), .A2(n692), .ZN(n917) );
  NAND2_X1 U779 ( .A1(G483), .A2(G661), .ZN(n694) );
  NOR2_X1 U780 ( .A1(n917), .A2(n694), .ZN(n835) );
  NAND2_X1 U781 ( .A1(n835), .A2(G36), .ZN(G176) );
  NOR2_X1 U782 ( .A1(G164), .A2(G1384), .ZN(n782) );
  INV_X1 U783 ( .A(n782), .ZN(n696) );
  NAND2_X1 U784 ( .A1(n695), .A2(G40), .ZN(n781) );
  NOR2_X1 U785 ( .A1(n696), .A2(n781), .ZN(n725) );
  INV_X1 U786 ( .A(n725), .ZN(n713) );
  NOR2_X1 U787 ( .A1(G1981), .A2(G305), .ZN(n697) );
  XOR2_X1 U788 ( .A(n697), .B(KEYINPUT24), .Z(n698) );
  NOR2_X1 U789 ( .A1(n773), .A2(n698), .ZN(n780) );
  INV_X1 U790 ( .A(G1996), .ZN(n847) );
  NOR2_X1 U791 ( .A1(n713), .A2(n847), .ZN(n699) );
  XOR2_X1 U792 ( .A(n699), .B(KEYINPUT26), .Z(n701) );
  BUF_X1 U793 ( .A(n713), .Z(n749) );
  NAND2_X1 U794 ( .A1(n749), .A2(G1341), .ZN(n700) );
  NAND2_X1 U795 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U796 ( .A1(n946), .A2(n702), .ZN(n703) );
  OR2_X1 U797 ( .A1(n940), .A2(n703), .ZN(n710) );
  NAND2_X1 U798 ( .A1(n940), .A2(n703), .ZN(n708) );
  NAND2_X1 U799 ( .A1(G1348), .A2(n749), .ZN(n705) );
  NAND2_X1 U800 ( .A1(G2067), .A2(n725), .ZN(n704) );
  NAND2_X1 U801 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U802 ( .A(KEYINPUT96), .B(n706), .ZN(n707) );
  NAND2_X1 U803 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U804 ( .A1(n710), .A2(n709), .ZN(n717) );
  INV_X1 U805 ( .A(G299), .ZN(n718) );
  AND2_X1 U806 ( .A1(G2072), .A2(n725), .ZN(n711) );
  XNOR2_X1 U807 ( .A(n711), .B(KEYINPUT95), .ZN(n712) );
  XNOR2_X1 U808 ( .A(n712), .B(KEYINPUT27), .ZN(n715) );
  AND2_X1 U809 ( .A1(n713), .A2(G1956), .ZN(n714) );
  NOR2_X1 U810 ( .A1(n715), .A2(n714), .ZN(n719) );
  NAND2_X1 U811 ( .A1(n718), .A2(n719), .ZN(n716) );
  NAND2_X1 U812 ( .A1(n717), .A2(n716), .ZN(n722) );
  NOR2_X1 U813 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U814 ( .A(n720), .B(KEYINPUT28), .Z(n721) );
  NAND2_X1 U815 ( .A1(n722), .A2(n721), .ZN(n724) );
  INV_X1 U816 ( .A(G1961), .ZN(n850) );
  NAND2_X1 U817 ( .A1(n749), .A2(n850), .ZN(n727) );
  XNOR2_X1 U818 ( .A(G2078), .B(KEYINPUT25), .ZN(n923) );
  NAND2_X1 U819 ( .A1(n725), .A2(n923), .ZN(n726) );
  NAND2_X1 U820 ( .A1(n727), .A2(n726), .ZN(n735) );
  AND2_X1 U821 ( .A1(n735), .A2(G171), .ZN(n728) );
  XOR2_X1 U822 ( .A(KEYINPUT94), .B(n728), .Z(n729) );
  NAND2_X1 U823 ( .A1(n730), .A2(n729), .ZN(n740) );
  NOR2_X1 U824 ( .A1(G2084), .A2(n749), .ZN(n745) );
  NOR2_X1 U825 ( .A1(G1966), .A2(n773), .ZN(n741) );
  NOR2_X1 U826 ( .A1(n745), .A2(n741), .ZN(n731) );
  NAND2_X1 U827 ( .A1(G8), .A2(n731), .ZN(n733) );
  NOR2_X1 U828 ( .A1(G168), .A2(n734), .ZN(n737) );
  NOR2_X1 U829 ( .A1(G171), .A2(n735), .ZN(n736) );
  NOR2_X1 U830 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U831 ( .A(KEYINPUT31), .B(n738), .Z(n739) );
  NAND2_X1 U832 ( .A1(n740), .A2(n739), .ZN(n748) );
  INV_X1 U833 ( .A(n748), .ZN(n742) );
  NOR2_X1 U834 ( .A1(n742), .A2(n741), .ZN(n744) );
  XNOR2_X1 U835 ( .A(n744), .B(n743), .ZN(n747) );
  NAND2_X1 U836 ( .A1(G8), .A2(n745), .ZN(n746) );
  NAND2_X1 U837 ( .A1(n747), .A2(n746), .ZN(n758) );
  NAND2_X1 U838 ( .A1(n748), .A2(G286), .ZN(n754) );
  NOR2_X1 U839 ( .A1(G1971), .A2(n773), .ZN(n751) );
  NOR2_X1 U840 ( .A1(G2090), .A2(n749), .ZN(n750) );
  NOR2_X1 U841 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U842 ( .A1(n752), .A2(G303), .ZN(n753) );
  NAND2_X1 U843 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U844 ( .A1(n755), .A2(G8), .ZN(n756) );
  XNOR2_X1 U845 ( .A(KEYINPUT32), .B(n756), .ZN(n757) );
  NAND2_X1 U846 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U847 ( .A(KEYINPUT100), .B(n759), .ZN(n771) );
  NOR2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n765) );
  NOR2_X1 U849 ( .A1(G1971), .A2(G303), .ZN(n760) );
  NOR2_X1 U850 ( .A1(n765), .A2(n760), .ZN(n948) );
  NAND2_X1 U851 ( .A1(n771), .A2(n948), .ZN(n762) );
  NAND2_X1 U852 ( .A1(G288), .A2(G1976), .ZN(n761) );
  XOR2_X1 U853 ( .A(KEYINPUT101), .B(n761), .Z(n947) );
  NAND2_X1 U854 ( .A1(n762), .A2(n947), .ZN(n763) );
  NAND2_X1 U855 ( .A1(n522), .A2(n764), .ZN(n769) );
  XOR2_X1 U856 ( .A(G1981), .B(G305), .Z(n959) );
  INV_X1 U857 ( .A(n959), .ZN(n768) );
  NAND2_X1 U858 ( .A1(n765), .A2(KEYINPUT33), .ZN(n766) );
  NOR2_X1 U859 ( .A1(n766), .A2(n773), .ZN(n767) );
  NAND2_X1 U860 ( .A1(n769), .A2(n521), .ZN(n777) );
  NOR2_X1 U861 ( .A1(G2090), .A2(G303), .ZN(n770) );
  NAND2_X1 U862 ( .A1(G8), .A2(n770), .ZN(n772) );
  NAND2_X1 U863 ( .A1(n772), .A2(n771), .ZN(n774) );
  NAND2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U865 ( .A(n775), .B(KEYINPUT102), .ZN(n776) );
  NAND2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U867 ( .A(KEYINPUT103), .B(n778), .Z(n779) );
  NOR2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n814) );
  NOR2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n827) );
  NAND2_X1 U870 ( .A1(n898), .A2(G140), .ZN(n783) );
  XOR2_X1 U871 ( .A(KEYINPUT87), .B(n783), .Z(n785) );
  NAND2_X1 U872 ( .A1(n897), .A2(G104), .ZN(n784) );
  NAND2_X1 U873 ( .A1(n785), .A2(n784), .ZN(n787) );
  XNOR2_X1 U874 ( .A(KEYINPUT88), .B(KEYINPUT34), .ZN(n786) );
  XNOR2_X1 U875 ( .A(n787), .B(n786), .ZN(n792) );
  NAND2_X1 U876 ( .A1(G116), .A2(n893), .ZN(n789) );
  NAND2_X1 U877 ( .A1(G128), .A2(n894), .ZN(n788) );
  NAND2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U879 ( .A(KEYINPUT35), .B(n790), .Z(n791) );
  NOR2_X1 U880 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U881 ( .A(KEYINPUT36), .B(n793), .ZN(n907) );
  XNOR2_X1 U882 ( .A(KEYINPUT37), .B(G2067), .ZN(n825) );
  NOR2_X1 U883 ( .A1(n907), .A2(n825), .ZN(n1020) );
  NAND2_X1 U884 ( .A1(n827), .A2(n1020), .ZN(n823) );
  NAND2_X1 U885 ( .A1(G95), .A2(n897), .ZN(n795) );
  NAND2_X1 U886 ( .A1(G119), .A2(n894), .ZN(n794) );
  NAND2_X1 U887 ( .A1(n795), .A2(n794), .ZN(n798) );
  NAND2_X1 U888 ( .A1(G107), .A2(n893), .ZN(n796) );
  XNOR2_X1 U889 ( .A(KEYINPUT89), .B(n796), .ZN(n797) );
  NOR2_X1 U890 ( .A1(n798), .A2(n797), .ZN(n800) );
  NAND2_X1 U891 ( .A1(n898), .A2(G131), .ZN(n799) );
  NAND2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n889) );
  XNOR2_X1 U893 ( .A(KEYINPUT90), .B(G1991), .ZN(n922) );
  AND2_X1 U894 ( .A1(n889), .A2(n922), .ZN(n801) );
  XNOR2_X1 U895 ( .A(n801), .B(KEYINPUT91), .ZN(n811) );
  NAND2_X1 U896 ( .A1(G105), .A2(n897), .ZN(n802) );
  XNOR2_X1 U897 ( .A(n802), .B(KEYINPUT38), .ZN(n809) );
  NAND2_X1 U898 ( .A1(G141), .A2(n898), .ZN(n804) );
  NAND2_X1 U899 ( .A1(G129), .A2(n894), .ZN(n803) );
  NAND2_X1 U900 ( .A1(n804), .A2(n803), .ZN(n807) );
  NAND2_X1 U901 ( .A1(n893), .A2(G117), .ZN(n805) );
  XOR2_X1 U902 ( .A(KEYINPUT92), .B(n805), .Z(n806) );
  NOR2_X1 U903 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n890) );
  NAND2_X1 U905 ( .A1(G1996), .A2(n890), .ZN(n810) );
  NAND2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n812) );
  XOR2_X1 U907 ( .A(KEYINPUT93), .B(n812), .Z(n998) );
  NAND2_X1 U908 ( .A1(n998), .A2(n827), .ZN(n817) );
  NAND2_X1 U909 ( .A1(n823), .A2(n817), .ZN(n813) );
  NOR2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n816) );
  XNOR2_X1 U911 ( .A(G1986), .B(G290), .ZN(n945) );
  NAND2_X1 U912 ( .A1(n945), .A2(n827), .ZN(n815) );
  NAND2_X1 U913 ( .A1(n816), .A2(n815), .ZN(n830) );
  NOR2_X1 U914 ( .A1(G1996), .A2(n890), .ZN(n1004) );
  INV_X1 U915 ( .A(n817), .ZN(n820) );
  NOR2_X1 U916 ( .A1(n889), .A2(n922), .ZN(n1000) );
  NOR2_X1 U917 ( .A1(G1986), .A2(G290), .ZN(n818) );
  NOR2_X1 U918 ( .A1(n1000), .A2(n818), .ZN(n819) );
  NOR2_X1 U919 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U920 ( .A1(n1004), .A2(n821), .ZN(n822) );
  XNOR2_X1 U921 ( .A(n822), .B(KEYINPUT39), .ZN(n824) );
  NAND2_X1 U922 ( .A1(n824), .A2(n823), .ZN(n826) );
  NAND2_X1 U923 ( .A1(n907), .A2(n825), .ZN(n1017) );
  NAND2_X1 U924 ( .A1(n826), .A2(n1017), .ZN(n828) );
  NAND2_X1 U925 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U926 ( .A1(n830), .A2(n829), .ZN(n831) );
  XNOR2_X1 U927 ( .A(KEYINPUT40), .B(n831), .ZN(G329) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n832), .ZN(G217) );
  INV_X1 U929 ( .A(n832), .ZN(G223) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U931 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U933 ( .A1(n835), .A2(n834), .ZN(G188) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  NOR2_X1 U936 ( .A1(n837), .A2(n836), .ZN(G325) );
  INV_X1 U937 ( .A(G325), .ZN(G261) );
  XOR2_X1 U938 ( .A(n838), .B(G301), .Z(n839) );
  XNOR2_X1 U939 ( .A(n839), .B(G286), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n946), .B(n840), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n843) );
  NOR2_X1 U942 ( .A1(G37), .A2(n843), .ZN(G397) );
  XOR2_X1 U943 ( .A(KEYINPUT107), .B(G1971), .Z(n845) );
  XNOR2_X1 U944 ( .A(G1986), .B(G1976), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U946 ( .A(n846), .B(KEYINPUT41), .Z(n849) );
  XOR2_X1 U947 ( .A(n847), .B(G1991), .Z(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n854) );
  XNOR2_X1 U949 ( .A(n850), .B(G1956), .ZN(n852) );
  XNOR2_X1 U950 ( .A(G1981), .B(G1966), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U952 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U953 ( .A(G2474), .B(KEYINPUT106), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(G229) );
  XOR2_X1 U955 ( .A(KEYINPUT105), .B(KEYINPUT104), .Z(n858) );
  XNOR2_X1 U956 ( .A(G2678), .B(KEYINPUT43), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U958 ( .A(KEYINPUT42), .B(G2090), .Z(n860) );
  XNOR2_X1 U959 ( .A(G2067), .B(G2072), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U961 ( .A(n862), .B(n861), .Z(n865) );
  XOR2_X1 U962 ( .A(G2096), .B(n863), .Z(n864) );
  XNOR2_X1 U963 ( .A(n865), .B(n864), .ZN(n867) );
  XOR2_X1 U964 ( .A(G2084), .B(G2078), .Z(n866) );
  XNOR2_X1 U965 ( .A(n867), .B(n866), .ZN(G227) );
  NAND2_X1 U966 ( .A1(G100), .A2(n897), .ZN(n869) );
  NAND2_X1 U967 ( .A1(G112), .A2(n893), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n875) );
  NAND2_X1 U969 ( .A1(n894), .A2(G124), .ZN(n870) );
  XNOR2_X1 U970 ( .A(n870), .B(KEYINPUT44), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n871), .B(KEYINPUT108), .ZN(n873) );
  NAND2_X1 U972 ( .A1(G136), .A2(n898), .ZN(n872) );
  NAND2_X1 U973 ( .A1(n873), .A2(n872), .ZN(n874) );
  NOR2_X1 U974 ( .A1(n875), .A2(n874), .ZN(G162) );
  NAND2_X1 U975 ( .A1(G103), .A2(n897), .ZN(n877) );
  NAND2_X1 U976 ( .A1(G139), .A2(n898), .ZN(n876) );
  NAND2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n882) );
  NAND2_X1 U978 ( .A1(G115), .A2(n893), .ZN(n879) );
  NAND2_X1 U979 ( .A1(G127), .A2(n894), .ZN(n878) );
  NAND2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U981 ( .A(KEYINPUT47), .B(n880), .Z(n881) );
  NOR2_X1 U982 ( .A1(n882), .A2(n881), .ZN(n1011) );
  XOR2_X1 U983 ( .A(KEYINPUT48), .B(KEYINPUT111), .Z(n884) );
  XNOR2_X1 U984 ( .A(G164), .B(KEYINPUT46), .ZN(n883) );
  XNOR2_X1 U985 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U986 ( .A(n885), .B(n999), .Z(n887) );
  XNOR2_X1 U987 ( .A(G160), .B(G162), .ZN(n886) );
  XNOR2_X1 U988 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U989 ( .A(n1011), .B(n888), .ZN(n892) );
  XOR2_X1 U990 ( .A(n890), .B(n889), .Z(n891) );
  XNOR2_X1 U991 ( .A(n892), .B(n891), .ZN(n909) );
  NAND2_X1 U992 ( .A1(G118), .A2(n893), .ZN(n896) );
  NAND2_X1 U993 ( .A1(G130), .A2(n894), .ZN(n895) );
  NAND2_X1 U994 ( .A1(n896), .A2(n895), .ZN(n905) );
  XNOR2_X1 U995 ( .A(KEYINPUT45), .B(KEYINPUT110), .ZN(n903) );
  NAND2_X1 U996 ( .A1(n897), .A2(G106), .ZN(n901) );
  NAND2_X1 U997 ( .A1(n898), .A2(G142), .ZN(n899) );
  XOR2_X1 U998 ( .A(KEYINPUT109), .B(n899), .Z(n900) );
  NAND2_X1 U999 ( .A1(n901), .A2(n900), .ZN(n902) );
  XOR2_X1 U1000 ( .A(n903), .B(n902), .Z(n904) );
  NOR2_X1 U1001 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n910), .ZN(G395) );
  NOR2_X1 U1005 ( .A1(G229), .A2(G227), .ZN(n911) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(n911), .ZN(n912) );
  NOR2_X1 U1007 ( .A1(G397), .A2(n912), .ZN(n916) );
  NOR2_X1 U1008 ( .A1(n917), .A2(G401), .ZN(n913) );
  XOR2_X1 U1009 ( .A(KEYINPUT112), .B(n913), .Z(n914) );
  NOR2_X1 U1010 ( .A1(G395), .A2(n914), .ZN(n915) );
  NAND2_X1 U1011 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(n917), .ZN(G319) );
  INV_X1 U1014 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1015 ( .A(G2084), .B(G34), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(n918), .B(KEYINPUT54), .ZN(n936) );
  XOR2_X1 U1017 ( .A(G32), .B(G1996), .Z(n919) );
  NAND2_X1 U1018 ( .A1(n919), .A2(G28), .ZN(n929) );
  XNOR2_X1 U1019 ( .A(G2067), .B(G26), .ZN(n921) );
  XNOR2_X1 U1020 ( .A(G33), .B(G2072), .ZN(n920) );
  NOR2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n927) );
  XNOR2_X1 U1022 ( .A(n922), .B(G25), .ZN(n925) );
  XOR2_X1 U1023 ( .A(n923), .B(G27), .Z(n924) );
  NOR2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1027 ( .A(KEYINPUT114), .B(n930), .Z(n931) );
  XOR2_X1 U1028 ( .A(KEYINPUT53), .B(n931), .Z(n933) );
  XNOR2_X1 U1029 ( .A(G2090), .B(G35), .ZN(n932) );
  NOR2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1031 ( .A(n934), .B(KEYINPUT115), .ZN(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1033 ( .A(KEYINPUT55), .B(n937), .Z(n938) );
  XNOR2_X1 U1034 ( .A(KEYINPUT116), .B(n938), .ZN(n939) );
  NOR2_X1 U1035 ( .A1(G29), .A2(n939), .ZN(n996) );
  XOR2_X1 U1036 ( .A(n940), .B(G1348), .Z(n942) );
  XOR2_X1 U1037 ( .A(G171), .B(G1961), .Z(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1039 ( .A(n943), .B(KEYINPUT119), .ZN(n944) );
  NOR2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n958) );
  XNOR2_X1 U1041 ( .A(n946), .B(G1341), .ZN(n956) );
  AND2_X1 U1042 ( .A1(G303), .A2(G1971), .ZN(n950) );
  NAND2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1045 ( .A(KEYINPUT120), .B(n951), .Z(n953) );
  XNOR2_X1 U1046 ( .A(G299), .B(G1956), .ZN(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(KEYINPUT121), .B(n954), .ZN(n955) );
  NOR2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1050 ( .A1(n958), .A2(n957), .ZN(n964) );
  XNOR2_X1 U1051 ( .A(G1966), .B(G168), .ZN(n960) );
  NAND2_X1 U1052 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1053 ( .A(KEYINPUT57), .B(n961), .Z(n962) );
  XNOR2_X1 U1054 ( .A(KEYINPUT118), .B(n962), .ZN(n963) );
  NOR2_X1 U1055 ( .A1(n964), .A2(n963), .ZN(n967) );
  XNOR2_X1 U1056 ( .A(G16), .B(KEYINPUT56), .ZN(n965) );
  XNOR2_X1 U1057 ( .A(KEYINPUT117), .B(n965), .ZN(n966) );
  NOR2_X1 U1058 ( .A1(n967), .A2(n966), .ZN(n993) );
  XOR2_X1 U1059 ( .A(G1966), .B(G21), .Z(n975) );
  XNOR2_X1 U1060 ( .A(G1986), .B(G24), .ZN(n972) );
  XNOR2_X1 U1061 ( .A(G1976), .B(G23), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(G22), .B(G1971), .ZN(n968) );
  NOR2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(KEYINPUT123), .B(n970), .ZN(n971) );
  NOR2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1066 ( .A(KEYINPUT58), .B(n973), .ZN(n974) );
  NAND2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n987) );
  XOR2_X1 U1068 ( .A(G20), .B(G1956), .Z(n979) );
  XNOR2_X1 U1069 ( .A(G1981), .B(G6), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(G19), .B(G1341), .ZN(n976) );
  NOR2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n982) );
  XOR2_X1 U1073 ( .A(KEYINPUT59), .B(G1348), .Z(n980) );
  XNOR2_X1 U1074 ( .A(G4), .B(n980), .ZN(n981) );
  NOR2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(n983), .B(KEYINPUT60), .ZN(n985) );
  XOR2_X1 U1077 ( .A(G1961), .B(G5), .Z(n984) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1080 ( .A(KEYINPUT61), .B(n988), .Z(n990) );
  XNOR2_X1 U1081 ( .A(G16), .B(KEYINPUT122), .ZN(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(KEYINPUT124), .B(n991), .ZN(n992) );
  NOR2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(G11), .A2(n994), .ZN(n995) );
  NOR2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(n997), .B(KEYINPUT125), .ZN(n1026) );
  INV_X1 U1088 ( .A(G29), .ZN(n1024) );
  INV_X1 U1089 ( .A(n998), .ZN(n1010) );
  XNOR2_X1 U1090 ( .A(G160), .B(G2084), .ZN(n1002) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1008) );
  XOR2_X1 U1093 ( .A(G2090), .B(G162), .Z(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1095 ( .A(KEYINPUT51), .B(n1005), .Z(n1006) );
  XNOR2_X1 U1096 ( .A(n1006), .B(KEYINPUT113), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1016) );
  XOR2_X1 U1099 ( .A(G2072), .B(n1011), .Z(n1013) );
  XOR2_X1 U1100 ( .A(G164), .B(G2078), .Z(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1102 ( .A(KEYINPUT50), .B(n1014), .Z(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1106 ( .A(KEYINPUT52), .B(n1021), .Z(n1022) );
  NOR2_X1 U1107 ( .A1(KEYINPUT55), .A2(n1022), .ZN(n1023) );
  NOR2_X1 U1108 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1109 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1110 ( .A(n1027), .B(KEYINPUT62), .ZN(n1028) );
  XNOR2_X1 U1111 ( .A(n1028), .B(KEYINPUT126), .ZN(G311) );
  XNOR2_X1 U1112 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

