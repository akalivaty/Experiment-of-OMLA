

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578;

  NOR2_X1 U318 ( .A1(n493), .A2(n437), .ZN(n557) );
  INV_X1 U319 ( .A(KEYINPUT32), .ZN(n375) );
  XNOR2_X1 U320 ( .A(n376), .B(n375), .ZN(n377) );
  NOR2_X1 U321 ( .A1(n491), .A2(n516), .ZN(n399) );
  XNOR2_X1 U322 ( .A(n378), .B(n377), .ZN(n382) );
  NOR2_X1 U323 ( .A1(n562), .A2(n448), .ZN(n435) );
  INV_X1 U324 ( .A(G190GAT), .ZN(n438) );
  XNOR2_X1 U325 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U326 ( .A(n441), .B(n440), .ZN(G1351GAT) );
  XOR2_X1 U327 ( .A(G120GAT), .B(G71GAT), .Z(n384) );
  XOR2_X1 U328 ( .A(G99GAT), .B(G190GAT), .Z(n287) );
  XNOR2_X1 U329 ( .A(G43GAT), .B(G15GAT), .ZN(n286) );
  XNOR2_X1 U330 ( .A(n287), .B(n286), .ZN(n288) );
  XOR2_X1 U331 ( .A(n384), .B(n288), .Z(n290) );
  NAND2_X1 U332 ( .A1(G227GAT), .A2(G233GAT), .ZN(n289) );
  XNOR2_X1 U333 ( .A(n290), .B(n289), .ZN(n304) );
  XOR2_X1 U334 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n292) );
  XNOR2_X1 U335 ( .A(G169GAT), .B(KEYINPUT20), .ZN(n291) );
  XNOR2_X1 U336 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U337 ( .A(G176GAT), .B(KEYINPUT65), .Z(n294) );
  XNOR2_X1 U338 ( .A(KEYINPUT83), .B(KEYINPUT86), .ZN(n293) );
  XNOR2_X1 U339 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U340 ( .A(n296), .B(n295), .Z(n302) );
  XOR2_X1 U341 ( .A(G127GAT), .B(KEYINPUT0), .Z(n298) );
  XNOR2_X1 U342 ( .A(G113GAT), .B(G134GAT), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n408) );
  XOR2_X1 U344 ( .A(G183GAT), .B(KEYINPUT17), .Z(n300) );
  XNOR2_X1 U345 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n315) );
  XNOR2_X1 U347 ( .A(n408), .B(n315), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U349 ( .A(n304), .B(n303), .ZN(n517) );
  INV_X1 U350 ( .A(n517), .ZN(n493) );
  XOR2_X1 U351 ( .A(KEYINPUT55), .B(KEYINPUT119), .Z(n436) );
  XOR2_X1 U352 ( .A(G211GAT), .B(KEYINPUT21), .Z(n306) );
  XNOR2_X1 U353 ( .A(G197GAT), .B(G218GAT), .ZN(n305) );
  XNOR2_X1 U354 ( .A(n306), .B(n305), .ZN(n428) );
  XOR2_X1 U355 ( .A(KEYINPUT92), .B(n428), .Z(n308) );
  NAND2_X1 U356 ( .A1(G226GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U358 ( .A(G36GAT), .B(G190GAT), .Z(n321) );
  XOR2_X1 U359 ( .A(n309), .B(n321), .Z(n313) );
  XOR2_X1 U360 ( .A(G169GAT), .B(G8GAT), .Z(n363) );
  XOR2_X1 U361 ( .A(G64GAT), .B(G92GAT), .Z(n311) );
  XNOR2_X1 U362 ( .A(G176GAT), .B(G204GAT), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n370) );
  XNOR2_X1 U364 ( .A(n363), .B(n370), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U366 ( .A(n315), .B(n314), .Z(n506) );
  INV_X1 U367 ( .A(n506), .ZN(n491) );
  XOR2_X1 U368 ( .A(KEYINPUT10), .B(KEYINPUT76), .Z(n317) );
  XNOR2_X1 U369 ( .A(G92GAT), .B(KEYINPUT11), .ZN(n316) );
  XNOR2_X1 U370 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U371 ( .A(G99GAT), .B(G85GAT), .Z(n369) );
  XOR2_X1 U372 ( .A(n318), .B(n369), .Z(n320) );
  XNOR2_X1 U373 ( .A(G218GAT), .B(G106GAT), .ZN(n319) );
  XNOR2_X1 U374 ( .A(n320), .B(n319), .ZN(n322) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U376 ( .A(G29GAT), .B(G43GAT), .Z(n324) );
  XNOR2_X1 U377 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n324), .B(n323), .ZN(n360) );
  XOR2_X1 U379 ( .A(G50GAT), .B(G162GAT), .Z(n421) );
  XOR2_X1 U380 ( .A(n360), .B(n421), .Z(n325) );
  XNOR2_X1 U381 ( .A(n326), .B(n325), .ZN(n330) );
  XOR2_X1 U382 ( .A(KEYINPUT75), .B(KEYINPUT66), .Z(n328) );
  NAND2_X1 U383 ( .A1(G232GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U384 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n330), .B(n329), .ZN(n335) );
  XOR2_X1 U386 ( .A(KEYINPUT77), .B(KEYINPUT74), .Z(n332) );
  XNOR2_X1 U387 ( .A(KEYINPUT67), .B(KEYINPUT9), .ZN(n331) );
  XNOR2_X1 U388 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U389 ( .A(G134GAT), .B(n333), .ZN(n334) );
  XNOR2_X1 U390 ( .A(n335), .B(n334), .ZN(n531) );
  INV_X1 U391 ( .A(n531), .ZN(n548) );
  XNOR2_X1 U392 ( .A(G22GAT), .B(G15GAT), .ZN(n336) );
  XNOR2_X1 U393 ( .A(n336), .B(G1GAT), .ZN(n359) );
  XOR2_X1 U394 ( .A(n359), .B(KEYINPUT78), .Z(n338) );
  NAND2_X1 U395 ( .A1(G231GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n338), .B(n337), .ZN(n353) );
  XOR2_X1 U397 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n340) );
  XNOR2_X1 U398 ( .A(G8GAT), .B(G64GAT), .ZN(n339) );
  XNOR2_X1 U399 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U400 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n342) );
  XNOR2_X1 U401 ( .A(KEYINPUT12), .B(KEYINPUT81), .ZN(n341) );
  XNOR2_X1 U402 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U403 ( .A(n344), .B(n343), .ZN(n351) );
  XOR2_X1 U404 ( .A(G211GAT), .B(G155GAT), .Z(n346) );
  XNOR2_X1 U405 ( .A(G183GAT), .B(G71GAT), .ZN(n345) );
  XNOR2_X1 U406 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U407 ( .A(G57GAT), .B(KEYINPUT13), .Z(n383) );
  XOR2_X1 U408 ( .A(n347), .B(n383), .Z(n349) );
  XNOR2_X1 U409 ( .A(G127GAT), .B(G78GAT), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U411 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U412 ( .A(n353), .B(n352), .Z(n572) );
  INV_X1 U413 ( .A(n572), .ZN(n545) );
  NAND2_X1 U414 ( .A1(n548), .A2(n545), .ZN(n391) );
  XNOR2_X1 U415 ( .A(KEYINPUT110), .B(KEYINPUT46), .ZN(n389) );
  XOR2_X1 U416 ( .A(KEYINPUT30), .B(G113GAT), .Z(n355) );
  XNOR2_X1 U417 ( .A(G197GAT), .B(G141GAT), .ZN(n354) );
  XNOR2_X1 U418 ( .A(n355), .B(n354), .ZN(n368) );
  XOR2_X1 U419 ( .A(KEYINPUT29), .B(KEYINPUT69), .Z(n357) );
  NAND2_X1 U420 ( .A1(G229GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U421 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U422 ( .A(n358), .B(KEYINPUT68), .Z(n362) );
  XNOR2_X1 U423 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U424 ( .A(n362), .B(n361), .ZN(n364) );
  XOR2_X1 U425 ( .A(n364), .B(n363), .Z(n366) );
  XNOR2_X1 U426 ( .A(G50GAT), .B(G36GAT), .ZN(n365) );
  XNOR2_X1 U427 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U428 ( .A(n368), .B(n367), .ZN(n563) );
  INV_X1 U429 ( .A(n563), .ZN(n537) );
  XOR2_X1 U430 ( .A(n370), .B(n369), .Z(n372) );
  NAND2_X1 U431 ( .A1(G230GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U432 ( .A(n372), .B(n371), .ZN(n378) );
  XOR2_X1 U433 ( .A(G78GAT), .B(G148GAT), .Z(n374) );
  XNOR2_X1 U434 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n374), .B(n373), .ZN(n427) );
  XNOR2_X1 U436 ( .A(n427), .B(KEYINPUT31), .ZN(n376) );
  XOR2_X1 U437 ( .A(KEYINPUT70), .B(KEYINPUT72), .Z(n380) );
  XNOR2_X1 U438 ( .A(KEYINPUT73), .B(KEYINPUT33), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U440 ( .A(n382), .B(n381), .Z(n386) );
  XNOR2_X1 U441 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n386), .B(n385), .ZN(n568) );
  XOR2_X1 U443 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n387) );
  XNOR2_X1 U444 ( .A(n568), .B(n387), .ZN(n542) );
  NOR2_X1 U445 ( .A1(n537), .A2(n542), .ZN(n388) );
  XNOR2_X1 U446 ( .A(n389), .B(n388), .ZN(n390) );
  NOR2_X1 U447 ( .A1(n391), .A2(n390), .ZN(n392) );
  XNOR2_X1 U448 ( .A(n392), .B(KEYINPUT47), .ZN(n397) );
  XOR2_X1 U449 ( .A(KEYINPUT36), .B(n531), .Z(n576) );
  NOR2_X1 U450 ( .A1(n576), .A2(n545), .ZN(n393) );
  XOR2_X1 U451 ( .A(KEYINPUT45), .B(n393), .Z(n394) );
  NOR2_X1 U452 ( .A1(n563), .A2(n394), .ZN(n395) );
  NAND2_X1 U453 ( .A1(n395), .A2(n568), .ZN(n396) );
  NAND2_X1 U454 ( .A1(n397), .A2(n396), .ZN(n398) );
  XOR2_X1 U455 ( .A(KEYINPUT48), .B(n398), .Z(n516) );
  XNOR2_X1 U456 ( .A(n399), .B(KEYINPUT54), .ZN(n417) );
  XOR2_X1 U457 ( .A(KEYINPUT5), .B(G57GAT), .Z(n401) );
  XNOR2_X1 U458 ( .A(G1GAT), .B(G120GAT), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n412) );
  XOR2_X1 U460 ( .A(G85GAT), .B(G162GAT), .Z(n403) );
  XNOR2_X1 U461 ( .A(G29GAT), .B(G148GAT), .ZN(n402) );
  XNOR2_X1 U462 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U463 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n405) );
  NAND2_X1 U464 ( .A1(G225GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U465 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U466 ( .A(n407), .B(n406), .Z(n410) );
  XNOR2_X1 U467 ( .A(n408), .B(KEYINPUT4), .ZN(n409) );
  XNOR2_X1 U468 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U469 ( .A(n412), .B(n411), .ZN(n416) );
  XOR2_X1 U470 ( .A(KEYINPUT2), .B(KEYINPUT89), .Z(n414) );
  XNOR2_X1 U471 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U473 ( .A(G141GAT), .B(n415), .ZN(n433) );
  XOR2_X1 U474 ( .A(n416), .B(n433), .Z(n503) );
  INV_X1 U475 ( .A(n503), .ZN(n485) );
  NAND2_X1 U476 ( .A1(n417), .A2(n485), .ZN(n562) );
  XOR2_X1 U477 ( .A(KEYINPUT87), .B(KEYINPUT22), .Z(n419) );
  XNOR2_X1 U478 ( .A(KEYINPUT88), .B(G204GAT), .ZN(n418) );
  XNOR2_X1 U479 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U480 ( .A(n420), .B(KEYINPUT24), .Z(n423) );
  XNOR2_X1 U481 ( .A(G22GAT), .B(n421), .ZN(n422) );
  XNOR2_X1 U482 ( .A(n423), .B(n422), .ZN(n432) );
  XOR2_X1 U483 ( .A(KEYINPUT90), .B(KEYINPUT23), .Z(n425) );
  NAND2_X1 U484 ( .A1(G228GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U485 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U486 ( .A(n426), .B(KEYINPUT91), .Z(n430) );
  XNOR2_X1 U487 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U488 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U489 ( .A(n432), .B(n431), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n434), .B(n433), .ZN(n448) );
  XNOR2_X1 U491 ( .A(n436), .B(n435), .ZN(n437) );
  NAND2_X1 U492 ( .A1(n557), .A2(n531), .ZN(n441) );
  XOR2_X1 U493 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n439) );
  XNOR2_X1 U494 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n462) );
  NAND2_X1 U495 ( .A1(n568), .A2(n563), .ZN(n472) );
  XOR2_X1 U496 ( .A(KEYINPUT16), .B(KEYINPUT82), .Z(n443) );
  NAND2_X1 U497 ( .A1(n572), .A2(n548), .ZN(n442) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n460) );
  XOR2_X1 U499 ( .A(KEYINPUT28), .B(n448), .Z(n496) );
  INV_X1 U500 ( .A(n496), .ZN(n519) );
  XNOR2_X1 U501 ( .A(KEYINPUT27), .B(n506), .ZN(n452) );
  NAND2_X1 U502 ( .A1(n503), .A2(n452), .ZN(n515) );
  NOR2_X1 U503 ( .A1(n519), .A2(n515), .ZN(n444) );
  NAND2_X1 U504 ( .A1(n493), .A2(n444), .ZN(n445) );
  XNOR2_X1 U505 ( .A(n445), .B(KEYINPUT93), .ZN(n458) );
  NOR2_X1 U506 ( .A1(n493), .A2(n491), .ZN(n446) );
  NOR2_X1 U507 ( .A1(n448), .A2(n446), .ZN(n447) );
  XNOR2_X1 U508 ( .A(n447), .B(KEYINPUT25), .ZN(n454) );
  XOR2_X1 U509 ( .A(KEYINPUT95), .B(KEYINPUT26), .Z(n450) );
  NAND2_X1 U510 ( .A1(n493), .A2(n448), .ZN(n449) );
  XNOR2_X1 U511 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U512 ( .A(KEYINPUT94), .B(n451), .ZN(n561) );
  INV_X1 U513 ( .A(n561), .ZN(n535) );
  NAND2_X1 U514 ( .A1(n535), .A2(n452), .ZN(n453) );
  NAND2_X1 U515 ( .A1(n454), .A2(n453), .ZN(n455) );
  XOR2_X1 U516 ( .A(KEYINPUT96), .B(n455), .Z(n456) );
  NOR2_X1 U517 ( .A1(n456), .A2(n503), .ZN(n457) );
  NOR2_X1 U518 ( .A1(n458), .A2(n457), .ZN(n469) );
  INV_X1 U519 ( .A(n469), .ZN(n459) );
  NAND2_X1 U520 ( .A1(n460), .A2(n459), .ZN(n483) );
  NOR2_X1 U521 ( .A1(n472), .A2(n483), .ZN(n467) );
  NAND2_X1 U522 ( .A1(n503), .A2(n467), .ZN(n461) );
  XNOR2_X1 U523 ( .A(n462), .B(n461), .ZN(G1324GAT) );
  NAND2_X1 U524 ( .A1(n467), .A2(n506), .ZN(n463) );
  XNOR2_X1 U525 ( .A(n463), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U526 ( .A(KEYINPUT97), .B(KEYINPUT35), .Z(n465) );
  NAND2_X1 U527 ( .A1(n467), .A2(n517), .ZN(n464) );
  XNOR2_X1 U528 ( .A(n465), .B(n464), .ZN(n466) );
  XOR2_X1 U529 ( .A(G15GAT), .B(n466), .Z(G1326GAT) );
  NAND2_X1 U530 ( .A1(n467), .A2(n519), .ZN(n468) );
  XNOR2_X1 U531 ( .A(n468), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U532 ( .A(G29GAT), .B(KEYINPUT39), .Z(n475) );
  NOR2_X1 U533 ( .A1(n469), .A2(n576), .ZN(n470) );
  NAND2_X1 U534 ( .A1(n470), .A2(n545), .ZN(n471) );
  XOR2_X1 U535 ( .A(KEYINPUT37), .B(n471), .Z(n500) );
  NOR2_X1 U536 ( .A1(n472), .A2(n500), .ZN(n473) );
  XNOR2_X1 U537 ( .A(n473), .B(KEYINPUT38), .ZN(n480) );
  NAND2_X1 U538 ( .A1(n503), .A2(n480), .ZN(n474) );
  XNOR2_X1 U539 ( .A(n475), .B(n474), .ZN(G1328GAT) );
  NAND2_X1 U540 ( .A1(n506), .A2(n480), .ZN(n476) );
  XNOR2_X1 U541 ( .A(G36GAT), .B(n476), .ZN(G1329GAT) );
  XOR2_X1 U542 ( .A(KEYINPUT40), .B(KEYINPUT98), .Z(n478) );
  NAND2_X1 U543 ( .A1(n480), .A2(n517), .ZN(n477) );
  XNOR2_X1 U544 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U545 ( .A(G43GAT), .B(n479), .Z(G1330GAT) );
  NAND2_X1 U546 ( .A1(n480), .A2(n519), .ZN(n481) );
  XNOR2_X1 U547 ( .A(n481), .B(G50GAT), .ZN(G1331GAT) );
  INV_X1 U548 ( .A(n542), .ZN(n554) );
  NAND2_X1 U549 ( .A1(n554), .A2(n537), .ZN(n482) );
  XNOR2_X1 U550 ( .A(n482), .B(KEYINPUT100), .ZN(n501) );
  NOR2_X1 U551 ( .A1(n501), .A2(n483), .ZN(n484) );
  XNOR2_X1 U552 ( .A(KEYINPUT101), .B(n484), .ZN(n495) );
  NOR2_X1 U553 ( .A1(n485), .A2(n495), .ZN(n490) );
  XOR2_X1 U554 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n487) );
  XNOR2_X1 U555 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n486) );
  XNOR2_X1 U556 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U557 ( .A(KEYINPUT99), .B(n488), .ZN(n489) );
  XNOR2_X1 U558 ( .A(n490), .B(n489), .ZN(G1332GAT) );
  NOR2_X1 U559 ( .A1(n491), .A2(n495), .ZN(n492) );
  XOR2_X1 U560 ( .A(G64GAT), .B(n492), .Z(G1333GAT) );
  NOR2_X1 U561 ( .A1(n493), .A2(n495), .ZN(n494) );
  XOR2_X1 U562 ( .A(G71GAT), .B(n494), .Z(G1334GAT) );
  NOR2_X1 U563 ( .A1(n496), .A2(n495), .ZN(n498) );
  XNOR2_X1 U564 ( .A(KEYINPUT104), .B(KEYINPUT43), .ZN(n497) );
  XNOR2_X1 U565 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U566 ( .A(G78GAT), .B(n499), .ZN(G1335GAT) );
  NOR2_X1 U567 ( .A1(n501), .A2(n500), .ZN(n502) );
  XOR2_X1 U568 ( .A(KEYINPUT105), .B(n502), .Z(n511) );
  NAND2_X1 U569 ( .A1(n511), .A2(n503), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n504), .B(KEYINPUT106), .ZN(n505) );
  XNOR2_X1 U571 ( .A(G85GAT), .B(n505), .ZN(G1336GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n508) );
  NAND2_X1 U573 ( .A1(n511), .A2(n506), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U575 ( .A(G92GAT), .B(n509), .ZN(G1337GAT) );
  NAND2_X1 U576 ( .A1(n517), .A2(n511), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n510), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT109), .B(KEYINPUT44), .Z(n513) );
  NAND2_X1 U579 ( .A1(n511), .A2(n519), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U581 ( .A(G106GAT), .B(n514), .ZN(G1339GAT) );
  XOR2_X1 U582 ( .A(G113GAT), .B(KEYINPUT113), .Z(n523) );
  NOR2_X1 U583 ( .A1(n516), .A2(n515), .ZN(n536) );
  NAND2_X1 U584 ( .A1(n536), .A2(n517), .ZN(n518) );
  XOR2_X1 U585 ( .A(KEYINPUT111), .B(n518), .Z(n520) );
  NOR2_X1 U586 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U587 ( .A(KEYINPUT112), .B(n521), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n532), .A2(n563), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(G1340GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n525) );
  NAND2_X1 U591 ( .A1(n554), .A2(n532), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U593 ( .A(G120GAT), .B(n526), .ZN(G1341GAT) );
  XNOR2_X1 U594 ( .A(G127GAT), .B(KEYINPUT115), .ZN(n530) );
  XOR2_X1 U595 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n528) );
  NAND2_X1 U596 ( .A1(n572), .A2(n532), .ZN(n527) );
  XNOR2_X1 U597 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U598 ( .A(n530), .B(n529), .ZN(G1342GAT) );
  XOR2_X1 U599 ( .A(G134GAT), .B(KEYINPUT51), .Z(n534) );
  NAND2_X1 U600 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U601 ( .A(n534), .B(n533), .ZN(G1343GAT) );
  NAND2_X1 U602 ( .A1(n536), .A2(n535), .ZN(n547) );
  NOR2_X1 U603 ( .A1(n537), .A2(n547), .ZN(n539) );
  XNOR2_X1 U604 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(G1344GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT52), .B(KEYINPUT118), .Z(n541) );
  XNOR2_X1 U607 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(n544) );
  NOR2_X1 U609 ( .A1(n542), .A2(n547), .ZN(n543) );
  XOR2_X1 U610 ( .A(n544), .B(n543), .Z(G1345GAT) );
  NOR2_X1 U611 ( .A1(n545), .A2(n547), .ZN(n546) );
  XOR2_X1 U612 ( .A(G155GAT), .B(n546), .Z(G1346GAT) );
  NOR2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U614 ( .A(G162GAT), .B(n549), .Z(G1347GAT) );
  NAND2_X1 U615 ( .A1(n563), .A2(n557), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n552) );
  XNOR2_X1 U618 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U620 ( .A(KEYINPUT56), .B(n553), .Z(n556) );
  NAND2_X1 U621 ( .A1(n557), .A2(n554), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1349GAT) );
  NAND2_X1 U623 ( .A1(n557), .A2(n572), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n560) );
  XNOR2_X1 U626 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n567) );
  XOR2_X1 U628 ( .A(G197GAT), .B(KEYINPUT59), .Z(n565) );
  NOR2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n573) );
  NAND2_X1 U630 ( .A1(n573), .A2(n563), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XOR2_X1 U632 ( .A(n567), .B(n566), .Z(G1352GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n570) );
  INV_X1 U634 ( .A(n573), .ZN(n575) );
  OR2_X1 U635 ( .A1(n575), .A2(n568), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(G204GAT), .B(n571), .ZN(G1353GAT) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U641 ( .A(KEYINPUT62), .B(n577), .Z(n578) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(n578), .ZN(G1355GAT) );
endmodule

