//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 0 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n830, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1029, new_n1030;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n202));
  INV_X1    g001(.A(G197gat), .ZN(new_n203));
  INV_X1    g002(.A(G204gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G197gat), .A2(G204gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT22), .ZN(new_n207));
  NAND2_X1  g006(.A1(G211gat), .A2(G218gat), .ZN(new_n208));
  AOI22_X1  g007(.A1(new_n205), .A2(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G211gat), .ZN(new_n210));
  INV_X1    g009(.A(G218gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n212), .A2(KEYINPUT72), .A3(new_n208), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n209), .A2(new_n213), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n202), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n205), .A2(new_n206), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n208), .A2(new_n207), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AND3_X1   g019(.A1(new_n212), .A2(KEYINPUT72), .A3(new_n208), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(KEYINPUT73), .A3(new_n214), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n217), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G226gat), .ZN(new_n225));
  INV_X1    g024(.A(G233gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(KEYINPUT29), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G190gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT66), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G190gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT28), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT27), .ZN(new_n236));
  INV_X1    g035(.A(G183gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT65), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G183gat), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n236), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n235), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n237), .A2(new_n230), .ZN(new_n244));
  AND2_X1   g043(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n231), .B(new_n233), .C1(new_n245), .C2(new_n242), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n244), .B1(new_n246), .B2(KEYINPUT28), .ZN(new_n247));
  INV_X1    g046(.A(G169gat), .ZN(new_n248));
  INV_X1    g047(.A(G176gat), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT26), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n248), .B(new_n249), .C1(new_n250), .C2(KEYINPUT67), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(KEYINPUT67), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G169gat), .A2(G176gat), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n250), .A2(new_n248), .A3(new_n249), .A4(KEYINPUT67), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n243), .A2(new_n247), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT68), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n243), .A2(new_n247), .A3(new_n259), .A4(new_n256), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NOR3_X1   g062(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n254), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n237), .A2(new_n230), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT24), .B1(new_n237), .B2(new_n230), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT24), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n268), .A2(G183gat), .A3(G190gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n265), .B1(new_n266), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n254), .B(KEYINPUT64), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n272), .B(KEYINPUT25), .C1(new_n263), .C2(new_n264), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n231), .A2(new_n233), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n238), .A2(new_n240), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n274), .A2(new_n275), .B1(new_n267), .B2(new_n269), .ZN(new_n276));
  OAI22_X1  g075(.A1(new_n271), .A2(KEYINPUT25), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n229), .B1(new_n261), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n257), .ZN(new_n279));
  INV_X1    g078(.A(new_n227), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n224), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n224), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n279), .A2(new_n228), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n261), .A2(new_n277), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n283), .B(new_n284), .C1(new_n285), .C2(new_n280), .ZN(new_n286));
  XOR2_X1   g085(.A(G8gat), .B(G36gat), .Z(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(KEYINPUT74), .ZN(new_n288));
  XNOR2_X1  g087(.A(G64gat), .B(G92gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n282), .A2(new_n286), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(KEYINPUT37), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n282), .A2(KEYINPUT37), .A3(new_n286), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT38), .ZN(new_n296));
  OR2_X1    g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n261), .A2(new_n227), .A3(new_n277), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n283), .B1(new_n298), .B2(new_n284), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n278), .A2(new_n281), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT37), .B1(new_n300), .B2(new_n224), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n293), .B(new_n296), .C1(new_n299), .C2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n290), .B1(new_n282), .B2(new_n286), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT5), .ZN(new_n306));
  NAND2_X1  g105(.A1(G225gat), .A2(G233gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT1), .ZN(new_n308));
  INV_X1    g107(.A(G134gat), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n308), .B1(new_n309), .B2(G127gat), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n310), .B1(G127gat), .B2(new_n309), .ZN(new_n311));
  OR2_X1    g110(.A1(G113gat), .A2(G120gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT71), .ZN(new_n313));
  NAND2_X1  g112(.A1(G113gat), .A2(G120gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G113gat), .B(G120gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT71), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n311), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  OR2_X1    g117(.A1(KEYINPUT69), .A2(G134gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(KEYINPUT69), .A2(G134gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(G127gat), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT70), .ZN(new_n322));
  INV_X1    g121(.A(G127gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G134gat), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n312), .A2(new_n308), .A3(new_n314), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n321), .A2(new_n324), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT70), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n318), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  AND2_X1   g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(G141gat), .A2(G148gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G155gat), .B(G162gat), .ZN(new_n334));
  INV_X1    g133(.A(G155gat), .ZN(new_n335));
  INV_X1    g134(.A(G162gat), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT2), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AND3_X1   g136(.A1(new_n333), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT76), .B(KEYINPUT2), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n334), .B1(new_n333), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT3), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  OR2_X1    g140(.A1(G141gat), .A2(G148gat), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT2), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT76), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT2), .ZN(new_n346));
  NAND2_X1  g145(.A1(G141gat), .A2(G148gat), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n342), .A2(new_n344), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  XOR2_X1   g147(.A(G155gat), .B(G162gat), .Z(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n333), .A2(new_n334), .A3(new_n337), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n341), .A2(new_n353), .ZN(new_n354));
  NOR3_X1   g153(.A1(new_n330), .A2(new_n354), .A3(KEYINPUT77), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n351), .B1(new_n350), .B2(new_n352), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n311), .A2(new_n315), .A3(new_n317), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n325), .A2(new_n326), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n322), .B1(new_n321), .B2(new_n324), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n356), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n306), .B(new_n307), .C1(new_n355), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n352), .ZN(new_n366));
  OAI211_X1 g165(.A(KEYINPUT80), .B(KEYINPUT4), .C1(new_n363), .C2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n329), .A2(new_n326), .A3(new_n325), .ZN(new_n368));
  INV_X1    g167(.A(new_n366), .ZN(new_n369));
  XOR2_X1   g168(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n370));
  NAND4_X1  g169(.A1(new_n368), .A2(new_n369), .A3(new_n360), .A4(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n368), .A2(new_n369), .A3(new_n360), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT80), .B1(new_n373), .B2(KEYINPUT4), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT81), .B1(new_n365), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT80), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n363), .A2(new_n366), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT4), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(new_n371), .A3(new_n367), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT81), .ZN(new_n382));
  INV_X1    g181(.A(new_n307), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT77), .B1(new_n330), .B2(new_n354), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n359), .A2(new_n356), .A3(new_n363), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n381), .A2(new_n382), .A3(new_n386), .A4(new_n306), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n376), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(KEYINPUT0), .ZN(new_n390));
  XNOR2_X1  g189(.A(G57gat), .B(G85gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n390), .B(new_n391), .Z(new_n392));
  AOI21_X1  g191(.A(new_n369), .B1(new_n368), .B2(new_n360), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n383), .B1(new_n378), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT5), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT79), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n373), .A2(new_n370), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n368), .A2(new_n369), .A3(KEYINPUT4), .A4(new_n360), .ZN(new_n398));
  AND2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n386), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT79), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n394), .A2(new_n401), .A3(KEYINPUT5), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n396), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n388), .A2(new_n392), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT82), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n388), .A2(new_n403), .ZN(new_n407));
  INV_X1    g206(.A(new_n392), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT6), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n392), .B1(new_n388), .B2(new_n403), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT6), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n388), .A2(KEYINPUT82), .A3(new_n403), .A4(new_n392), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n297), .B(new_n305), .C1(new_n410), .C2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(G22gat), .ZN(new_n416));
  AND2_X1   g215(.A1(G228gat), .A2(G233gat), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT29), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n353), .A2(new_n419), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n224), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n212), .A2(new_n208), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n220), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n419), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n220), .A2(new_n422), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n351), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n426), .A2(new_n366), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n418), .B1(new_n421), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT29), .B1(new_n222), .B2(new_n214), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n351), .B1(new_n429), .B2(KEYINPUT83), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT83), .ZN(new_n431));
  AOI211_X1 g230(.A(new_n431), .B(KEYINPUT29), .C1(new_n222), .C2(new_n214), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n366), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n418), .B1(new_n224), .B2(new_n420), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT84), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n435), .B1(new_n433), .B2(new_n434), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n416), .B(new_n428), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT85), .ZN(new_n439));
  XNOR2_X1  g238(.A(G78gat), .B(G106gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT31), .B(G50gat), .ZN(new_n441));
  XOR2_X1   g240(.A(new_n440), .B(new_n441), .Z(new_n442));
  NAND2_X1  g241(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n428), .B1(new_n436), .B2(new_n437), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(G22gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n438), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT85), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n445), .A2(new_n448), .A3(new_n438), .A4(new_n442), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT75), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT30), .B1(new_n303), .B2(new_n451), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n452), .A2(new_n291), .ZN(new_n453));
  OR3_X1    g252(.A1(new_n303), .A2(new_n451), .A3(KEYINPUT30), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n411), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n384), .A2(new_n385), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n307), .B1(new_n381), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT39), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n392), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT40), .ZN(new_n461));
  OR2_X1    g260(.A1(new_n378), .A2(new_n393), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT39), .B1(new_n462), .B2(new_n383), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  NOR3_X1   g263(.A1(new_n460), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n464), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n408), .B1(new_n457), .B2(new_n458), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT40), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n450), .B1(new_n455), .B2(new_n469), .ZN(new_n470));
  XOR2_X1   g269(.A(G15gat), .B(G43gat), .Z(new_n471));
  XNOR2_X1  g270(.A(G71gat), .B(G99gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n471), .B(new_n472), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n261), .A2(new_n363), .A3(new_n277), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n363), .B1(new_n261), .B2(new_n277), .ZN(new_n475));
  INV_X1    g274(.A(G227gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n476), .A2(new_n226), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  NOR3_X1   g277(.A1(new_n474), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n473), .B1(new_n479), .B2(KEYINPUT33), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n478), .B1(new_n474), .B2(new_n475), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT34), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT34), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n483), .B(new_n478), .C1(new_n474), .C2(new_n475), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n473), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n285), .A2(new_n330), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n261), .A2(new_n363), .A3(new_n277), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n477), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT33), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n486), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n487), .A2(new_n488), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n483), .B1(new_n492), .B2(new_n478), .ZN(new_n493));
  INV_X1    g292(.A(new_n484), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n485), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n489), .A2(KEYINPUT32), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n497), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n485), .A2(new_n495), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(KEYINPUT36), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT36), .ZN(new_n502));
  INV_X1    g301(.A(new_n500), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n499), .B1(new_n485), .B2(new_n495), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n415), .A2(new_n470), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  AOI22_X1  g305(.A1(KEYINPUT79), .A2(new_n395), .B1(new_n386), .B2(new_n399), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n376), .A2(new_n387), .B1(new_n507), .B2(new_n402), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT82), .B1(new_n508), .B2(new_n392), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n412), .B1(new_n509), .B2(new_n411), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n413), .A2(new_n412), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(new_n409), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n454), .A2(new_n291), .A3(new_n452), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n510), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n450), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n506), .A2(new_n516), .ZN(new_n517));
  NOR3_X1   g316(.A1(new_n410), .A2(new_n414), .A3(new_n513), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n498), .A2(new_n449), .A3(new_n447), .A4(new_n500), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT86), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n518), .A2(new_n520), .A3(new_n521), .A4(KEYINPUT35), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n519), .A2(KEYINPUT35), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT35), .ZN(new_n524));
  INV_X1    g323(.A(new_n449), .ZN(new_n525));
  AOI22_X1  g324(.A1(new_n439), .A2(new_n442), .B1(new_n445), .B2(new_n438), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n527), .A2(new_n521), .A3(new_n500), .A4(new_n498), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n523), .B(new_n524), .C1(new_n515), .C2(new_n528), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n517), .A2(KEYINPUT87), .A3(new_n522), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n505), .A2(new_n501), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n302), .B(new_n304), .C1(new_n295), .C2(new_n296), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n532), .B1(new_n510), .B2(new_n512), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n461), .B1(new_n460), .B2(new_n464), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n466), .A2(KEYINPUT40), .A3(new_n467), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n513), .A2(new_n409), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(new_n527), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n531), .B1(new_n533), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n518), .A2(new_n527), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n529), .B(new_n522), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT87), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT15), .ZN(new_n543));
  XOR2_X1   g342(.A(KEYINPUT90), .B(G43gat), .Z(new_n544));
  NOR2_X1   g343(.A1(new_n544), .A2(G50gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT91), .B(G50gat), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n546), .A2(G43gat), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n543), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G43gat), .B(G50gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT15), .ZN(new_n550));
  OR3_X1    g349(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G29gat), .A2(G36gat), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n550), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n548), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT88), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g357(.A(KEYINPUT88), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n558), .A2(new_n551), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n550), .B1(new_n560), .B2(new_n554), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n561), .A2(KEYINPUT89), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(KEYINPUT89), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n556), .B(KEYINPUT17), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G15gat), .B(G22gat), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT16), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n565), .B1(new_n566), .B2(G1gat), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n567), .B1(G1gat), .B2(new_n565), .ZN(new_n568));
  INV_X1    g367(.A(G8gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n561), .A2(KEYINPUT89), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n561), .A2(KEYINPUT89), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n571), .A2(new_n572), .B1(new_n548), .B2(new_n555), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT92), .B(KEYINPUT17), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n564), .B(new_n570), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n570), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n556), .B1(new_n562), .B2(new_n563), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT93), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n574), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n581), .A2(KEYINPUT93), .A3(new_n564), .A4(new_n570), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G229gat), .A2(G233gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT18), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n585), .A2(KEYINPUT94), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT94), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n579), .A2(new_n582), .B1(G229gat), .B2(G233gat), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n588), .B1(new_n589), .B2(KEYINPUT18), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n577), .B(new_n570), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n584), .B(KEYINPUT13), .Z(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n594), .B1(new_n589), .B2(KEYINPUT18), .ZN(new_n595));
  XNOR2_X1  g394(.A(G113gat), .B(G141gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(G197gat), .ZN(new_n597));
  XOR2_X1   g396(.A(KEYINPUT11), .B(G169gat), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n599), .B(KEYINPUT12), .Z(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n587), .A2(new_n590), .A3(new_n595), .A4(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n583), .A2(KEYINPUT18), .A3(new_n584), .ZN(new_n603));
  INV_X1    g402(.A(new_n594), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n589), .A2(KEYINPUT18), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n600), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT95), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n602), .A2(new_n607), .A3(KEYINPUT95), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(G64gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(G57gat), .ZN(new_n614));
  INV_X1    g413(.A(G57gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(G64gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT9), .ZN(new_n618));
  OR2_X1    g417(.A1(G71gat), .A2(G78gat), .ZN(new_n619));
  NAND2_X1  g418(.A1(G71gat), .A2(G78gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT96), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n618), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT9), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n625), .B1(new_n614), .B2(new_n616), .ZN(new_n626));
  OAI21_X1  g425(.A(KEYINPUT96), .B1(new_n626), .B2(new_n621), .ZN(new_n627));
  XOR2_X1   g426(.A(KEYINPUT97), .B(G57gat), .Z(new_n628));
  OAI21_X1  g427(.A(new_n614), .B1(new_n628), .B2(new_n613), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n620), .B1(new_n619), .B2(new_n625), .ZN(new_n630));
  AOI22_X1  g429(.A1(new_n624), .A2(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n631), .A2(KEYINPUT21), .ZN(new_n632));
  NAND2_X1  g431(.A1(G231gat), .A2(G233gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G127gat), .B(G155gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT98), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n634), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(G183gat), .B(G211gat), .Z(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n637), .B(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n576), .B1(KEYINPUT21), .B2(new_n631), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n640), .B(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT99), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT100), .B(G92gat), .ZN(new_n646));
  INV_X1    g445(.A(G85gat), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G85gat), .A2(G92gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT7), .ZN(new_n650));
  INV_X1    g449(.A(G99gat), .ZN(new_n651));
  INV_X1    g450(.A(G106gat), .ZN(new_n652));
  OAI21_X1  g451(.A(KEYINPUT8), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n648), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g453(.A(G99gat), .B(G106gat), .Z(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n655), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n657), .A2(new_n648), .A3(new_n650), .A4(new_n653), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n581), .A2(new_n564), .A3(new_n659), .ZN(new_n660));
  AND3_X1   g459(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n661));
  INV_X1    g460(.A(new_n659), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n661), .B1(new_n577), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT101), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT101), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n660), .A2(new_n666), .A3(new_n663), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(G190gat), .B(G218gat), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n645), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n669), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n665), .A2(new_n667), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(G134gat), .B(G162gat), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n674), .B(new_n675), .Z(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n670), .A2(new_n672), .A3(new_n676), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n631), .A2(new_n658), .A3(new_n656), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT10), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n624), .A2(new_n627), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n629), .A2(new_n630), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n659), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n687), .A2(new_n681), .A3(KEYINPUT102), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT102), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n662), .A2(new_n689), .A3(new_n631), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n683), .B1(new_n691), .B2(new_n682), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(KEYINPUT103), .ZN(new_n693));
  NAND2_X1  g492(.A1(G230gat), .A2(G233gat), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT10), .B1(new_n688), .B2(new_n690), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n695), .B1(new_n696), .B2(new_n683), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n693), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n694), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n688), .A2(new_n699), .A3(new_n690), .ZN(new_n700));
  XNOR2_X1  g499(.A(G120gat), .B(G148gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(G176gat), .B(G204gat), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n701), .B(new_n702), .Z(new_n703));
  AND2_X1   g502(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n698), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n700), .B1(new_n692), .B2(new_n699), .ZN(new_n706));
  INV_X1    g505(.A(new_n703), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n644), .A2(new_n680), .A3(new_n709), .ZN(new_n710));
  AND4_X1   g509(.A1(new_n530), .A2(new_n542), .A3(new_n612), .A4(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n410), .A2(new_n414), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g514(.A(new_n569), .B1(new_n711), .B2(new_n513), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n542), .A2(new_n530), .A3(new_n612), .A4(new_n710), .ZN(new_n717));
  XNOR2_X1  g516(.A(KEYINPUT16), .B(G8gat), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n717), .A2(new_n514), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(KEYINPUT42), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n542), .A2(new_n530), .A3(new_n612), .ZN(new_n722));
  INV_X1    g521(.A(new_n718), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n722), .A2(new_n513), .A3(new_n710), .A4(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT42), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n720), .A2(new_n721), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G8gat), .B1(new_n717), .B2(new_n514), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n725), .B1(new_n724), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n719), .A2(KEYINPUT42), .ZN(new_n730));
  OAI21_X1  g529(.A(KEYINPUT104), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n727), .A2(new_n731), .ZN(G1325gat));
  OAI21_X1  g531(.A(G15gat), .B1(new_n717), .B2(new_n531), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n503), .A2(new_n504), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n735), .A2(G15gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n733), .B1(new_n717), .B2(new_n736), .ZN(G1326gat));
  NOR2_X1   g536(.A1(new_n717), .A2(new_n527), .ZN(new_n738));
  XOR2_X1   g537(.A(KEYINPUT43), .B(G22gat), .Z(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(G1327gat));
  INV_X1    g539(.A(KEYINPUT45), .ZN(new_n741));
  INV_X1    g540(.A(new_n709), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n644), .A2(new_n680), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT105), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n722), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n712), .A2(G29gat), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n741), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n722), .A2(KEYINPUT45), .A3(new_n744), .A4(new_n746), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT106), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(new_n518), .B2(new_n527), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n515), .A2(KEYINPUT106), .A3(new_n450), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n506), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n753), .A2(new_n522), .A3(new_n529), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n680), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n542), .A2(new_n530), .A3(KEYINPUT44), .A4(new_n680), .ZN(new_n758));
  INV_X1    g557(.A(new_n644), .ZN(new_n759));
  INV_X1    g558(.A(new_n608), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n759), .A2(new_n760), .A3(new_n709), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n757), .A2(new_n758), .A3(new_n713), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(KEYINPUT107), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G29gat), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n762), .A2(KEYINPUT107), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n748), .B(new_n749), .C1(new_n764), .C2(new_n765), .ZN(G1328gat));
  AOI21_X1  g565(.A(G36gat), .B1(KEYINPUT108), .B2(KEYINPUT46), .ZN(new_n767));
  AND4_X1   g566(.A1(new_n513), .A2(new_n722), .A3(new_n744), .A4(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n757), .A2(new_n758), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n771), .A2(new_n513), .A3(new_n761), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G36gat), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n768), .A2(new_n769), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n770), .A2(new_n773), .A3(new_n774), .ZN(G1329gat));
  INV_X1    g574(.A(KEYINPUT47), .ZN(new_n776));
  INV_X1    g575(.A(new_n531), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n757), .A2(new_n758), .A3(new_n777), .A4(new_n761), .ZN(new_n778));
  INV_X1    g577(.A(new_n544), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n734), .A2(new_n544), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n745), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n776), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n778), .A2(new_n779), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n784), .B(KEYINPUT47), .C1(new_n745), .C2(new_n781), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(G1330gat));
  OAI21_X1  g585(.A(new_n546), .B1(new_n745), .B2(new_n527), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n527), .A2(new_n546), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n757), .A2(new_n758), .A3(new_n761), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT48), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT48), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n787), .A2(new_n792), .A3(new_n789), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(G1331gat));
  NOR2_X1   g593(.A1(new_n644), .A2(new_n680), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n795), .A2(new_n760), .A3(new_n709), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT109), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT109), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n795), .A2(new_n798), .A3(new_n760), .A4(new_n709), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n754), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT110), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n754), .A2(new_n800), .A3(KEYINPUT110), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n713), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(new_n628), .ZN(G1332gat));
  INV_X1    g606(.A(KEYINPUT49), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n613), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT111), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n514), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n810), .B1(new_n805), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n803), .A2(new_n804), .ZN(new_n813));
  INV_X1    g612(.A(new_n811), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n813), .A2(KEYINPUT111), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n809), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n805), .A2(new_n810), .A3(new_n811), .ZN(new_n817));
  OAI21_X1  g616(.A(KEYINPUT111), .B1(new_n813), .B2(new_n814), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n817), .A2(new_n808), .A3(new_n818), .A4(new_n613), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n816), .A2(new_n819), .ZN(G1333gat));
  INV_X1    g619(.A(KEYINPUT50), .ZN(new_n821));
  INV_X1    g620(.A(G71gat), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n822), .B1(new_n805), .B2(new_n777), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n734), .A2(new_n822), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n813), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n821), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(G71gat), .B1(new_n813), .B2(new_n531), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n827), .B(KEYINPUT50), .C1(new_n813), .C2(new_n824), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(G1334gat));
  NAND2_X1  g628(.A1(new_n805), .A2(new_n450), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g630(.A1(new_n759), .A2(new_n608), .A3(new_n742), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n771), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(G85gat), .B1(new_n833), .B2(new_n712), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n759), .A2(new_n608), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n506), .A2(new_n751), .A3(new_n752), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n529), .A2(new_n522), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n680), .B(new_n835), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT51), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n754), .A2(KEYINPUT51), .A3(new_n680), .A4(new_n835), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n713), .A2(new_n647), .A3(new_n709), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n834), .B1(new_n843), .B2(new_n844), .ZN(G1336gat));
  INV_X1    g644(.A(KEYINPUT112), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n840), .A2(new_n846), .A3(new_n841), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n838), .A2(KEYINPUT112), .A3(new_n839), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n514), .A2(new_n742), .A3(G92gat), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n757), .A2(new_n758), .A3(new_n513), .A4(new_n832), .ZN(new_n851));
  INV_X1    g650(.A(new_n646), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT52), .ZN(new_n855));
  AOI21_X1  g654(.A(KEYINPUT52), .B1(new_n842), .B2(new_n849), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n853), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n857), .ZN(G1337gat));
  OAI21_X1  g657(.A(G99gat), .B1(new_n833), .B2(new_n531), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n734), .A2(new_n651), .A3(new_n709), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT113), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n859), .B1(new_n843), .B2(new_n861), .ZN(G1338gat));
  NOR3_X1   g661(.A1(new_n527), .A2(new_n742), .A3(G106gat), .ZN(new_n863));
  XOR2_X1   g662(.A(new_n863), .B(KEYINPUT114), .Z(new_n864));
  NAND3_X1  g663(.A1(new_n847), .A2(new_n848), .A3(new_n864), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n757), .A2(new_n758), .A3(new_n450), .A4(new_n832), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(G106gat), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT53), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT53), .B1(new_n842), .B2(new_n863), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n867), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(G1339gat));
  INV_X1    g671(.A(new_n705), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n874), .B1(new_n692), .B2(new_n699), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n697), .A2(new_n694), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n696), .A2(new_n695), .A3(new_n683), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n874), .B(new_n694), .C1(new_n696), .C2(new_n683), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT115), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n880), .A3(new_n707), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n880), .B1(new_n879), .B2(new_n707), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n878), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT55), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n873), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n698), .B2(new_n875), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n879), .A2(new_n707), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT115), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n881), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n887), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n891), .B1(new_n887), .B2(new_n890), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n886), .B(new_n608), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n591), .A2(new_n593), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n895), .B1(new_n583), .B2(new_n584), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n599), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n602), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n709), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n680), .B1(new_n894), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n680), .A2(new_n898), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n886), .B1(new_n892), .B2(new_n893), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n644), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n795), .A2(new_n760), .A3(new_n742), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n519), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n712), .A2(new_n513), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n909), .A2(G113gat), .A3(new_n612), .ZN(new_n910));
  AOI21_X1  g709(.A(G113gat), .B1(new_n909), .B2(new_n608), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n910), .A2(new_n911), .ZN(G1340gat));
  NAND2_X1  g711(.A1(new_n909), .A2(new_n709), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(G120gat), .ZN(G1341gat));
  NOR2_X1   g713(.A1(new_n908), .A2(new_n644), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(new_n323), .ZN(G1342gat));
  NAND2_X1  g715(.A1(new_n909), .A2(new_n680), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n319), .A2(new_n320), .ZN(new_n918));
  OR3_X1    g717(.A1(new_n917), .A2(KEYINPUT56), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(G134gat), .ZN(new_n920));
  OAI21_X1  g719(.A(KEYINPUT56), .B1(new_n917), .B2(new_n918), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(G1343gat));
  INV_X1    g721(.A(new_n905), .ZN(new_n923));
  AOI22_X1  g722(.A1(new_n889), .A2(new_n881), .B1(new_n698), .B2(new_n875), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n705), .B1(new_n924), .B2(KEYINPUT55), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n887), .A2(new_n890), .A3(new_n891), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n887), .A2(new_n890), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT116), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n925), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  AOI22_X1  g728(.A1(new_n929), .A2(new_n612), .B1(new_n709), .B2(new_n898), .ZN(new_n930));
  OAI22_X1  g729(.A1(new_n930), .A2(new_n680), .B1(new_n902), .B2(new_n901), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n923), .B1(new_n931), .B2(new_n644), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT57), .B1(new_n932), .B2(new_n527), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n907), .A2(new_n531), .ZN(new_n934));
  XOR2_X1   g733(.A(new_n934), .B(KEYINPUT117), .Z(new_n935));
  AOI21_X1  g734(.A(new_n527), .B1(new_n904), .B2(new_n905), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT57), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n933), .A2(new_n938), .A3(new_n612), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(G141gat), .ZN(new_n940));
  AOI211_X1 g739(.A(new_n527), .B(new_n777), .C1(new_n904), .C2(new_n905), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n907), .ZN(new_n942));
  INV_X1    g741(.A(new_n612), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n943), .A2(G141gat), .ZN(new_n944));
  XOR2_X1   g743(.A(new_n944), .B(KEYINPUT118), .Z(new_n945));
  NOR2_X1   g744(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  XNOR2_X1  g746(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n940), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT58), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n933), .A2(new_n938), .A3(new_n608), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n946), .B1(new_n951), .B2(G141gat), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n949), .B1(new_n950), .B2(new_n952), .ZN(G1344gat));
  OR3_X1    g752(.A1(new_n942), .A2(G148gat), .A3(new_n742), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT59), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n931), .A2(new_n644), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n710), .A2(new_n943), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n527), .A2(KEYINPUT57), .ZN(new_n959));
  INV_X1    g758(.A(new_n936), .ZN(new_n960));
  AOI22_X1  g759(.A1(new_n958), .A2(new_n959), .B1(new_n960), .B2(KEYINPUT57), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n935), .A2(new_n742), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n955), .B1(new_n963), .B2(G148gat), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n955), .A2(G148gat), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n933), .A2(new_n938), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n965), .B1(new_n966), .B2(new_n709), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n954), .B1(new_n964), .B2(new_n967), .ZN(G1345gat));
  AOI21_X1  g767(.A(new_n335), .B1(new_n966), .B2(new_n759), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n942), .A2(G155gat), .A3(new_n644), .ZN(new_n970));
  OR2_X1    g769(.A1(new_n969), .A2(new_n970), .ZN(G1346gat));
  NAND2_X1  g770(.A1(new_n680), .A2(new_n336), .ZN(new_n972));
  OR3_X1    g771(.A1(new_n942), .A2(KEYINPUT120), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g772(.A(KEYINPUT120), .B1(new_n942), .B2(new_n972), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n966), .A2(new_n680), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n975), .B1(new_n976), .B2(new_n336), .ZN(G1347gat));
  NOR2_X1   g776(.A1(new_n713), .A2(new_n514), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n906), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n979), .A2(new_n248), .A3(new_n608), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT121), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n248), .B1(new_n979), .B2(new_n612), .ZN(new_n982));
  OR2_X1    g781(.A1(new_n982), .A2(KEYINPUT122), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(KEYINPUT122), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n981), .A2(new_n983), .A3(new_n984), .ZN(G1348gat));
  NAND2_X1  g784(.A1(new_n979), .A2(new_n709), .ZN(new_n986));
  XNOR2_X1  g785(.A(new_n986), .B(G176gat), .ZN(G1349gat));
  INV_X1    g786(.A(KEYINPUT125), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n904), .A2(new_n905), .ZN(new_n989));
  NAND4_X1  g788(.A1(new_n989), .A2(new_n520), .A3(new_n759), .A4(new_n978), .ZN(new_n990));
  INV_X1    g789(.A(new_n275), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n991), .A2(KEYINPUT123), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n245), .A2(new_n242), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n994), .B1(new_n275), .B2(KEYINPUT123), .ZN(new_n995));
  INV_X1    g794(.A(new_n995), .ZN(new_n996));
  NAND4_X1  g795(.A1(new_n906), .A2(new_n759), .A3(new_n978), .A4(new_n996), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n988), .B1(new_n993), .B2(new_n997), .ZN(new_n998));
  NOR3_X1   g797(.A1(new_n998), .A2(KEYINPUT124), .A3(KEYINPUT60), .ZN(new_n999));
  OR2_X1    g798(.A1(new_n998), .A2(KEYINPUT124), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT60), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n993), .A2(new_n997), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n1001), .B1(new_n1002), .B2(KEYINPUT124), .ZN(new_n1003));
  AOI21_X1  g802(.A(new_n999), .B1(new_n1000), .B2(new_n1003), .ZN(G1350gat));
  AOI21_X1  g803(.A(new_n230), .B1(new_n979), .B2(new_n680), .ZN(new_n1005));
  OR2_X1    g804(.A1(new_n1005), .A2(KEYINPUT61), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1005), .A2(KEYINPUT61), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n979), .A2(new_n274), .A3(new_n680), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(G1351gat));
  AND2_X1   g808(.A1(new_n941), .A2(new_n978), .ZN(new_n1010));
  AOI21_X1  g809(.A(G197gat), .B1(new_n1010), .B2(new_n608), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n978), .A2(new_n531), .ZN(new_n1012));
  XNOR2_X1  g811(.A(new_n1012), .B(KEYINPUT126), .ZN(new_n1013));
  AND2_X1   g812(.A1(new_n961), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g813(.A1(new_n943), .A2(new_n203), .ZN(new_n1015));
  AOI21_X1  g814(.A(new_n1011), .B1(new_n1014), .B2(new_n1015), .ZN(G1352gat));
  NAND4_X1  g815(.A1(new_n941), .A2(new_n204), .A3(new_n709), .A4(new_n978), .ZN(new_n1017));
  XOR2_X1   g816(.A(new_n1017), .B(KEYINPUT62), .Z(new_n1018));
  AND3_X1   g817(.A1(new_n961), .A2(new_n709), .A3(new_n1013), .ZN(new_n1019));
  OAI21_X1  g818(.A(new_n1018), .B1(new_n1019), .B2(new_n204), .ZN(G1353gat));
  NAND3_X1  g819(.A1(new_n1010), .A2(new_n210), .A3(new_n759), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n958), .A2(new_n959), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n960), .A2(KEYINPUT57), .ZN(new_n1023));
  NOR2_X1   g822(.A1(new_n1012), .A2(new_n644), .ZN(new_n1024));
  NAND3_X1  g823(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  AND3_X1   g824(.A1(new_n1025), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1026));
  AOI21_X1  g825(.A(KEYINPUT63), .B1(new_n1025), .B2(G211gat), .ZN(new_n1027));
  OAI21_X1  g826(.A(new_n1021), .B1(new_n1026), .B2(new_n1027), .ZN(G1354gat));
  NAND3_X1  g827(.A1(new_n1010), .A2(new_n211), .A3(new_n680), .ZN(new_n1029));
  AND3_X1   g828(.A1(new_n961), .A2(new_n680), .A3(new_n1013), .ZN(new_n1030));
  OAI21_X1  g829(.A(new_n1029), .B1(new_n1030), .B2(new_n211), .ZN(G1355gat));
endmodule


