//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1206,
    new_n1207, new_n1208, new_n1210, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  AND2_X1   g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G20), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n207), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n210), .B1(new_n212), .B2(new_n213), .C1(KEYINPUT1), .C2(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(KEYINPUT1), .B2(new_n220), .ZN(G361));
  XNOR2_X1  g0022(.A(G238), .B(G244), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(G232), .ZN(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT2), .B(G226), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(G264), .B(G270), .Z(new_n227));
  XNOR2_X1  g0027(.A(G250), .B(G257), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n226), .B(new_n229), .ZN(G358));
  XOR2_X1   g0030(.A(G87), .B(G97), .Z(new_n231));
  XNOR2_X1  g0031(.A(G107), .B(G116), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n201), .A2(G68), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n203), .A2(G50), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G58), .B(G77), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n233), .B(new_n238), .ZN(G351));
  NAND2_X1  g0039(.A1(G33), .A2(G41), .ZN(new_n240));
  NAND3_X1  g0040(.A1(new_n240), .A2(G1), .A3(G13), .ZN(new_n241));
  INV_X1    g0041(.A(G1), .ZN(new_n242));
  OAI21_X1  g0042(.A(new_n242), .B1(G41), .B2(G45), .ZN(new_n243));
  AND3_X1   g0043(.A1(new_n241), .A2(G226), .A3(new_n243), .ZN(new_n244));
  AND2_X1   g0044(.A1(G33), .A2(G41), .ZN(new_n245));
  NAND2_X1  g0045(.A1(G1), .A2(G13), .ZN(new_n246));
  OAI21_X1  g0046(.A(G274), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g0047(.A(KEYINPUT64), .B1(new_n247), .B2(new_n243), .ZN(new_n248));
  INV_X1    g0048(.A(G274), .ZN(new_n249));
  AOI21_X1  g0049(.A(new_n249), .B1(new_n211), .B2(new_n240), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT64), .ZN(new_n251));
  INV_X1    g0051(.A(new_n243), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n244), .B1(new_n248), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  AND2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  OAI211_X1 g0057(.A(G222), .B(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  OAI211_X1 g0058(.A(G223), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n259));
  OR2_X1    g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n260), .A2(G77), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n258), .A2(new_n259), .A3(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n245), .A2(new_n246), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AND3_X1   g0065(.A1(new_n254), .A2(KEYINPUT65), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(KEYINPUT65), .B1(new_n254), .B2(new_n265), .ZN(new_n267));
  OAI21_X1  g0067(.A(G190), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT9), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n246), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT66), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT66), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n270), .A2(new_n273), .A3(new_n246), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G13), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(G1), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G20), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n201), .B1(new_n242), .B2(G20), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n275), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT8), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(new_n202), .B2(KEYINPUT67), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT67), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(KEYINPUT8), .A3(G58), .ZN(new_n284));
  INV_X1    g0084(.A(G20), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n282), .A2(new_n284), .A3(new_n285), .A4(G33), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n275), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n280), .B1(new_n289), .B2(KEYINPUT68), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n286), .ZN(new_n291));
  AND3_X1   g0091(.A1(new_n270), .A2(new_n273), .A3(new_n246), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n273), .B1(new_n270), .B2(new_n246), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n291), .A2(KEYINPUT68), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n278), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n201), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n269), .B1(new_n290), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n291), .A2(new_n294), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT68), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n294), .A2(new_n296), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n300), .A2(new_n301), .B1(new_n302), .B2(new_n279), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n295), .A2(new_n297), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n303), .A2(new_n304), .A3(KEYINPUT9), .ZN(new_n305));
  AND3_X1   g0105(.A1(new_n268), .A2(new_n299), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(KEYINPUT69), .A2(KEYINPUT70), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT10), .ZN(new_n308));
  INV_X1    g0108(.A(G200), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n266), .A2(new_n267), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT10), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT69), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n308), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n306), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n268), .A2(new_n299), .A3(new_n305), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n310), .B1(new_n315), .B2(KEYINPUT70), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n314), .B1(new_n316), .B2(new_n311), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n266), .A2(new_n267), .ZN(new_n318));
  INV_X1    g0118(.A(G169), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n303), .A2(new_n304), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n320), .B(new_n321), .C1(G179), .C2(new_n318), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(G20), .A2(G77), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT15), .B(G87), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n285), .A2(G33), .ZN(new_n326));
  INV_X1    g0126(.A(new_n287), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT8), .B(G58), .ZN(new_n328));
  OAI221_X1 g0128(.A(new_n324), .B1(new_n325), .B2(new_n326), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G77), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n329), .A2(new_n294), .B1(new_n330), .B2(new_n296), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n242), .A2(G20), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n302), .A2(G77), .A3(new_n332), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n260), .A2(new_n261), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(G232), .A3(new_n255), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(G238), .A3(G1698), .ZN(new_n337));
  INV_X1    g0137(.A(G107), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n336), .B(new_n337), .C1(new_n338), .C2(new_n335), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n264), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n248), .A2(new_n253), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n264), .A2(new_n252), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G244), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n340), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n334), .B1(new_n344), .B2(new_n319), .ZN(new_n345));
  OR2_X1    g0145(.A1(new_n344), .A2(G179), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n344), .A2(G200), .ZN(new_n348));
  INV_X1    g0148(.A(G190), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n334), .B1(new_n344), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n347), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n323), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n296), .A2(KEYINPUT76), .A3(new_n203), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT12), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT76), .B1(new_n296), .B2(new_n203), .ZN(new_n355));
  XOR2_X1   g0155(.A(new_n354), .B(new_n355), .Z(new_n356));
  AOI22_X1  g0156(.A1(new_n287), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n330), .B2(new_n326), .ZN(new_n358));
  AND3_X1   g0158(.A1(new_n294), .A2(new_n358), .A3(KEYINPUT11), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT11), .B1(new_n294), .B2(new_n358), .ZN(new_n360));
  OR3_X1    g0160(.A1(new_n359), .A2(new_n360), .A3(KEYINPUT74), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT74), .B1(new_n359), .B2(new_n360), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n275), .A2(G68), .A3(new_n278), .A4(new_n332), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT75), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n363), .B(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n356), .A2(new_n361), .A3(new_n362), .A4(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT72), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n341), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n248), .A2(KEYINPUT72), .A3(new_n253), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G232), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(G1698), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(G226), .B2(G1698), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n256), .A2(new_n257), .ZN(new_n374));
  INV_X1    g0174(.A(G33), .ZN(new_n375));
  INV_X1    g0175(.A(G97), .ZN(new_n376));
  OAI22_X1  g0176(.A1(new_n373), .A2(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n377), .A2(KEYINPUT71), .A3(new_n264), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n264), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT71), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n379), .A2(new_n380), .B1(G238), .B2(new_n342), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n370), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n349), .B1(new_n382), .B2(KEYINPUT13), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT13), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n370), .A2(new_n381), .A3(new_n384), .A4(new_n378), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n366), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n369), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT72), .B1(new_n248), .B2(new_n253), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(G226), .A2(G1698), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n371), .B2(G1698), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n391), .A2(new_n335), .B1(G33), .B2(G97), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n380), .B1(new_n392), .B2(new_n241), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n342), .A2(G238), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(new_n378), .A3(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT13), .B1(new_n389), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(new_n385), .A3(KEYINPUT73), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT73), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n382), .A2(new_n398), .A3(KEYINPUT13), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(G200), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n386), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n397), .A2(G169), .A3(new_n399), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT14), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n396), .A2(new_n385), .A3(G179), .ZN(new_n405));
  XNOR2_X1  g0205(.A(KEYINPUT77), .B(KEYINPUT14), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n397), .A2(G169), .A3(new_n399), .A4(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n404), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n402), .B1(new_n408), .B2(new_n366), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n282), .A2(new_n284), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n332), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n413), .A2(new_n302), .B1(new_n296), .B2(new_n410), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n202), .A2(new_n203), .ZN(new_n416));
  NOR2_X1   g0216(.A1(G58), .A2(G68), .ZN(new_n417));
  OAI21_X1  g0217(.A(G20), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n287), .A2(G159), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT7), .ZN(new_n422));
  NOR4_X1   g0222(.A1(new_n256), .A2(new_n257), .A3(new_n422), .A4(G20), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n260), .A2(KEYINPUT78), .A3(new_n261), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT78), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n256), .B2(new_n257), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n424), .A2(new_n426), .A3(new_n285), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n423), .B1(new_n427), .B2(new_n422), .ZN(new_n428));
  OAI211_X1 g0228(.A(KEYINPUT16), .B(new_n421), .C1(new_n428), .C2(new_n203), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT16), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n422), .B1(new_n335), .B2(G20), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n374), .A2(KEYINPUT7), .A3(new_n285), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n203), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n430), .B1(new_n433), .B2(new_n420), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n429), .A2(new_n294), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT79), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT7), .B1(new_n374), .B2(new_n285), .ZN(new_n438));
  OAI21_X1  g0238(.A(G68), .B1(new_n438), .B2(new_n423), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n421), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n275), .B1(new_n440), .B2(new_n430), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n441), .A2(KEYINPUT79), .A3(new_n429), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n415), .B1(new_n437), .B2(new_n442), .ZN(new_n443));
  OR2_X1    g0243(.A1(G223), .A2(G1698), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(G226), .B2(new_n255), .ZN(new_n445));
  INV_X1    g0245(.A(G87), .ZN(new_n446));
  OAI22_X1  g0246(.A1(new_n445), .A2(new_n374), .B1(new_n375), .B2(new_n446), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n447), .A2(new_n264), .B1(G232), .B2(new_n342), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n341), .ZN(new_n449));
  NOR3_X1   g0249(.A1(new_n449), .A2(KEYINPUT80), .A3(G179), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT80), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n448), .A2(new_n341), .ZN(new_n452));
  INV_X1    g0252(.A(G179), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n449), .A2(new_n319), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n450), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT18), .B1(new_n443), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n449), .A2(new_n309), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(G190), .B2(new_n449), .ZN(new_n459));
  AND4_X1   g0259(.A1(KEYINPUT79), .A2(new_n429), .A3(new_n294), .A4(new_n434), .ZN(new_n460));
  AOI21_X1  g0260(.A(KEYINPUT79), .B1(new_n441), .B2(new_n429), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n414), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT17), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n414), .B1(new_n460), .B2(new_n461), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT18), .ZN(new_n466));
  INV_X1    g0266(.A(new_n450), .ZN(new_n467));
  INV_X1    g0267(.A(new_n455), .ZN(new_n468));
  OAI21_X1  g0268(.A(KEYINPUT80), .B1(new_n449), .B2(G179), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n465), .A2(new_n466), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n437), .A2(new_n442), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n472), .A2(KEYINPUT17), .A3(new_n414), .A4(new_n459), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n457), .A2(new_n464), .A3(new_n471), .A4(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n352), .A2(new_n409), .A3(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n242), .A2(G45), .ZN(new_n478));
  OR2_X1    g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  NAND2_X1  g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(KEYINPUT81), .A3(new_n250), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT81), .ZN(new_n483));
  INV_X1    g0283(.A(G45), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(G1), .ZN(new_n485));
  INV_X1    g0285(.A(new_n480), .ZN(new_n486));
  NOR2_X1   g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n483), .B1(new_n488), .B2(new_n247), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n481), .A2(new_n264), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n482), .A2(new_n489), .B1(new_n490), .B2(G270), .ZN(new_n491));
  OAI211_X1 g0291(.A(G264), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n492));
  OAI211_X1 g0292(.A(G257), .B(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n493));
  INV_X1    g0293(.A(G303), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n492), .B(new_n493), .C1(new_n494), .C2(new_n335), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n264), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n319), .B1(new_n491), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G283), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n498), .B(new_n285), .C1(G33), .C2(new_n376), .ZN(new_n499));
  INV_X1    g0299(.A(G116), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G20), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n499), .A2(new_n271), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT20), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n499), .A2(KEYINPUT20), .A3(new_n271), .A4(new_n501), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n277), .A2(G20), .A3(new_n500), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n242), .A2(G33), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n275), .A2(new_n278), .A3(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n506), .B(new_n507), .C1(new_n509), .C2(new_n500), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n497), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT21), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n510), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n489), .A2(new_n482), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n490), .A2(G270), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n496), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G200), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n491), .A2(G190), .A3(new_n496), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n514), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AND4_X1   g0320(.A1(G179), .A2(new_n496), .A3(new_n515), .A4(new_n516), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n510), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n510), .A2(KEYINPUT21), .A3(new_n517), .A4(G169), .ZN(new_n523));
  AND4_X1   g0323(.A1(new_n513), .A2(new_n520), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n285), .B(G87), .C1(new_n256), .C2(new_n257), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT22), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT22), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n335), .A2(new_n527), .A3(new_n285), .A4(G87), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT24), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G116), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(G20), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT23), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n285), .B2(G107), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n338), .A2(KEYINPUT23), .A3(G20), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n529), .A2(new_n530), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n530), .B1(new_n529), .B2(new_n536), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n294), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n296), .A2(new_n338), .ZN(new_n540));
  XNOR2_X1  g0340(.A(new_n540), .B(KEYINPUT25), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n509), .A2(new_n338), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n488), .A2(G264), .A3(new_n241), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT82), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n488), .A2(KEYINPUT82), .A3(G264), .A4(new_n241), .ZN(new_n547));
  OAI211_X1 g0347(.A(G257), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n548));
  OAI211_X1 g0348(.A(G250), .B(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n549));
  INV_X1    g0349(.A(G294), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n548), .B(new_n549), .C1(new_n375), .C2(new_n550), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n546), .A2(new_n547), .B1(new_n551), .B2(new_n264), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n552), .A2(G179), .A3(new_n515), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n264), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n554), .A2(new_n515), .A3(new_n544), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G169), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n539), .A2(new_n543), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(G244), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n558));
  OAI211_X1 g0358(.A(G238), .B(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(new_n559), .A3(new_n531), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n264), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n478), .A2(G250), .ZN(new_n562));
  OAI22_X1  g0362(.A1(new_n247), .A2(new_n478), .B1(new_n264), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n561), .A2(new_n564), .A3(G179), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n563), .B1(new_n264), .B2(new_n560), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n565), .B1(new_n319), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n285), .ZN(new_n569));
  NOR2_X1   g0369(.A1(G97), .A2(G107), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n446), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n285), .B(G68), .C1(new_n256), .C2(new_n257), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n326), .A2(new_n376), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n572), .B(new_n573), .C1(KEYINPUT19), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n294), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n296), .A2(new_n325), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n576), .B(new_n577), .C1(new_n509), .C2(new_n325), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n567), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n309), .B1(new_n561), .B2(new_n564), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n275), .A2(G87), .A3(new_n278), .A4(new_n508), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n576), .A2(new_n577), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n566), .A2(G190), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n579), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n557), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n482), .A2(new_n489), .B1(new_n490), .B2(G257), .ZN(new_n588));
  OAI211_X1 g0388(.A(G250), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n589));
  OAI211_X1 g0389(.A(G244), .B(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT4), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n498), .B(new_n589), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n590), .A2(new_n591), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n264), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G200), .ZN(new_n596));
  OAI21_X1  g0396(.A(G107), .B1(new_n438), .B2(new_n423), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n287), .A2(G77), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT6), .ZN(new_n599));
  AND2_X1   g0399(.A1(G97), .A2(G107), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n599), .B1(new_n600), .B2(new_n570), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n338), .A2(KEYINPUT6), .A3(G97), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(G20), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n597), .A2(new_n598), .A3(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n605), .A2(new_n294), .B1(new_n376), .B2(new_n296), .ZN(new_n606));
  INV_X1    g0406(.A(new_n509), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G97), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n588), .A2(new_n594), .A3(G190), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n596), .A2(new_n606), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n604), .A2(new_n598), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n338), .B1(new_n431), .B2(new_n432), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n294), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n296), .A2(new_n376), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n608), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n595), .A2(new_n319), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n588), .A2(new_n594), .A3(new_n453), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n610), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(G200), .B1(new_n552), .B2(new_n515), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n555), .A2(G190), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n539), .B(new_n543), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n524), .A2(new_n587), .A3(new_n619), .A4(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n477), .A2(new_n623), .ZN(G372));
  AND2_X1   g0424(.A1(new_n457), .A2(new_n471), .ZN(new_n625));
  INV_X1    g0425(.A(new_n347), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n408), .A2(new_n366), .B1(new_n401), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n464), .A2(new_n473), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT85), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT85), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n631), .B(new_n625), .C1(new_n627), .C2(new_n628), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n630), .A2(new_n317), .A3(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n633), .A2(new_n322), .ZN(new_n634));
  INV_X1    g0434(.A(new_n578), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n561), .A2(G179), .A3(new_n564), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n319), .B1(new_n561), .B2(new_n564), .ZN(new_n637));
  OAI21_X1  g0437(.A(KEYINPUT83), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT83), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n565), .B(new_n639), .C1(new_n319), .C2(new_n566), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n635), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n585), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n641), .A2(new_n618), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(KEYINPUT84), .B1(new_n643), .B2(KEYINPUT26), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n638), .A2(new_n640), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n578), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(new_n647), .A3(new_n585), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT84), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n580), .B1(G190), .B2(new_n566), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n652), .A2(new_n583), .B1(new_n578), .B2(new_n567), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n647), .A2(new_n653), .A3(KEYINPUT26), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n644), .A2(new_n651), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n522), .A2(new_n523), .ZN(new_n656));
  AOI21_X1  g0456(.A(KEYINPUT21), .B1(new_n497), .B2(new_n510), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n557), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n622), .A2(new_n610), .A3(new_n618), .A4(new_n585), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n646), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n634), .B1(new_n477), .B2(new_n662), .ZN(G369));
  OR2_X1    g0463(.A1(new_n524), .A2(KEYINPUT86), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n524), .A2(KEYINPUT86), .ZN(new_n665));
  INV_X1    g0465(.A(new_n277), .ZN(new_n666));
  OR3_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .A3(G20), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT27), .B1(new_n666), .B2(G20), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n664), .B(new_n665), .C1(new_n514), .C2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n656), .A2(new_n657), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n514), .A2(new_n672), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(G330), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n539), .A2(new_n543), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n671), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n557), .B1(new_n681), .B2(new_n622), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n557), .A2(new_n672), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n674), .A2(new_n671), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n683), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n685), .A2(new_n687), .ZN(G399));
  INV_X1    g0488(.A(new_n208), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(G41), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n571), .A2(G116), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G1), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n213), .B2(new_n691), .ZN(new_n694));
  XOR2_X1   g0494(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n695));
  XNOR2_X1  g0495(.A(new_n694), .B(new_n695), .ZN(new_n696));
  AOI211_X1 g0496(.A(KEYINPUT29), .B(new_n671), .C1(new_n655), .C2(new_n661), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT26), .B1(new_n647), .B2(new_n653), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n698), .B1(KEYINPUT26), .B2(new_n643), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n672), .B1(new_n699), .B2(new_n660), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n700), .A2(KEYINPUT29), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n552), .A2(new_n566), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n588), .A2(new_n594), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n703), .A2(KEYINPUT30), .A3(new_n521), .A4(new_n704), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n588), .A2(new_n594), .B1(new_n566), .B2(KEYINPUT88), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n566), .A2(KEYINPUT88), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n552), .A2(new_n515), .ZN(new_n708));
  AOI21_X1  g0508(.A(G179), .B1(new_n491), .B2(new_n496), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n706), .A2(new_n707), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n705), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT31), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT89), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n703), .A2(new_n521), .A3(new_n704), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT30), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n552), .A2(new_n594), .A3(new_n588), .A4(new_n566), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n491), .A2(G179), .A3(new_n496), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n713), .B(new_n715), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n711), .B(new_n712), .C1(new_n716), .C2(new_n720), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n623), .A2(KEYINPUT31), .B1(new_n721), .B2(new_n671), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n671), .A2(KEYINPUT31), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n714), .A2(new_n715), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n723), .B1(new_n711), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(G330), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n702), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n696), .B1(new_n727), .B2(G1), .ZN(G364));
  AOI21_X1  g0528(.A(G330), .B1(new_n673), .B2(new_n676), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n276), .A2(G20), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n242), .B1(new_n730), .B2(G45), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n690), .A2(new_n732), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n679), .A2(new_n729), .A3(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G13), .A2(G33), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G20), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n677), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n733), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n246), .B1(G20), .B2(new_n319), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n453), .A2(new_n309), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT92), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n285), .A2(G190), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G159), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT32), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n743), .A2(G190), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n376), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n285), .A2(new_n349), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n453), .A2(G200), .ZN(new_n755));
  AND3_X1   g0555(.A1(new_n754), .A2(KEYINPUT91), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(KEYINPUT91), .B1(new_n754), .B2(new_n755), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G58), .ZN(new_n760));
  NAND3_X1  g0560(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G190), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n761), .A2(new_n349), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n763), .A2(new_n203), .B1(new_n765), .B2(new_n201), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n755), .A2(new_n744), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n309), .A2(G179), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n744), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n330), .A2(new_n767), .B1(new_n769), .B2(new_n338), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n754), .A2(new_n768), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n335), .B1(new_n771), .B2(new_n446), .ZN(new_n772));
  NOR3_X1   g0572(.A1(new_n766), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n748), .A2(new_n753), .A3(new_n760), .A4(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n745), .ZN(new_n775));
  AOI22_X1  g0575(.A1(G329), .A2(new_n775), .B1(new_n759), .B2(G322), .ZN(new_n776));
  INV_X1    g0576(.A(G283), .ZN(new_n777));
  INV_X1    g0577(.A(G311), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n777), .A2(new_n769), .B1(new_n767), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n771), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n335), .B(new_n779), .C1(G303), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n750), .A2(G294), .ZN(new_n782));
  XNOR2_X1  g0582(.A(KEYINPUT33), .B(G317), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n762), .A2(new_n783), .B1(new_n764), .B2(G326), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n776), .A2(new_n781), .A3(new_n782), .A4(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n741), .B1(new_n774), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n689), .A2(new_n374), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n787), .A2(G355), .B1(new_n500), .B2(new_n689), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n424), .A2(new_n426), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n689), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(G45), .B2(new_n213), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n238), .A2(new_n484), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n788), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n793), .A2(KEYINPUT90), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n737), .B(new_n740), .C1(new_n793), .C2(KEYINPUT90), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n739), .B(new_n786), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n734), .B1(new_n738), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(G396));
  AOI21_X1  g0598(.A(new_n671), .B1(new_n655), .B2(new_n661), .ZN(new_n799));
  AND3_X1   g0599(.A1(new_n345), .A2(new_n346), .A3(new_n672), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n350), .A2(new_n348), .B1(new_n334), .B2(new_n672), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n800), .B1(new_n801), .B2(new_n347), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n799), .B(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n733), .B1(new_n803), .B2(new_n726), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n726), .B2(new_n803), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n740), .A2(new_n735), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n739), .B1(new_n330), .B2(new_n806), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n763), .A2(new_n777), .B1(new_n765), .B2(new_n494), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n758), .A2(new_n550), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n374), .B1(new_n767), .B2(new_n500), .C1(new_n338), .C2(new_n771), .ZN(new_n810));
  NOR4_X1   g0610(.A1(new_n752), .A2(new_n808), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n745), .A2(new_n778), .B1(new_n446), .B2(new_n769), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT93), .ZN(new_n813));
  INV_X1    g0613(.A(new_n767), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n814), .A2(G159), .B1(G137), .B2(new_n764), .ZN(new_n815));
  INV_X1    g0615(.A(G150), .ZN(new_n816));
  INV_X1    g0616(.A(G143), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n815), .B1(new_n816), .B2(new_n763), .C1(new_n758), .C2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT34), .ZN(new_n819));
  INV_X1    g0619(.A(new_n769), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n780), .A2(G50), .B1(new_n820), .B2(G68), .ZN(new_n821));
  INV_X1    g0621(.A(G132), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n821), .B(new_n789), .C1(new_n822), .C2(new_n745), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(G58), .B2(new_n750), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n811), .A2(new_n813), .B1(new_n819), .B2(new_n824), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n807), .B1(new_n825), .B2(new_n741), .C1(new_n802), .C2(new_n736), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n805), .A2(new_n826), .ZN(G384));
  NAND2_X1  g0627(.A1(new_n408), .A2(new_n366), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n366), .A2(new_n671), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n828), .A2(new_n401), .A3(new_n829), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n366), .B(new_n671), .C1(new_n408), .C2(new_n402), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n801), .A2(new_n347), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n347), .B2(new_n671), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n623), .A2(KEYINPUT31), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n721), .A2(new_n671), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n711), .B1(new_n716), .B2(new_n720), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n838), .A2(KEYINPUT31), .A3(new_n671), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n834), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n421), .B1(new_n428), .B2(new_n203), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n430), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n842), .A2(new_n294), .A3(new_n429), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n669), .B1(new_n843), .B2(new_n414), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n474), .A2(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n456), .A2(new_n669), .B1(new_n414), .B2(new_n843), .ZN(new_n846));
  INV_X1    g0646(.A(new_n462), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT37), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n465), .A2(new_n470), .ZN(new_n849));
  INV_X1    g0649(.A(new_n669), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n465), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT37), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n849), .A2(new_n851), .A3(new_n852), .A4(new_n462), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n848), .A2(new_n853), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n845), .A2(KEYINPUT38), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT38), .B1(new_n845), .B2(new_n854), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n832), .B(new_n840), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT40), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n845), .A2(KEYINPUT38), .A3(new_n854), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n849), .A2(new_n851), .A3(new_n462), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT37), .ZN(new_n862));
  INV_X1    g0662(.A(new_n851), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n862), .A2(new_n853), .B1(new_n474), .B2(new_n863), .ZN(new_n864));
  XNOR2_X1  g0664(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n860), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n867), .A2(KEYINPUT40), .A3(new_n832), .A4(new_n840), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n859), .A2(new_n868), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n869), .B(KEYINPUT96), .Z(new_n870));
  NAND2_X1  g0670(.A1(new_n837), .A2(new_n839), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n476), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n678), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n870), .B2(new_n872), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n476), .B1(new_n697), .B2(new_n701), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n634), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT39), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n867), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n856), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(KEYINPUT39), .A3(new_n860), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n408), .A2(new_n366), .A3(new_n672), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n878), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n671), .B(new_n834), .C1(new_n655), .C2(new_n661), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n800), .B(KEYINPUT94), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  OAI221_X1 g0686(.A(new_n832), .B1(new_n855), .B2(new_n856), .C1(new_n884), .C2(new_n886), .ZN(new_n887));
  OR2_X1    g0687(.A1(new_n625), .A2(new_n850), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n883), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n876), .B(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n874), .A2(new_n890), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n891), .A2(KEYINPUT97), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n891), .A2(KEYINPUT97), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n874), .A2(new_n890), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n730), .A2(new_n242), .ZN(new_n895));
  NOR4_X1   g0695(.A1(new_n892), .A2(new_n893), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n603), .A2(KEYINPUT35), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n603), .A2(KEYINPUT35), .ZN(new_n898));
  NOR4_X1   g0698(.A1(new_n897), .A2(new_n898), .A3(new_n500), .A4(new_n212), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT36), .ZN(new_n900));
  OR3_X1    g0700(.A1(new_n416), .A2(new_n213), .A3(new_n330), .ZN(new_n901));
  AOI211_X1 g0701(.A(new_n242), .B(G13), .C1(new_n901), .C2(new_n234), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n896), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n903), .B(KEYINPUT98), .ZN(G367));
  NAND2_X1  g0704(.A1(new_n615), .A2(new_n671), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n619), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n647), .A2(new_n671), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n685), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n908), .B(KEYINPUT99), .Z(new_n909));
  NAND3_X1  g0709(.A1(new_n619), .A2(new_n557), .A3(new_n905), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n671), .B1(new_n910), .B2(new_n618), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n906), .A2(new_n907), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n912), .A2(new_n684), .A3(new_n686), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n911), .B1(new_n913), .B2(KEYINPUT42), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(KEYINPUT42), .B2(new_n913), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT43), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n672), .A2(new_n583), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n646), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n641), .A2(new_n642), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n918), .B1(new_n919), .B2(new_n917), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n915), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n920), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n921), .B(new_n924), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n909), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n925), .B1(KEYINPUT99), .B2(new_n908), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n687), .A2(new_n912), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT45), .Z(new_n930));
  NOR2_X1   g0730(.A1(new_n687), .A2(new_n912), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT44), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(new_n685), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n684), .B(new_n686), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n679), .B(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n727), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n727), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n690), .B(KEYINPUT41), .Z(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n732), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n928), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n737), .A2(new_n740), .ZN(new_n945));
  INV_X1    g0745(.A(new_n790), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n945), .B1(new_n208), .B2(new_n325), .C1(new_n946), .C2(new_n229), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT100), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n376), .A2(new_n769), .B1(new_n767), .B2(new_n777), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n789), .B(new_n949), .C1(new_n759), .C2(G303), .ZN(new_n950));
  INV_X1    g0750(.A(G317), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n950), .B1(new_n951), .B2(new_n745), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n780), .A2(G116), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT46), .ZN(new_n954));
  AOI22_X1  g0754(.A1(G294), .A2(new_n762), .B1(new_n764), .B2(G311), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n954), .B(new_n955), .C1(new_n751), .C2(new_n338), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n750), .A2(G68), .B1(new_n759), .B2(G150), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT101), .Z(new_n959));
  OAI22_X1  g0759(.A1(new_n763), .A2(new_n746), .B1(new_n765), .B2(new_n817), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n769), .A2(new_n330), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(G50), .B2(new_n814), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n962), .B(new_n335), .C1(new_n202), .C2(new_n771), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n960), .B(new_n963), .C1(G137), .C2(new_n775), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n957), .B1(new_n959), .B2(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT47), .Z(new_n966));
  AOI211_X1 g0766(.A(new_n739), .B(new_n948), .C1(new_n966), .C2(new_n740), .ZN(new_n967));
  INV_X1    g0767(.A(new_n737), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n967), .B1(new_n968), .B2(new_n922), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT102), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n944), .A2(new_n971), .ZN(G387));
  INV_X1    g0772(.A(new_n692), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n973), .A2(new_n787), .B1(new_n338), .B2(new_n689), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n226), .A2(new_n484), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n328), .A2(G50), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT50), .Z(new_n977));
  OAI211_X1 g0777(.A(new_n692), .B(new_n484), .C1(new_n203), .C2(new_n330), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n790), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n974), .B1(new_n975), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n739), .B1(new_n980), .B2(new_n945), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n684), .B2(new_n968), .ZN(new_n982));
  XNOR2_X1  g0782(.A(KEYINPUT103), .B(G150), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n745), .A2(new_n983), .B1(new_n330), .B2(new_n771), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT104), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n410), .A2(new_n763), .B1(new_n765), .B2(new_n746), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n789), .B1(new_n203), .B2(new_n767), .C1(new_n376), .C2(new_n769), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n986), .B(new_n987), .C1(G50), .C2(new_n759), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n751), .A2(new_n325), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n985), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n750), .A2(G283), .B1(G294), .B2(new_n780), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n758), .A2(new_n951), .B1(new_n494), .B2(new_n767), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n992), .A2(KEYINPUT105), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(KEYINPUT105), .ZN(new_n994));
  AOI22_X1  g0794(.A1(G311), .A2(new_n762), .B1(new_n764), .B2(G322), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT48), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n991), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT106), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n996), .A2(new_n997), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n999), .A2(KEYINPUT49), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n789), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n500), .B2(new_n769), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G326), .B2(new_n775), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(KEYINPUT49), .B1(new_n999), .B2(new_n1000), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n990), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n982), .B1(new_n1007), .B2(new_n740), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(new_n936), .B2(new_n732), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n937), .A2(new_n690), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n936), .A2(new_n727), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(G393));
  NAND2_X1  g0812(.A1(new_n939), .A2(new_n690), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n934), .A2(new_n938), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n934), .A2(new_n732), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n912), .A2(new_n968), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT107), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n945), .B1(new_n376), .B2(new_n208), .C1(new_n946), .C2(new_n233), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n771), .A2(new_n777), .B1(new_n767), .B2(new_n550), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n335), .B(new_n1020), .C1(G107), .C2(new_n820), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n775), .A2(G322), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(new_n494), .C2(new_n763), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G116), .B2(new_n750), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n758), .A2(new_n778), .B1(new_n951), .B2(new_n765), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT52), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1002), .B1(G50), .B2(new_n762), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n328), .A2(new_n767), .B1(new_n769), .B2(new_n446), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G68), .B2(new_n780), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1027), .B(new_n1029), .C1(new_n817), .C2(new_n745), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G77), .B2(new_n750), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n758), .A2(new_n746), .B1(new_n816), .B2(new_n765), .ZN(new_n1032));
  XOR2_X1   g0832(.A(KEYINPUT108), .B(KEYINPUT51), .Z(new_n1033));
  XNOR2_X1  g0833(.A(new_n1032), .B(new_n1033), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n1024), .A2(new_n1026), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n733), .B(new_n1019), .C1(new_n1035), .C2(new_n741), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1016), .B1(new_n1018), .B2(new_n1036), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1015), .A2(new_n1037), .ZN(G390));
  NAND3_X1  g0838(.A1(new_n476), .A2(G330), .A3(new_n871), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n633), .A2(new_n322), .A3(new_n875), .A4(new_n1039), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n884), .A2(new_n886), .ZN(new_n1041));
  OAI211_X1 g0841(.A(G330), .B(new_n802), .C1(new_n722), .C2(new_n725), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1042), .A2(KEYINPUT110), .A3(new_n830), .A4(new_n831), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n832), .A2(new_n840), .A3(G330), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n830), .A2(new_n831), .ZN(new_n1046));
  AOI21_X1  g0846(.A(KEYINPUT110), .B1(new_n1046), .B2(new_n1042), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1041), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1046), .A2(new_n1042), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n672), .B(new_n802), .C1(new_n699), .C2(new_n660), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n885), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(KEYINPUT109), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT109), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1050), .A2(new_n1053), .A3(new_n885), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n840), .A2(G330), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n1046), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1049), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1040), .B1(new_n1048), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1044), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n832), .B1(new_n884), .B2(new_n886), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n878), .A2(new_n880), .B1(new_n1061), .B2(new_n881), .ZN(new_n1062));
  AND3_X1   g0862(.A1(new_n1052), .A2(new_n832), .A3(new_n1054), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n867), .A2(new_n881), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1060), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n878), .A2(new_n880), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1061), .A2(new_n881), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n881), .B(new_n867), .C1(new_n1055), .C2(new_n1046), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1069), .A2(new_n1070), .A3(new_n1049), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1059), .A2(new_n1066), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1066), .A2(new_n1071), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1059), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT111), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(KEYINPUT111), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n690), .B(new_n1072), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1067), .A2(new_n735), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n739), .B1(new_n410), .B2(new_n806), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n765), .A2(new_n777), .B1(new_n767), .B2(new_n376), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(G107), .B2(new_n762), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT113), .Z(new_n1084));
  OAI221_X1 g0884(.A(new_n374), .B1(new_n769), .B2(new_n203), .C1(new_n446), .C2(new_n771), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n758), .A2(new_n500), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(G294), .C2(new_n775), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1084), .B(new_n1087), .C1(new_n330), .C2(new_n751), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1088), .A2(KEYINPUT114), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1088), .A2(KEYINPUT114), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n771), .A2(new_n983), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT53), .Z(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G125), .B2(new_n775), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n374), .B1(new_n820), .B2(G50), .ZN(new_n1094));
  INV_X1    g0894(.A(G128), .ZN(new_n1095));
  INV_X1    g0895(.A(G137), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1094), .B1(new_n765), .B2(new_n1095), .C1(new_n1096), .C2(new_n763), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G159), .B2(new_n750), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(KEYINPUT54), .B(G143), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT112), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n759), .A2(G132), .B1(new_n814), .B2(new_n1100), .ZN(new_n1101));
  AND3_X1   g0901(.A1(new_n1093), .A2(new_n1098), .A3(new_n1101), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n1089), .A2(new_n1090), .A3(new_n1102), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1080), .B(new_n1081), .C1(new_n741), .C2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n1073), .B2(new_n731), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n1105), .A2(KEYINPUT115), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(KEYINPUT115), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1079), .A2(new_n1106), .A3(new_n1107), .ZN(G378));
  NAND2_X1  g0908(.A1(new_n321), .A2(new_n850), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT55), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT117), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n317), .A2(new_n1112), .A3(new_n322), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1112), .B1(new_n317), .B2(new_n322), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1111), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n323), .A2(KEYINPUT117), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n317), .A2(new_n1112), .A3(new_n322), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n1110), .A3(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1119));
  AND3_X1   g0919(.A1(new_n1115), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1119), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n735), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1002), .B1(new_n765), .B2(new_n500), .C1(new_n376), .C2(new_n763), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(G68), .B2(new_n750), .ZN(new_n1125));
  INV_X1    g0925(.A(G41), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n771), .B2(new_n330), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n325), .A2(new_n767), .B1(new_n769), .B2(new_n202), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1127), .B(new_n1128), .C1(new_n775), .C2(G283), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1125), .B(new_n1129), .C1(new_n338), .C2(new_n758), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT58), .ZN(new_n1131));
  AOI21_X1  g0931(.A(G41), .B1(new_n789), .B2(G33), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n759), .A2(G128), .B1(new_n780), .B2(new_n1100), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n764), .A2(G125), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n1096), .B2(new_n767), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G132), .B2(new_n762), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1133), .B(new_n1136), .C1(new_n816), .C2(new_n751), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1137), .A2(KEYINPUT59), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(KEYINPUT59), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n375), .B(new_n1126), .C1(new_n769), .C2(new_n746), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n775), .B2(G124), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1131), .B1(G50), .B2(new_n1132), .C1(new_n1138), .C2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n741), .B1(new_n1143), .B2(KEYINPUT116), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(KEYINPUT116), .B2(new_n1143), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n739), .B1(new_n201), .B2(new_n806), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1123), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT119), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n859), .A2(G330), .A3(new_n868), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1122), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n678), .B1(new_n857), .B2(new_n858), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1153), .A2(new_n868), .A3(new_n1122), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1152), .A2(new_n889), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n889), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1149), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n889), .ZN(new_n1158));
  AND4_X1   g0958(.A1(G330), .A2(new_n859), .A3(new_n1122), .A4(new_n868), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1122), .B1(new_n1153), .B2(new_n868), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1152), .A2(new_n889), .A3(new_n1154), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1161), .A2(KEYINPUT119), .A3(new_n1162), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n1157), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1148), .B1(new_n1164), .B2(new_n732), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT57), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1040), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1166), .B1(new_n1072), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT120), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1156), .A2(KEYINPUT120), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1168), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1172), .A2(KEYINPUT121), .A3(new_n690), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1072), .A2(new_n1167), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1157), .A2(new_n1174), .A3(new_n1163), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n1166), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(KEYINPUT121), .B1(new_n1172), .B2(new_n690), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1165), .B1(new_n1177), .B2(new_n1178), .ZN(G375));
  NAND2_X1  g0979(.A1(new_n1048), .A2(new_n1058), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(KEYINPUT122), .B1(new_n1181), .B2(new_n731), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT122), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1180), .A2(new_n1183), .A3(new_n732), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n759), .A2(G283), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n775), .A2(G303), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n335), .B(new_n961), .C1(G97), .C2(new_n780), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n989), .A2(new_n1185), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n765), .A2(new_n550), .B1(new_n767), .B2(new_n338), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G116), .B2(new_n762), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT123), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1100), .A2(new_n762), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1192), .B1(new_n1095), .B2(new_n745), .C1(new_n1096), .C2(new_n758), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n202), .A2(new_n769), .B1(new_n767), .B2(new_n816), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G159), .B2(new_n780), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1002), .B1(G132), .B2(new_n764), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1195), .B(new_n1196), .C1(new_n751), .C2(new_n201), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n1188), .A2(new_n1191), .B1(new_n1193), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n740), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n739), .B1(new_n203), .B2(new_n806), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(new_n832), .C2(new_n736), .ZN(new_n1201));
  AND3_X1   g1001(.A1(new_n1182), .A2(new_n1184), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1181), .A2(new_n1040), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1203), .A2(new_n1074), .A3(new_n942), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1202), .A2(new_n1204), .ZN(G381));
  OR2_X1    g1005(.A1(G393), .A2(G396), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(G390), .A2(G384), .A3(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1207), .A2(new_n971), .A3(new_n944), .ZN(new_n1208));
  OR4_X1    g1008(.A1(G378), .A2(new_n1208), .A3(G375), .A4(G381), .ZN(G407));
  OR2_X1    g1009(.A1(G375), .A2(G378), .ZN(new_n1210));
  OAI211_X1 g1010(.A(G407), .B(G213), .C1(G343), .C2(new_n1210), .ZN(G409));
  OAI211_X1 g1011(.A(G378), .B(new_n1165), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n732), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1147), .B(new_n1213), .C1(new_n1175), .C2(new_n941), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1214), .A2(new_n1079), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1212), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n670), .A2(G213), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1074), .A2(KEYINPUT60), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n1203), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1048), .A2(new_n1040), .A3(new_n1058), .A4(KEYINPUT60), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n690), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1220), .A2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1224), .A2(new_n1202), .A3(G384), .ZN(new_n1225));
  INV_X1    g1025(.A(G384), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1222), .B1(new_n1219), .B2(new_n1203), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1182), .A2(new_n1184), .A3(new_n1201), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1226), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1225), .A2(new_n1229), .A3(KEYINPUT124), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1217), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n1231), .A2(G2897), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1225), .A2(new_n1229), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT124), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1233), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1234), .A2(new_n1235), .A3(new_n1232), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT61), .B1(new_n1218), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1234), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1216), .A2(new_n1217), .A3(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT63), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1206), .ZN(new_n1245));
  AND2_X1   g1045(.A1(G393), .A2(G396), .ZN(new_n1246));
  OAI21_X1  g1046(.A(KEYINPUT125), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G390), .B(new_n971), .C1(new_n943), .C2(new_n928), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(G390), .B1(new_n944), .B2(new_n971), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1247), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(G390), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G387), .A2(new_n1252), .ZN(new_n1253));
  OR3_X1    g1053(.A1(new_n1245), .A2(KEYINPUT125), .A3(new_n1246), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1247), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1253), .A2(new_n1255), .A3(new_n1248), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1251), .A2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1231), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(KEYINPUT63), .A3(new_n1241), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1240), .A2(new_n1244), .A3(new_n1257), .A4(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT61), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1261), .B1(new_n1258), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT62), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1242), .A2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1258), .A2(KEYINPUT62), .A3(new_n1241), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1263), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1257), .B(KEYINPUT126), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1260), .B1(new_n1267), .B2(new_n1268), .ZN(G405));
  INV_X1    g1069(.A(KEYINPUT127), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1251), .A2(new_n1256), .A3(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1270), .B1(new_n1251), .B2(new_n1256), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G375), .A2(G378), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1210), .A2(new_n1234), .A3(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1234), .B1(new_n1210), .B2(new_n1274), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1273), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1277), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1279), .A2(new_n1271), .A3(new_n1275), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1278), .A2(new_n1280), .ZN(G402));
endmodule


