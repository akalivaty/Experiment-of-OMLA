//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 0 0 1 1 0 1 0 0 1 1 0 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1205, new_n1206, new_n1207;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT67), .B(G57), .Z(G237));
  XOR2_X1   g015(.A(KEYINPUT68), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT69), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g025(.A1(G221), .A2(G218), .A3(G219), .A4(G220), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n452), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OR2_X1    g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n471), .A2(G137), .B1(G101), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  NOR2_X1   g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT70), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n472), .B1(new_n469), .B2(new_n470), .ZN(new_n480));
  AOI22_X1  g055(.A1(G124), .A2(new_n480), .B1(new_n471), .B2(G136), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n479), .A2(new_n481), .ZN(G162));
  OAI211_X1 g057(.A(G138), .B(new_n472), .C1(new_n462), .C2(new_n463), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT4), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n469), .A2(new_n470), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n485), .A2(new_n486), .A3(G138), .A4(new_n472), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  OR2_X1    g063(.A1(new_n472), .A2(G114), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  AOI22_X1  g066(.A1(new_n480), .A2(G126), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AND3_X1   g067(.A1(new_n488), .A2(KEYINPUT71), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(KEYINPUT71), .B1(new_n488), .B2(new_n492), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  NAND2_X1  g071(.A1(G75), .A2(G543), .ZN(new_n497));
  INV_X1    g072(.A(G62), .ZN(new_n498));
  OR2_X1    g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT73), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n497), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT5), .B(G543), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(new_n502), .A3(G62), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  OAI21_X1  g081(.A(G651), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT74), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  OAI21_X1  g086(.A(G62), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(KEYINPUT73), .B1(G75), .B2(G543), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n509), .B1(new_n513), .B2(new_n505), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT74), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n517), .B1(new_n509), .B2(KEYINPUT6), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n519), .A2(KEYINPUT72), .A3(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n509), .A2(KEYINPUT6), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n521), .A2(G88), .A3(new_n504), .A4(new_n522), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n521), .A2(G50), .A3(G543), .A4(new_n522), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n508), .A2(new_n516), .A3(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(G166));
  AOI22_X1  g102(.A1(new_n518), .A2(new_n520), .B1(KEYINPUT6), .B2(new_n509), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n528), .A2(G51), .A3(G543), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n528), .A2(G89), .A3(new_n504), .ZN(new_n530));
  AND2_X1   g105(.A1(G63), .A2(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT7), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n534), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n504), .A2(new_n531), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  AND3_X1   g111(.A1(new_n529), .A2(new_n530), .A3(new_n536), .ZN(G168));
  AOI22_X1  g112(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(new_n509), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n521), .A2(G52), .A3(G543), .A4(new_n522), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n521), .A2(G90), .A3(new_n504), .A4(new_n522), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT75), .ZN(new_n542));
  AND3_X1   g117(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n542), .B1(new_n540), .B2(new_n541), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n539), .B1(new_n543), .B2(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  INV_X1    g121(.A(G56), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n547), .B1(new_n499), .B2(new_n500), .ZN(new_n548));
  AND2_X1   g123(.A1(G68), .A2(G543), .ZN(new_n549));
  OAI21_X1  g124(.A(G651), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND4_X1  g125(.A1(new_n521), .A2(G81), .A3(new_n504), .A4(new_n522), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n521), .A2(G43), .A3(G543), .A4(new_n522), .ZN(new_n552));
  AND3_X1   g127(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  NAND4_X1  g133(.A1(new_n521), .A2(G53), .A3(G543), .A4(new_n522), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT9), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n504), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n561), .A2(new_n509), .ZN(new_n562));
  AND3_X1   g137(.A1(new_n519), .A2(KEYINPUT72), .A3(G651), .ZN(new_n563));
  AOI21_X1  g138(.A(KEYINPUT72), .B1(new_n519), .B2(G651), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n504), .B(new_n522), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(KEYINPUT76), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n528), .A2(new_n567), .A3(new_n504), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(G91), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n560), .A2(new_n562), .A3(new_n569), .ZN(G299));
  NAND3_X1  g145(.A1(new_n529), .A2(new_n530), .A3(new_n536), .ZN(G286));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n525), .B1(new_n514), .B2(new_n515), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n507), .A2(KEYINPUT74), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n508), .A2(new_n516), .A3(KEYINPUT77), .A4(new_n525), .ZN(new_n576));
  AND2_X1   g151(.A1(new_n575), .A2(new_n576), .ZN(G303));
  NAND3_X1  g152(.A1(new_n521), .A2(G543), .A3(new_n522), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n504), .A2(G74), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n579), .A2(G49), .B1(G651), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n566), .A2(G87), .A3(new_n568), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G288));
  OAI21_X1  g158(.A(G61), .B1(new_n510), .B2(new_n511), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n509), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n586), .A2(KEYINPUT78), .ZN(new_n587));
  AND2_X1   g162(.A1(G48), .A2(G543), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n586), .A2(KEYINPUT78), .B1(new_n528), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n566), .A2(G86), .A3(new_n568), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G305));
  INV_X1    g167(.A(G47), .ZN(new_n593));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n593), .A2(new_n578), .B1(new_n565), .B2(new_n594), .ZN(new_n595));
  AND2_X1   g170(.A1(new_n595), .A2(KEYINPUT79), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n595), .A2(KEYINPUT79), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  OAI22_X1  g173(.A1(new_n596), .A2(new_n597), .B1(new_n509), .B2(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n504), .A2(G66), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G651), .ZN(new_n604));
  INV_X1    g179(.A(G54), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n578), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n566), .A2(G92), .A3(new_n568), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n566), .A2(KEYINPUT10), .A3(new_n568), .A4(G92), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n600), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n600), .B1(new_n611), .B2(G868), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT80), .Z(new_n615));
  INV_X1    g190(.A(G299), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(G868), .B2(new_n616), .ZN(G297));
  OAI21_X1  g192(.A(new_n615), .B1(G868), .B2(new_n616), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n611), .B1(new_n619), .B2(G860), .ZN(G148));
  INV_X1    g195(.A(new_n553), .ZN(new_n621));
  INV_X1    g196(.A(G868), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n609), .A2(new_n610), .ZN(new_n624));
  INV_X1    g199(.A(new_n606), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n626), .A2(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n623), .B1(new_n627), .B2(new_n622), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g204(.A1(new_n485), .A2(new_n473), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  INV_X1    g207(.A(G2100), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n471), .A2(G135), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n480), .A2(G123), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n472), .A2(G111), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n636), .B(new_n637), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(G2096), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n634), .A2(new_n635), .A3(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2427), .B(G2430), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(KEYINPUT14), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT81), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n649), .B1(new_n645), .B2(new_n646), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n654), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(new_n658), .A3(G14), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(G401));
  INV_X1    g235(.A(KEYINPUT18), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n661), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT82), .B(G2100), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2072), .B(G2078), .Z(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n664), .B2(KEYINPUT18), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(new_n641), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n669), .B(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1956), .B(G2474), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT83), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1961), .B(G1966), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT20), .Z(new_n682));
  NOR2_X1   g257(.A1(new_n675), .A2(new_n677), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n684), .A2(new_n680), .A3(new_n678), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n682), .B(new_n685), .C1(new_n680), .C2(new_n684), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n690), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(G229));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G32), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n480), .A2(G129), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT91), .Z(new_n698));
  AND2_X1   g273(.A1(new_n473), .A2(G105), .ZN(new_n699));
  NAND3_X1  g274(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT26), .ZN(new_n701));
  AOI211_X1 g276(.A(new_n699), .B(new_n701), .C1(G141), .C2(new_n471), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n696), .B1(new_n704), .B2(new_n695), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT92), .Z(new_n706));
  XOR2_X1   g281(.A(KEYINPUT27), .B(G1996), .Z(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NOR2_X1   g284(.A1(G171), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G5), .B2(new_n709), .ZN(new_n711));
  INV_X1    g286(.A(G1961), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT24), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n714), .A2(G34), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n695), .B1(new_n714), .B2(G34), .ZN(new_n716));
  OAI22_X1  g291(.A1(new_n475), .A2(new_n695), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G2084), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n708), .A2(new_n713), .A3(new_n719), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT95), .Z(new_n721));
  NOR2_X1   g296(.A1(G4), .A2(G16), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n611), .B2(G16), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT86), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT87), .B(G1348), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n695), .A2(G35), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G162), .B2(new_n695), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT29), .Z(new_n729));
  INV_X1    g304(.A(G2090), .ZN(new_n730));
  NOR2_X1   g305(.A1(G16), .A2(G19), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n553), .B2(G16), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n729), .A2(new_n730), .B1(G1341), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n709), .A2(G21), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G168), .B2(new_n709), .ZN(new_n735));
  INV_X1    g310(.A(G1966), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n733), .B(new_n737), .C1(new_n712), .C2(new_n711), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT30), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT94), .ZN(new_n740));
  AND3_X1   g315(.A1(new_n740), .A2(new_n739), .A3(G28), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n740), .B1(new_n739), .B2(G28), .ZN(new_n742));
  OAI221_X1 g317(.A(new_n695), .B1(new_n739), .B2(G28), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT31), .B(G11), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n640), .A2(new_n695), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(KEYINPUT93), .ZN(new_n747));
  OAI221_X1 g322(.A(new_n747), .B1(KEYINPUT93), .B2(new_n746), .C1(new_n718), .C2(new_n717), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n695), .A2(G26), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n471), .A2(G140), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n480), .A2(G128), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n472), .A2(G116), .ZN(new_n754));
  OAI21_X1  g329(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n752), .B(new_n753), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n751), .B1(new_n756), .B2(G29), .ZN(new_n757));
  INV_X1    g332(.A(G2067), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n748), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n695), .A2(G27), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G164), .B2(new_n695), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G2078), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n695), .A2(G33), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT89), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT25), .ZN(new_n767));
  NAND2_X1  g342(.A1(G115), .A2(G2104), .ZN(new_n768));
  INV_X1    g343(.A(G127), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n464), .B2(new_n769), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n770), .A2(G2105), .B1(G139), .B2(new_n471), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT90), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n764), .B1(new_n774), .B2(new_n695), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n763), .B1(new_n775), .B2(G2072), .ZN(new_n776));
  OAI22_X1  g351(.A1(new_n729), .A2(new_n730), .B1(G1341), .B2(new_n732), .ZN(new_n777));
  NOR4_X1   g352(.A1(new_n738), .A2(new_n760), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n709), .A2(G20), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT23), .Z(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G299), .B2(G16), .ZN(new_n781));
  INV_X1    g356(.A(G1956), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  OAI22_X1  g358(.A1(new_n706), .A2(new_n707), .B1(G2078), .B2(new_n762), .ZN(new_n784));
  AOI211_X1 g359(.A(new_n783), .B(new_n784), .C1(G2072), .C2(new_n775), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n721), .A2(new_n726), .A3(new_n778), .A4(new_n785), .ZN(new_n786));
  MUX2_X1   g361(.A(G6), .B(G305), .S(G16), .Z(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT32), .B(G1981), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n709), .A2(G22), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G166), .B2(new_n709), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n789), .B1(G1971), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n709), .A2(G23), .ZN(new_n793));
  INV_X1    g368(.A(G288), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(new_n709), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT33), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G1976), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n792), .B(new_n797), .C1(G1971), .C2(new_n791), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n798), .A2(KEYINPUT34), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(KEYINPUT34), .ZN(new_n800));
  INV_X1    g375(.A(G290), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT84), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n801), .A2(new_n802), .ZN(new_n805));
  OAI21_X1  g380(.A(G16), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G16), .B2(G24), .ZN(new_n807));
  INV_X1    g382(.A(G1986), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n471), .A2(G131), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n480), .A2(G119), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n472), .A2(G107), .ZN(new_n812));
  OAI21_X1  g387(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n810), .B(new_n811), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  MUX2_X1   g389(.A(G25), .B(new_n814), .S(G29), .Z(new_n815));
  XOR2_X1   g390(.A(KEYINPUT35), .B(G1991), .Z(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n815), .B(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n809), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n799), .A2(new_n800), .A3(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT85), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n820), .A2(new_n821), .A3(KEYINPUT36), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(KEYINPUT36), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n799), .A2(new_n823), .A3(new_n800), .A4(new_n819), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n786), .B1(new_n822), .B2(new_n824), .ZN(G311));
  INV_X1    g400(.A(G311), .ZN(G150));
  NAND2_X1  g401(.A1(new_n611), .A2(G559), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT96), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT38), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n521), .A2(G93), .A3(new_n504), .A4(new_n522), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n521), .A2(G55), .A3(G543), .A4(new_n522), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n830), .B(new_n831), .C1(new_n509), .C2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n553), .B(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n829), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(KEYINPUT39), .ZN(new_n836));
  INV_X1    g411(.A(new_n834), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n829), .B(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT39), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(G860), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n836), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n833), .A2(G860), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT37), .Z(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT97), .ZN(G145));
  XNOR2_X1  g421(.A(new_n774), .B(new_n703), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n480), .A2(G130), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n472), .A2(G118), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(G142), .B2(new_n471), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(new_n631), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n847), .B(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT98), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n484), .A2(new_n487), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n855), .B1(new_n484), .B2(new_n487), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n492), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n756), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n814), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n475), .B(new_n640), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(G162), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n854), .A2(new_n860), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n861), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(G37), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n863), .B1(new_n861), .B2(new_n864), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT40), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(G395));
  NAND2_X1  g446(.A1(new_n833), .A2(new_n622), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT100), .ZN(new_n873));
  AND2_X1   g448(.A1(G290), .A2(G288), .ZN(new_n874));
  NOR2_X1   g449(.A1(G290), .A2(G288), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n801), .A2(new_n794), .ZN(new_n877));
  NAND2_X1  g452(.A1(G290), .A2(G288), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n877), .A2(KEYINPUT100), .A3(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(G305), .B(new_n526), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n876), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n880), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n877), .A2(new_n878), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n883), .A3(new_n873), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT42), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n624), .A2(G299), .A3(new_n625), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n611), .A2(G299), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT41), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n890), .B1(new_n887), .B2(new_n888), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n626), .A2(new_n616), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n611), .A2(G299), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(KEYINPUT41), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(new_n894), .A3(KEYINPUT99), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT99), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n889), .A2(new_n896), .A3(KEYINPUT41), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n627), .B(new_n837), .ZN(new_n899));
  MUX2_X1   g474(.A(new_n889), .B(new_n898), .S(new_n899), .Z(new_n900));
  XNOR2_X1  g475(.A(new_n886), .B(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n872), .B1(new_n901), .B2(new_n622), .ZN(G295));
  OAI21_X1  g477(.A(new_n872), .B1(new_n901), .B2(new_n622), .ZN(G331));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n904));
  NAND2_X1  g479(.A1(G168), .A2(KEYINPUT101), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT101), .ZN(new_n906));
  NAND2_X1  g481(.A1(G286), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(G301), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n540), .A2(new_n541), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT75), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n912), .A2(KEYINPUT101), .A3(G168), .A4(new_n539), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n834), .B1(new_n908), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n908), .A2(new_n913), .A3(new_n834), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(KEYINPUT102), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT102), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n908), .A2(new_n913), .A3(new_n834), .A4(new_n918), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n895), .A2(new_n897), .A3(new_n917), .A4(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT104), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n892), .A2(new_n893), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n916), .A2(KEYINPUT103), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n923), .A2(new_n914), .ZN(new_n924));
  AOI211_X1 g499(.A(KEYINPUT103), .B(new_n834), .C1(new_n913), .C2(new_n908), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n921), .B(new_n922), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n920), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n915), .A2(KEYINPUT103), .A3(new_n916), .ZN(new_n928));
  INV_X1    g503(.A(new_n925), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n921), .B1(new_n930), .B2(new_n922), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n885), .B1(new_n927), .B2(new_n931), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n881), .A2(new_n884), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT104), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n933), .A2(new_n935), .A3(new_n920), .A4(new_n926), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n932), .A2(new_n866), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n891), .A2(KEYINPUT105), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n922), .A2(new_n941), .A3(new_n890), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n930), .B1(new_n943), .B2(new_n894), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n889), .B1(new_n917), .B2(new_n919), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n885), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n946), .A2(new_n936), .A3(KEYINPUT43), .A4(new_n866), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n904), .B1(new_n939), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n946), .A2(new_n936), .A3(new_n938), .A4(new_n866), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT44), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT106), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n935), .A2(new_n920), .A3(new_n926), .ZN(new_n953));
  AOI21_X1  g528(.A(G37), .B1(new_n953), .B2(new_n885), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT43), .B1(new_n954), .B2(new_n936), .ZN(new_n955));
  INV_X1    g530(.A(new_n947), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT44), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n938), .B1(new_n954), .B2(new_n936), .ZN(new_n958));
  INV_X1    g533(.A(new_n950), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n904), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n957), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n952), .A2(new_n962), .ZN(G397));
  NAND2_X1  g538(.A1(new_n616), .A2(KEYINPUT57), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT117), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n569), .A2(new_n965), .A3(new_n562), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n965), .B1(new_n569), .B2(new_n562), .ZN(new_n967));
  XOR2_X1   g542(.A(new_n559), .B(KEYINPUT9), .Z(new_n968));
  NOR3_X1   g543(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n964), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n486), .B1(new_n471), .B2(G138), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n483), .A2(KEYINPUT4), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n492), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT71), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT50), .ZN(new_n978));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n488), .A2(KEYINPUT71), .A3(new_n492), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n977), .A2(new_n978), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n468), .A2(G40), .A3(new_n474), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n978), .B1(new_n858), .B2(new_n979), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n782), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n977), .A2(new_n979), .A3(new_n980), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n988), .A2(G1384), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n982), .B1(new_n858), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(KEYINPUT56), .B(G2072), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n989), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n972), .B1(new_n986), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n858), .A2(new_n979), .A3(new_n983), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n995), .A2(G2067), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n858), .A2(new_n978), .A3(new_n979), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n493), .A2(new_n494), .A3(G1384), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n997), .B(new_n983), .C1(new_n998), .C2(new_n978), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n996), .B1(new_n999), .B2(new_n725), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(new_n626), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n972), .A2(new_n986), .A3(new_n993), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n994), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT61), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n986), .A2(new_n993), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n967), .A2(new_n968), .ZN(new_n1006));
  INV_X1    g581(.A(new_n966), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n1008), .A2(new_n970), .B1(KEYINPUT57), .B2(new_n616), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1004), .B1(new_n1010), .B2(new_n994), .ZN(new_n1011));
  AOI211_X1 g586(.A(new_n611), .B(new_n996), .C1(new_n999), .C2(new_n725), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT60), .B1(new_n1001), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT60), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1000), .A2(new_n1014), .A3(new_n611), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1016), .A2(KEYINPUT61), .A3(new_n1002), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1011), .A2(new_n1013), .A3(new_n1015), .A4(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT59), .ZN(new_n1019));
  INV_X1    g594(.A(G1996), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n989), .A2(new_n1020), .A3(new_n991), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT118), .ZN(new_n1022));
  XOR2_X1   g597(.A(KEYINPUT58), .B(G1341), .Z(new_n1023));
  AOI22_X1  g598(.A1(new_n1021), .A2(new_n1022), .B1(new_n995), .B2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n989), .A2(KEYINPUT118), .A3(new_n991), .A4(new_n1020), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1019), .B1(new_n1026), .B2(new_n553), .ZN(new_n1027));
  AOI211_X1 g602(.A(KEYINPUT59), .B(new_n621), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1003), .B1(new_n1018), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT119), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT119), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1032), .B(new_n1003), .C1(new_n1018), .C2(new_n1029), .ZN(new_n1033));
  XOR2_X1   g608(.A(KEYINPUT123), .B(KEYINPUT54), .Z(new_n1034));
  XNOR2_X1  g609(.A(KEYINPUT125), .B(KEYINPUT53), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n989), .A2(new_n991), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1035), .B1(new_n1036), .B2(G2078), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT98), .B1(new_n973), .B2(new_n974), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n484), .A2(new_n487), .A3(new_n855), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1384), .B1(new_n1040), .B2(new_n492), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n982), .B1(new_n1041), .B2(new_n978), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n987), .A2(KEYINPUT50), .ZN(new_n1043));
  AOI21_X1  g618(.A(G1961), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT124), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n977), .A2(new_n980), .A3(new_n990), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n983), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT45), .B1(new_n858), .B2(new_n979), .ZN(new_n1048));
  INV_X1    g623(.A(G2078), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT53), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1047), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n1044), .A2(new_n1045), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n999), .A2(new_n712), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1048), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1050), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1054), .A2(new_n983), .A3(new_n1046), .A4(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT124), .B1(new_n1053), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1037), .B1(new_n1052), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(G171), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1054), .A2(new_n991), .A3(new_n1055), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1037), .A2(new_n1053), .A3(new_n1060), .ZN(new_n1061));
  OR2_X1    g636(.A1(new_n1061), .A2(G171), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1034), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n575), .A2(G8), .A3(new_n576), .ZN(new_n1064));
  NAND2_X1  g639(.A1(KEYINPUT111), .A2(KEYINPUT55), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  XOR2_X1   g641(.A(KEYINPUT111), .B(KEYINPUT55), .Z(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n575), .A2(G8), .A3(new_n576), .A4(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  XOR2_X1   g645(.A(KEYINPUT109), .B(G1971), .Z(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT45), .B1(new_n495), .B2(new_n979), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n858), .A2(new_n990), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n983), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1072), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT110), .B(G2090), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1043), .A2(new_n1077), .A3(new_n983), .A4(new_n997), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1070), .A2(G8), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1976), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n995), .B(G8), .C1(new_n1081), .C2(G288), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT52), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT52), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n794), .B2(G1976), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n995), .A2(G8), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n586), .B1(new_n528), .B2(new_n588), .ZN(new_n1089));
  INV_X1    g664(.A(G86), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1089), .B1(new_n1090), .B2(new_n565), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1091), .A2(G1981), .ZN(new_n1092));
  XOR2_X1   g667(.A(KEYINPUT112), .B(G1981), .Z(new_n1093));
  NAND4_X1  g668(.A1(new_n590), .A2(KEYINPUT113), .A3(new_n591), .A4(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n591), .A2(new_n587), .A3(new_n589), .A4(new_n1093), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT113), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1092), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1088), .B1(new_n1098), .B2(KEYINPUT49), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT49), .ZN(new_n1100));
  AOI211_X1 g675(.A(new_n1100), .B(new_n1092), .C1(new_n1097), .C2(new_n1094), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1083), .B(new_n1086), .C1(new_n1099), .C2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1080), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT114), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1077), .ZN(new_n1105));
  NOR3_X1   g680(.A1(new_n984), .A2(new_n1105), .A3(new_n985), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1071), .B1(new_n989), .B2(new_n991), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1104), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n858), .A2(new_n979), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(KEYINPUT50), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1110), .A2(new_n1077), .A3(new_n983), .A4(new_n981), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1076), .A2(KEYINPUT114), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1108), .A2(G8), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1070), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1035), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1116), .B1(new_n1117), .B2(new_n1049), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1045), .B1(new_n1044), .B2(new_n1051), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1053), .A2(KEYINPUT124), .A3(new_n1056), .ZN(new_n1120));
  AOI211_X1 g695(.A(G171), .B(new_n1118), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1061), .A2(G171), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT54), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1103), .B(new_n1115), .C1(new_n1121), .C2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1063), .A2(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT120), .B(KEYINPUT51), .ZN(new_n1126));
  INV_X1    g701(.A(G8), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n736), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1043), .A2(new_n718), .A3(new_n983), .A4(new_n997), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1127), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(G168), .A2(new_n1127), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1126), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g709(.A(KEYINPUT121), .B(new_n1126), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1130), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1136), .A2(KEYINPUT122), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1131), .A2(KEYINPUT51), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1138), .B1(new_n1130), .B2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1134), .B(new_n1135), .C1(new_n1137), .C2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n1131), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1031), .A2(new_n1033), .A3(new_n1125), .A4(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1099), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1101), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(G288), .A2(G1976), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1148), .A2(new_n1149), .B1(new_n1097), .B2(new_n1094), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1070), .A2(new_n1079), .A3(G8), .ZN(new_n1151));
  OAI22_X1  g726(.A1(new_n1150), .A2(new_n1087), .B1(new_n1151), .B2(new_n1102), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1083), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1153), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1136), .A2(G286), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1115), .A2(new_n1151), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(KEYINPUT115), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT63), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT115), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1103), .A2(new_n1159), .A3(new_n1115), .A4(new_n1155), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1157), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1079), .A2(G8), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(new_n1114), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1103), .A2(KEYINPUT63), .A3(new_n1155), .A4(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1152), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1144), .A2(KEYINPUT62), .ZN(new_n1166));
  AND4_X1   g741(.A1(G171), .A2(new_n1103), .A3(new_n1115), .A4(new_n1058), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT62), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1141), .A2(new_n1168), .A3(new_n1143), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1166), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1145), .A2(new_n1165), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1048), .A2(new_n983), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1172), .A2(new_n1020), .A3(new_n704), .ZN(new_n1173));
  OR2_X1    g748(.A1(new_n1173), .A2(KEYINPUT108), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(KEYINPUT108), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1172), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n756), .B(new_n758), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1177), .B1(new_n703), .B2(G1996), .ZN(new_n1178));
  AOI22_X1  g753(.A1(new_n1174), .A2(new_n1175), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n814), .B(new_n816), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1179), .B1(new_n1172), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n801), .A2(new_n808), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1182), .B(KEYINPUT107), .Z(new_n1183));
  OAI21_X1  g758(.A(new_n1183), .B1(new_n808), .B2(new_n801), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1181), .B1(new_n1176), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1171), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1172), .B1(new_n704), .B2(new_n1177), .ZN(new_n1187));
  OR3_X1    g762(.A1(new_n1172), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1188));
  OAI21_X1  g763(.A(KEYINPUT46), .B1(new_n1172), .B2(G1996), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1187), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  XOR2_X1   g765(.A(new_n1190), .B(KEYINPUT47), .Z(new_n1191));
  NOR2_X1   g766(.A1(new_n1183), .A2(new_n1172), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1192), .B(KEYINPUT48), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1191), .B1(new_n1193), .B2(new_n1181), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n756), .A2(G2067), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n814), .A2(new_n817), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n1196), .B(KEYINPUT126), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1195), .B1(new_n1179), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT127), .ZN(new_n1199));
  OR2_X1    g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1172), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1194), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1186), .A2(new_n1202), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g778(.A1(new_n460), .A2(G227), .ZN(new_n1205));
  NAND3_X1  g779(.A1(new_n693), .A2(new_n659), .A3(new_n1205), .ZN(new_n1206));
  NOR2_X1   g780(.A1(new_n958), .A2(new_n959), .ZN(new_n1207));
  NOR3_X1   g781(.A1(new_n1206), .A2(new_n869), .A3(new_n1207), .ZN(G308));
  OR3_X1    g782(.A1(new_n1206), .A2(new_n869), .A3(new_n1207), .ZN(G225));
endmodule


