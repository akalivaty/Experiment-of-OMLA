//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n554, new_n555, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT66), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT67), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n459), .A2(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n462), .A2(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT68), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n462), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n468), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n466), .B1(new_n472), .B2(G2105), .ZN(G160));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n459), .ZN(new_n475));
  NAND2_X1  g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n463), .B1(new_n475), .B2(new_n476), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  NAND3_X1  g059(.A1(new_n462), .A2(G126), .A3(G2105), .ZN(new_n485));
  OR2_X1    g060(.A1(G102), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n476), .ZN(new_n489));
  NOR2_X1   g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  OAI211_X1 g065(.A(G138), .B(new_n463), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n477), .A2(new_n493), .A3(G138), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n488), .B1(new_n492), .B2(new_n494), .ZN(G164));
  NAND2_X1  g070(.A1(G75), .A2(G543), .ZN(new_n496));
  AND2_X1   g071(.A1(KEYINPUT5), .A2(G543), .ZN(new_n497));
  NOR2_X1   g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G62), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n496), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G651), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(new_n508), .A3(G88), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n508), .A2(G50), .A3(G543), .ZN(new_n510));
  AND3_X1   g085(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT69), .ZN(new_n511));
  AOI21_X1  g086(.A(KEYINPUT69), .B1(new_n509), .B2(new_n510), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n502), .B1(new_n511), .B2(new_n512), .ZN(G303));
  INV_X1    g088(.A(G303), .ZN(G166));
  XOR2_X1   g089(.A(KEYINPUT70), .B(KEYINPUT7), .Z(new_n515));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT70), .B(KEYINPUT7), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n518), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n519));
  AND2_X1   g094(.A1(G63), .A2(G651), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n517), .A2(new_n519), .B1(new_n507), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n523), .A2(new_n524), .B1(new_n505), .B2(new_n506), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n504), .B1(new_n523), .B2(new_n524), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n525), .A2(G89), .B1(new_n526), .B2(G51), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n521), .A2(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n530));
  INV_X1    g105(.A(G64), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n531), .B1(new_n505), .B2(new_n506), .ZN(new_n532));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n530), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g110(.A(KEYINPUT71), .B(new_n533), .C1(new_n499), .C2(new_n531), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n535), .A2(G651), .A3(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n525), .A2(G90), .B1(new_n526), .B2(G52), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  AOI22_X1  g115(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G651), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n508), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G43), .ZN(new_n545));
  AND2_X1   g120(.A1(KEYINPUT6), .A2(G651), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n498), .A2(new_n497), .B1(new_n546), .B2(new_n522), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n544), .A2(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n543), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(new_n551));
  XOR2_X1   g126(.A(new_n551), .B(KEYINPUT72), .Z(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  OAI211_X1 g131(.A(G53), .B(G543), .C1(new_n546), .C2(new_n522), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(KEYINPUT9), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n508), .A2(new_n559), .A3(G53), .A4(G543), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n562), .B1(new_n505), .B2(new_n506), .ZN(new_n563));
  AND2_X1   g138(.A1(G78), .A2(G543), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n525), .A2(G91), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n561), .A2(new_n565), .A3(new_n566), .ZN(G299));
  NAND2_X1  g142(.A1(new_n525), .A2(G87), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n526), .A2(G49), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G288));
  AOI22_X1  g146(.A1(new_n525), .A2(G86), .B1(new_n526), .B2(G48), .ZN(new_n572));
  OAI21_X1  g147(.A(G61), .B1(new_n497), .B2(new_n498), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n573), .A2(KEYINPUT73), .B1(G73), .B2(G543), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT73), .ZN(new_n575));
  OAI211_X1 g150(.A(new_n575), .B(G61), .C1(new_n497), .C2(new_n498), .ZN(new_n576));
  AOI211_X1 g151(.A(KEYINPUT74), .B(new_n542), .C1(new_n574), .C2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n573), .A2(KEYINPUT73), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n579), .A2(new_n576), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n578), .B1(new_n581), .B2(G651), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n572), .B1(new_n577), .B2(new_n582), .ZN(G305));
  XNOR2_X1  g158(.A(KEYINPUT75), .B(G85), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n525), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n526), .A2(G47), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OAI211_X1 g162(.A(new_n585), .B(new_n586), .C1(new_n542), .C2(new_n587), .ZN(G290));
  NAND3_X1  g163(.A1(new_n525), .A2(KEYINPUT10), .A3(G92), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n590));
  INV_X1    g165(.A(G92), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n547), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n499), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(G54), .B2(new_n526), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(KEYINPUT76), .B1(new_n598), .B2(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  MUX2_X1   g175(.A(KEYINPUT76), .B(new_n599), .S(new_n600), .Z(G284));
  MUX2_X1   g176(.A(KEYINPUT76), .B(new_n599), .S(new_n600), .Z(G321));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(G299), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G168), .B2(new_n603), .ZN(G280));
  XNOR2_X1  g180(.A(G280), .B(KEYINPUT77), .ZN(G297));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n598), .B1(new_n607), .B2(G860), .ZN(G148));
  OR2_X1    g183(.A1(new_n543), .A2(new_n549), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(new_n603), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n593), .A2(new_n597), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n611), .A2(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n610), .B1(new_n612), .B2(new_n603), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g189(.A1(new_n477), .A2(G135), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n479), .A2(G123), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n463), .A2(G111), .ZN(new_n617));
  OAI21_X1  g192(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n615), .B(new_n616), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(G2096), .Z(new_n620));
  NAND3_X1  g195(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  XOR2_X1   g198(.A(KEYINPUT78), .B(G2100), .Z(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n620), .A2(new_n625), .A3(new_n626), .ZN(G156));
  XNOR2_X1  g202(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  INV_X1    g207(.A(G2430), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n632), .A2(new_n633), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n631), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n632), .A2(new_n633), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n638), .A2(new_n630), .A3(new_n634), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n637), .A2(KEYINPUT14), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(KEYINPUT80), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT80), .ZN(new_n642));
  NAND4_X1  g217(.A1(new_n637), .A2(new_n642), .A3(KEYINPUT14), .A4(new_n639), .ZN(new_n643));
  XOR2_X1   g218(.A(G2443), .B(G2446), .Z(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  AND3_X1   g222(.A1(new_n641), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n647), .B1(new_n641), .B2(new_n643), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n629), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n641), .A2(new_n643), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(new_n646), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n641), .A2(new_n643), .A3(new_n647), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(new_n628), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1341), .B(G1348), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n650), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n656), .A2(G14), .ZN(new_n657));
  INV_X1    g232(.A(KEYINPUT81), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n650), .A2(new_n654), .ZN(new_n659));
  INV_X1    g234(.A(new_n655), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI211_X1 g236(.A(KEYINPUT81), .B(new_n655), .C1(new_n650), .C2(new_n654), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n657), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n665), .B1(new_n668), .B2(KEYINPUT18), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT82), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2100), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT18), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n668), .A2(KEYINPUT17), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n666), .A2(new_n667), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2096), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n671), .B(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(G1991), .B(G1996), .Z(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT84), .B(KEYINPUT20), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1961), .B(G1966), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT83), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1956), .B(G2474), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n683), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1971), .B(G1976), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n680), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT19), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n688), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n681), .B(KEYINPUT83), .ZN(new_n693));
  NAND4_X1  g268(.A1(new_n692), .A2(new_n693), .A3(new_n686), .A4(new_n679), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n683), .A2(new_n684), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n696), .A2(new_n692), .A3(new_n685), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n685), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n698), .A2(new_n689), .A3(new_n687), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n695), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(KEYINPUT85), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT85), .ZN(new_n702));
  NAND4_X1  g277(.A1(new_n695), .A2(new_n702), .A3(new_n697), .A4(new_n699), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n701), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n704), .B1(new_n701), .B2(new_n703), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n678), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n701), .A2(new_n703), .ZN(new_n709));
  INV_X1    g284(.A(new_n704), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n678), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n711), .A2(new_n712), .A3(new_n705), .ZN(new_n713));
  XNOR2_X1  g288(.A(G1981), .B(G1986), .ZN(new_n714));
  AND3_X1   g289(.A1(new_n708), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n714), .B1(new_n708), .B2(new_n713), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(G229));
  XNOR2_X1  g293(.A(KEYINPUT95), .B(KEYINPUT25), .ZN(new_n719));
  AND3_X1   g294(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G139), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(new_n464), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n724), .A2(new_n463), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n727), .B2(G33), .ZN(new_n729));
  INV_X1    g304(.A(G2072), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(G16), .A2(G19), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n550), .B2(G16), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(G1341), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n733), .A2(G1341), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT86), .B(G29), .Z(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G27), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G164), .B2(new_n736), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G2078), .ZN(new_n739));
  NOR4_X1   g314(.A1(new_n731), .A2(new_n734), .A3(new_n735), .A4(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G16), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G20), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT23), .ZN(new_n743));
  INV_X1    g318(.A(G299), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(new_n741), .ZN(new_n745));
  INV_X1    g320(.A(G1956), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n736), .A2(G35), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT100), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G162), .B2(new_n736), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT101), .B(KEYINPUT29), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n740), .B(new_n747), .C1(G2090), .C2(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n729), .A2(new_n730), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT97), .ZN(new_n755));
  NOR2_X1   g330(.A1(G4), .A2(G16), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n598), .B2(G16), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT94), .ZN(new_n758));
  INV_X1    g333(.A(G1348), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n752), .A2(G2090), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n741), .A2(G5), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G171), .B2(new_n741), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT99), .B(G1961), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n755), .A2(new_n760), .A3(new_n761), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n727), .A2(G32), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n477), .A2(G141), .B1(G105), .B2(new_n460), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n479), .A2(G129), .ZN(new_n769));
  NAND3_X1  g344(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT26), .Z(new_n771));
  NAND3_X1  g346(.A1(new_n768), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n767), .B1(new_n773), .B2(new_n727), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT27), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1996), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT30), .B(G28), .ZN(new_n777));
  OR2_X1    g352(.A1(KEYINPUT31), .A2(G11), .ZN(new_n778));
  NAND2_X1  g353(.A1(KEYINPUT31), .A2(G11), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n777), .A2(new_n727), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n619), .B2(new_n736), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT98), .Z(new_n782));
  NAND2_X1  g357(.A1(new_n736), .A2(G26), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT28), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n477), .A2(G140), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n479), .A2(G128), .ZN(new_n786));
  OR2_X1    g361(.A1(G104), .A2(G2105), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n787), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n785), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n784), .B1(new_n790), .B2(new_n727), .ZN(new_n791));
  INV_X1    g366(.A(G2067), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n741), .A2(G21), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G168), .B2(new_n741), .ZN(new_n795));
  INV_X1    g370(.A(G1966), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n776), .A2(new_n782), .A3(new_n793), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(G160), .A2(G29), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT24), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(G34), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(G34), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n736), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT96), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G2084), .ZN(new_n806));
  NOR4_X1   g381(.A1(new_n753), .A2(new_n766), .A3(new_n798), .A4(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n741), .A2(G23), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G288), .B2(G16), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT33), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G1976), .ZN(new_n816));
  INV_X1    g391(.A(G1976), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n813), .A2(new_n817), .A3(new_n814), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n741), .A2(G22), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT91), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G303), .B2(G16), .ZN(new_n823));
  INV_X1    g398(.A(G1971), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n823), .A2(new_n824), .ZN(new_n827));
  OAI21_X1  g402(.A(KEYINPUT92), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n827), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT92), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n829), .A2(new_n830), .A3(new_n825), .ZN(new_n831));
  AND3_X1   g406(.A1(new_n819), .A2(new_n828), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(G305), .A2(G16), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n741), .A2(G6), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(KEYINPUT32), .B(G1981), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(KEYINPUT90), .ZN(new_n838));
  INV_X1    g413(.A(new_n836), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n835), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT90), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n832), .A2(new_n838), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(KEYINPUT34), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT34), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n832), .A2(new_n838), .A3(new_n842), .A4(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT93), .ZN(new_n847));
  INV_X1    g422(.A(G290), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(KEYINPUT88), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT88), .ZN(new_n850));
  NAND2_X1  g425(.A1(G290), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n741), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(G16), .A2(G24), .ZN(new_n853));
  OR3_X1    g428(.A1(new_n852), .A2(KEYINPUT89), .A3(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(G1986), .ZN(new_n855));
  OAI21_X1  g430(.A(KEYINPUT89), .B1(new_n852), .B2(new_n853), .ZN(new_n856));
  AND3_X1   g431(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n855), .B1(new_n854), .B2(new_n856), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n477), .A2(G131), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n479), .A2(G119), .ZN(new_n860));
  OR2_X1    g435(.A1(G95), .A2(G2105), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n861), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT87), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT87), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n859), .A2(new_n860), .A3(new_n865), .A4(new_n862), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n736), .ZN(new_n868));
  MUX2_X1   g443(.A(G25), .B(new_n867), .S(new_n868), .Z(new_n869));
  XOR2_X1   g444(.A(KEYINPUT35), .B(G1991), .Z(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n869), .B(new_n871), .ZN(new_n872));
  NOR3_X1   g447(.A1(new_n857), .A2(new_n858), .A3(new_n872), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n846), .A2(new_n847), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n847), .B1(new_n846), .B2(new_n873), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n844), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT36), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT36), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n878), .B(new_n844), .C1(new_n874), .C2(new_n875), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n808), .B1(new_n877), .B2(new_n879), .ZN(G311));
  NAND2_X1  g455(.A1(new_n877), .A2(new_n879), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n807), .ZN(G150));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n883));
  INV_X1    g458(.A(G67), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(new_n505), .B2(new_n506), .ZN(new_n885));
  NAND2_X1  g460(.A1(G80), .A2(G543), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n883), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  OAI211_X1 g463(.A(KEYINPUT102), .B(new_n886), .C1(new_n499), .C2(new_n884), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(G651), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n891));
  XNOR2_X1  g466(.A(KEYINPUT103), .B(G55), .ZN(new_n892));
  AOI22_X1  g467(.A1(new_n525), .A2(G93), .B1(new_n526), .B2(new_n892), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n891), .B1(new_n890), .B2(new_n893), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n609), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n890), .A2(new_n893), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT104), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n890), .A2(new_n893), .A3(new_n891), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(new_n550), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT38), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n611), .A2(new_n607), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n902), .B(new_n903), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n904), .A2(KEYINPUT39), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(KEYINPUT39), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n905), .A2(new_n906), .A3(G860), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n897), .A2(G860), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT37), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n907), .A2(new_n909), .ZN(G145));
  XNOR2_X1  g485(.A(G160), .B(new_n619), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(G162), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT106), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n479), .A2(G130), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n477), .A2(G142), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n917), .B1(new_n463), .B2(G118), .ZN(new_n918));
  INV_X1    g493(.A(G118), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n919), .A2(KEYINPUT105), .A3(G2105), .ZN(new_n920));
  OR2_X1    g495(.A1(G106), .A2(G2105), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n918), .A2(new_n920), .A3(new_n921), .A4(G2104), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n915), .A2(new_n916), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n622), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n622), .A2(new_n915), .A3(new_n916), .A4(new_n922), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n925), .A2(new_n864), .A3(new_n866), .A4(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n925), .A2(new_n926), .B1(new_n864), .B2(new_n866), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n914), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n925), .A2(new_n926), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n867), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n932), .A2(KEYINPUT106), .A3(new_n927), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n723), .A2(new_n725), .ZN(new_n935));
  INV_X1    g510(.A(new_n488), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n494), .A2(new_n492), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n938), .A2(new_n789), .ZN(new_n939));
  NOR2_X1   g514(.A1(G164), .A2(new_n790), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n935), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n938), .A2(new_n789), .ZN(new_n942));
  NAND2_X1  g517(.A1(G164), .A2(new_n790), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n726), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n941), .A2(new_n772), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n941), .A2(new_n944), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n773), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n934), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n941), .A2(new_n772), .A3(new_n944), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n772), .B1(new_n941), .B2(new_n944), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n949), .A2(new_n950), .A3(new_n930), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n913), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G37), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n930), .B(new_n933), .C1(new_n949), .C2(new_n950), .ZN(new_n955));
  INV_X1    g530(.A(new_n930), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n947), .A2(new_n956), .A3(new_n945), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n955), .A2(new_n912), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT107), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n955), .A2(new_n960), .A3(new_n957), .A4(new_n912), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n954), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n963), .B(new_n964), .ZN(G395));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n581), .A2(G651), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT74), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n542), .B1(new_n574), .B2(new_n576), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n578), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(G290), .B1(new_n971), .B2(new_n572), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n572), .B(G290), .C1(new_n577), .C2(new_n582), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G288), .ZN(new_n975));
  NAND2_X1  g550(.A1(G303), .A2(new_n975), .ZN(new_n976));
  OAI211_X1 g551(.A(G288), .B(new_n502), .C1(new_n511), .C2(new_n512), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n972), .A2(new_n974), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(G305), .A2(new_n848), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n980), .A2(new_n973), .B1(new_n977), .B2(new_n976), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n966), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n978), .B1(new_n972), .B2(new_n974), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n980), .A2(new_n977), .A3(new_n976), .A4(new_n973), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n983), .A2(KEYINPUT110), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT42), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n979), .A2(new_n981), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n987), .B1(KEYINPUT42), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n901), .B(new_n612), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n561), .A2(KEYINPUT109), .A3(new_n565), .A4(new_n566), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n991), .A2(new_n593), .A3(new_n597), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n566), .A2(new_n565), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT109), .B1(new_n993), .B2(new_n561), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT109), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n611), .A2(G299), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n990), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(G299), .A2(new_n996), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n598), .A2(new_n1001), .A3(new_n991), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT41), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n1002), .A2(new_n1003), .A3(new_n997), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1003), .B1(new_n1002), .B2(new_n997), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1000), .B1(new_n990), .B2(new_n1006), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n989), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n989), .A2(new_n1007), .ZN(new_n1009));
  OAI21_X1  g584(.A(G868), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n897), .A2(new_n603), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(G295));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1011), .ZN(G331));
  AND4_X1   g588(.A1(new_n521), .A2(new_n537), .A3(new_n527), .A4(new_n538), .ZN(new_n1014));
  AOI22_X1  g589(.A1(new_n537), .A2(new_n538), .B1(new_n521), .B2(new_n527), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n1016), .A2(new_n896), .A3(new_n900), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1015), .ZN(new_n1018));
  NAND2_X1  g593(.A1(G171), .A2(G168), .ZN(new_n1019));
  AOI22_X1  g594(.A1(new_n896), .A2(new_n900), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI22_X1  g595(.A1(new_n1017), .A2(new_n1020), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1018), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n894), .A2(new_n895), .A3(new_n609), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n550), .B1(new_n898), .B2(new_n899), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1022), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1016), .A2(new_n896), .A3(new_n900), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n999), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1021), .A2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n986), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(G37), .B1(new_n986), .B2(new_n1028), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1029), .B1(new_n1030), .B2(KEYINPUT111), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n985), .A2(new_n982), .B1(new_n1021), .B2(new_n1027), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1032), .B1(new_n1033), .B2(G37), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT43), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n953), .B1(new_n986), .B2(new_n1028), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT43), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT41), .B1(new_n995), .B2(new_n998), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1002), .A2(new_n1003), .A3(new_n997), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1004), .A2(KEYINPUT112), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1038), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n1044), .A2(new_n1027), .B1(new_n982), .B2(new_n985), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n1036), .A2(new_n1037), .A3(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT44), .B1(new_n1035), .B2(new_n1046), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n1036), .A2(KEYINPUT43), .A3(new_n1045), .ZN(new_n1048));
  INV_X1    g623(.A(new_n985), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT110), .B1(new_n983), .B2(new_n984), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1025), .A2(new_n999), .A3(new_n1026), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1025), .A2(new_n1026), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1052));
  OAI22_X1  g627(.A1(new_n1049), .A2(new_n1050), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1053), .A2(KEYINPUT111), .A3(new_n953), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1029), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1034), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1048), .B1(new_n1056), .B2(KEYINPUT43), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1047), .B1(KEYINPUT44), .B2(new_n1057), .ZN(G397));
  NAND2_X1  g633(.A1(new_n472), .A2(G2105), .ZN(new_n1059));
  INV_X1    g634(.A(new_n466), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(G40), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G1384), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n938), .A2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT116), .B(G8), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n975), .A2(new_n817), .ZN(new_n1067));
  XNOR2_X1  g642(.A(new_n1067), .B(KEYINPUT117), .ZN(new_n1068));
  INV_X1    g643(.A(G1981), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1069), .B(new_n572), .C1(new_n577), .C2(new_n582), .ZN(new_n1070));
  INV_X1    g645(.A(new_n572), .ZN(new_n1071));
  OAI21_X1  g646(.A(G1981), .B1(new_n1071), .B2(new_n969), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT49), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1070), .A2(KEYINPUT49), .A3(new_n1072), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1068), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1070), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1066), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(G1384), .B1(new_n936), .B2(new_n937), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT113), .B1(new_n1080), .B2(KEYINPUT45), .ZN(new_n1081));
  INV_X1    g656(.A(G40), .ZN(new_n1082));
  AOI211_X1 g657(.A(new_n1082), .B(new_n466), .C1(new_n472), .C2(G2105), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT45), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1084), .B(new_n1085), .C1(G164), .C2(G1384), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n938), .A2(KEYINPUT45), .A3(new_n1062), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1081), .A2(new_n1083), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT114), .B(G1971), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT50), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n938), .A2(new_n1092), .A3(new_n1062), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1083), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT115), .B(G2090), .Z(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1090), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(G303), .A2(G8), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1098), .B(KEYINPUT55), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1097), .A2(G8), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1075), .A2(new_n1066), .A3(new_n1076), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n975), .A2(G1976), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT52), .B1(G288), .B2(new_n817), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1066), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1083), .A2(new_n1080), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1065), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(new_n1107), .A3(new_n1103), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT52), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1102), .A2(new_n1105), .A3(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1079), .B1(new_n1101), .B2(new_n1110), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1102), .A2(new_n1105), .A3(new_n1109), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1088), .A2(new_n1089), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1099), .B1(new_n1113), .B2(new_n1065), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT53), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n1088), .B2(G2078), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1085), .B1(G164), .B2(G1384), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1083), .A2(new_n1117), .A3(new_n1087), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1115), .A2(G2078), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1083), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1120));
  INV_X1    g695(.A(G1961), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1118), .A2(new_n1119), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(G301), .B1(new_n1116), .B2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1112), .A2(new_n1114), .A3(new_n1101), .A4(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G8), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1083), .A2(new_n1117), .A3(new_n1087), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n796), .ZN(new_n1127));
  INV_X1    g702(.A(G2084), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1083), .A2(new_n1091), .A3(new_n1093), .A4(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1125), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(G168), .A2(new_n1065), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT51), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1065), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1131), .A2(KEYINPUT51), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT123), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1094), .A2(new_n1128), .B1(new_n1126), .B2(new_n796), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1137), .B(new_n1134), .C1(new_n1138), .C2(new_n1065), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1132), .A2(new_n1136), .A3(new_n1139), .ZN(new_n1140));
  OR3_X1    g715(.A1(new_n1138), .A2(G168), .A3(new_n1065), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1124), .B1(new_n1142), .B2(KEYINPUT62), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1140), .A2(new_n1144), .A3(new_n1141), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1111), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1113), .A2(new_n1125), .A3(new_n1099), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1147), .A2(new_n1110), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1138), .A2(G286), .A3(new_n1065), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1148), .A2(KEYINPUT118), .A3(new_n1114), .A4(new_n1149), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1112), .A2(new_n1114), .A3(new_n1101), .A4(new_n1149), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT118), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT63), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1150), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1097), .A2(G8), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1154), .B1(new_n1156), .B2(new_n1099), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1148), .A2(new_n1149), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  NOR3_X1   g734(.A1(G164), .A2(new_n1085), .A3(G1384), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1160), .A2(new_n1061), .ZN(new_n1161));
  XNOR2_X1  g736(.A(KEYINPUT56), .B(G2072), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT120), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1161), .A2(new_n1086), .A3(new_n1081), .A4(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n993), .A2(KEYINPUT119), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT57), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(new_n744), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1120), .A2(new_n746), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1164), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1168), .B1(new_n1164), .B2(new_n1169), .ZN(new_n1171));
  AOI22_X1  g746(.A1(new_n759), .A2(new_n1120), .B1(new_n1064), .B2(new_n792), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1172), .A2(new_n611), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1170), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n598), .B1(new_n1172), .B2(KEYINPUT60), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT122), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1176), .B1(new_n1172), .B2(KEYINPUT60), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1120), .A2(new_n759), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1064), .A2(new_n792), .ZN(new_n1179));
  AND4_X1   g754(.A1(new_n1176), .A2(new_n1178), .A3(KEYINPUT60), .A4(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1175), .B1(new_n1177), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT60), .ZN(new_n1183));
  OAI21_X1  g758(.A(KEYINPUT122), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n611), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1172), .A2(new_n1176), .A3(KEYINPUT60), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1164), .A2(new_n1169), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1168), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1190), .A2(KEYINPUT61), .A3(new_n1170), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1181), .A2(new_n1187), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n1193));
  AND3_X1   g768(.A1(new_n1164), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1193), .B1(new_n1194), .B2(new_n1171), .ZN(new_n1195));
  XOR2_X1   g770(.A(KEYINPUT58), .B(G1341), .Z(new_n1196));
  OAI21_X1  g771(.A(new_n1196), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT121), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1106), .A2(KEYINPUT121), .A3(new_n1196), .ZN(new_n1200));
  OAI211_X1 g775(.A(new_n1199), .B(new_n1200), .C1(G1996), .C2(new_n1088), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n550), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT59), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1201), .A2(KEYINPUT59), .A3(new_n550), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1195), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1174), .B1(new_n1192), .B2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1112), .A2(new_n1114), .A3(new_n1101), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1208), .B1(new_n1141), .B2(new_n1140), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1116), .A2(new_n1122), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1210), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1211));
  NAND4_X1  g786(.A1(new_n1116), .A2(new_n1122), .A3(KEYINPUT124), .A4(G301), .ZN(new_n1212));
  AND3_X1   g787(.A1(new_n1211), .A2(KEYINPUT54), .A3(new_n1212), .ZN(new_n1213));
  AOI21_X1  g788(.A(KEYINPUT54), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1214));
  NOR2_X1   g789(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1207), .A2(new_n1209), .A3(new_n1215), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1146), .A2(new_n1159), .A3(new_n1216), .ZN(new_n1217));
  NOR2_X1   g792(.A1(new_n1117), .A2(new_n1061), .ZN(new_n1218));
  INV_X1    g793(.A(G1996), .ZN(new_n1219));
  XNOR2_X1  g794(.A(new_n772), .B(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g795(.A(new_n789), .B(new_n792), .ZN(new_n1221));
  AND2_X1   g796(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n867), .A2(new_n871), .ZN(new_n1223));
  NOR2_X1   g798(.A1(new_n867), .A2(new_n871), .ZN(new_n1224));
  INV_X1    g799(.A(new_n1224), .ZN(new_n1225));
  NAND3_X1  g800(.A1(new_n1222), .A2(new_n1223), .A3(new_n1225), .ZN(new_n1226));
  XNOR2_X1  g801(.A(G290), .B(G1986), .ZN(new_n1227));
  OAI21_X1  g802(.A(new_n1218), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1217), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g804(.A1(new_n1218), .A2(new_n855), .A3(new_n848), .ZN(new_n1230));
  INV_X1    g805(.A(new_n1230), .ZN(new_n1231));
  NOR2_X1   g806(.A1(new_n1231), .A2(KEYINPUT48), .ZN(new_n1232));
  AND2_X1   g807(.A1(new_n1231), .A2(KEYINPUT48), .ZN(new_n1233));
  AOI211_X1 g808(.A(new_n1232), .B(new_n1233), .C1(new_n1218), .C2(new_n1226), .ZN(new_n1234));
  AOI21_X1  g809(.A(KEYINPUT46), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1235));
  INV_X1    g810(.A(KEYINPUT126), .ZN(new_n1236));
  AND2_X1   g811(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NOR2_X1   g812(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1238));
  INV_X1    g813(.A(new_n1218), .ZN(new_n1239));
  AOI21_X1  g814(.A(new_n772), .B1(KEYINPUT46), .B2(new_n1219), .ZN(new_n1240));
  AND2_X1   g815(.A1(new_n1221), .A2(new_n1240), .ZN(new_n1241));
  OAI22_X1  g816(.A1(new_n1237), .A2(new_n1238), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1242));
  XOR2_X1   g817(.A(new_n1242), .B(KEYINPUT47), .Z(new_n1243));
  INV_X1    g818(.A(KEYINPUT125), .ZN(new_n1244));
  OAI21_X1  g819(.A(new_n1222), .B1(new_n1244), .B2(new_n1224), .ZN(new_n1245));
  NOR2_X1   g820(.A1(new_n1225), .A2(KEYINPUT125), .ZN(new_n1246));
  OAI22_X1  g821(.A1(new_n1245), .A2(new_n1246), .B1(G2067), .B2(new_n789), .ZN(new_n1247));
  AOI211_X1 g822(.A(new_n1234), .B(new_n1243), .C1(new_n1218), .C2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g823(.A1(new_n1229), .A2(new_n1248), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g824(.A(KEYINPUT127), .ZN(new_n1251));
  NOR2_X1   g825(.A1(G227), .A2(new_n457), .ZN(new_n1252));
  AND2_X1   g826(.A1(new_n663), .A2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g827(.A1(new_n963), .A2(new_n717), .A3(new_n1253), .ZN(new_n1254));
  OAI21_X1  g828(.A(new_n1251), .B1(new_n1057), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g829(.A1(new_n952), .A2(new_n953), .ZN(new_n1256));
  AOI21_X1  g830(.A(new_n1256), .B1(new_n959), .B2(new_n961), .ZN(new_n1257));
  OAI211_X1 g831(.A(new_n663), .B(new_n1252), .C1(new_n715), .C2(new_n716), .ZN(new_n1258));
  NOR2_X1   g832(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g833(.A(new_n1037), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1260));
  OAI211_X1 g834(.A(new_n1259), .B(KEYINPUT127), .C1(new_n1260), .C2(new_n1048), .ZN(new_n1261));
  AND2_X1   g835(.A1(new_n1255), .A2(new_n1261), .ZN(G308));
  NAND2_X1  g836(.A1(new_n1255), .A2(new_n1261), .ZN(G225));
endmodule


