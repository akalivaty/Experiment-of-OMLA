

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580;

  NOR2_X1 U321 ( .A1(n478), .A2(n452), .ZN(n444) );
  XOR2_X1 U322 ( .A(KEYINPUT119), .B(KEYINPUT55), .Z(n289) );
  XOR2_X1 U323 ( .A(n323), .B(G176GAT), .Z(n290) );
  XOR2_X1 U324 ( .A(n344), .B(KEYINPUT32), .Z(n291) );
  XNOR2_X1 U325 ( .A(G85GAT), .B(KEYINPUT70), .ZN(n302) );
  NOR2_X1 U326 ( .A1(n534), .A2(n448), .ZN(n449) );
  INV_X1 U327 ( .A(KEYINPUT47), .ZN(n372) );
  XNOR2_X1 U328 ( .A(n372), .B(KEYINPUT107), .ZN(n373) );
  XNOR2_X1 U329 ( .A(n374), .B(n373), .ZN(n380) );
  XNOR2_X1 U330 ( .A(n381), .B(KEYINPUT48), .ZN(n382) );
  NOR2_X1 U331 ( .A1(n456), .A2(n455), .ZN(n468) );
  XNOR2_X1 U332 ( .A(n383), .B(n382), .ZN(n516) );
  XNOR2_X1 U333 ( .A(n355), .B(n354), .ZN(n568) );
  INV_X1 U334 ( .A(G190GAT), .ZN(n438) );
  XNOR2_X1 U335 ( .A(n568), .B(KEYINPUT41), .ZN(n550) );
  INV_X1 U336 ( .A(G43GAT), .ZN(n461) );
  XNOR2_X1 U337 ( .A(KEYINPUT38), .B(n460), .ZN(n490) );
  XNOR2_X1 U338 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U339 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U340 ( .A(n441), .B(n440), .ZN(G1351GAT) );
  XNOR2_X1 U341 ( .A(n464), .B(n463), .ZN(G1330GAT) );
  XNOR2_X1 U342 ( .A(G43GAT), .B(G50GAT), .ZN(n292) );
  XNOR2_X1 U343 ( .A(n292), .B(KEYINPUT8), .ZN(n293) );
  XOR2_X1 U344 ( .A(n293), .B(KEYINPUT7), .Z(n295) );
  XNOR2_X1 U345 ( .A(G29GAT), .B(G36GAT), .ZN(n294) );
  XOR2_X1 U346 ( .A(n295), .B(n294), .Z(n366) );
  XOR2_X1 U347 ( .A(KEYINPUT9), .B(KEYINPUT65), .Z(n297) );
  XNOR2_X1 U348 ( .A(G134GAT), .B(KEYINPUT10), .ZN(n296) );
  XNOR2_X1 U349 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U350 ( .A(n366), .B(n298), .Z(n309) );
  XOR2_X1 U351 ( .A(G92GAT), .B(G106GAT), .Z(n300) );
  XOR2_X1 U352 ( .A(G162GAT), .B(KEYINPUT73), .Z(n409) );
  XOR2_X1 U353 ( .A(G218GAT), .B(G190GAT), .Z(n393) );
  XNOR2_X1 U354 ( .A(n409), .B(n393), .ZN(n299) );
  XNOR2_X1 U355 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U356 ( .A(n301), .B(KEYINPUT11), .Z(n307) );
  XNOR2_X1 U357 ( .A(n302), .B(G99GAT), .ZN(n344) );
  XOR2_X1 U358 ( .A(n344), .B(KEYINPUT74), .Z(n304) );
  NAND2_X1 U359 ( .A1(G232GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U360 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U361 ( .A(n305), .B(KEYINPUT75), .ZN(n306) );
  XNOR2_X1 U362 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U363 ( .A(n309), .B(n308), .Z(n528) );
  XOR2_X1 U364 ( .A(G190GAT), .B(G43GAT), .Z(n311) );
  NAND2_X1 U365 ( .A1(G227GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U366 ( .A(n311), .B(n310), .ZN(n314) );
  XOR2_X1 U367 ( .A(G169GAT), .B(KEYINPUT19), .Z(n313) );
  XNOR2_X1 U368 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n313), .B(n312), .ZN(n386) );
  XOR2_X1 U370 ( .A(n314), .B(n386), .Z(n322) );
  XOR2_X1 U371 ( .A(KEYINPUT81), .B(KEYINPUT79), .Z(n316) );
  XNOR2_X1 U372 ( .A(G99GAT), .B(KEYINPUT20), .ZN(n315) );
  XNOR2_X1 U373 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U374 ( .A(KEYINPUT80), .B(G183GAT), .Z(n318) );
  XNOR2_X1 U375 ( .A(G71GAT), .B(G15GAT), .ZN(n317) );
  XNOR2_X1 U376 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U377 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U378 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U379 ( .A(G113GAT), .B(G120GAT), .Z(n325) );
  XNOR2_X1 U380 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n325), .B(n324), .ZN(n422) );
  XNOR2_X1 U382 ( .A(n422), .B(G127GAT), .ZN(n326) );
  XOR2_X1 U383 ( .A(n290), .B(n326), .Z(n519) );
  INV_X1 U384 ( .A(n519), .ZN(n478) );
  XOR2_X1 U385 ( .A(G78GAT), .B(G71GAT), .Z(n328) );
  XNOR2_X1 U386 ( .A(KEYINPUT13), .B(KEYINPUT68), .ZN(n327) );
  XNOR2_X1 U387 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U388 ( .A(G57GAT), .B(n329), .ZN(n354) );
  XOR2_X1 U389 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n331) );
  XNOR2_X1 U390 ( .A(G64GAT), .B(KEYINPUT76), .ZN(n330) );
  XNOR2_X1 U391 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U392 ( .A(n354), .B(n332), .Z(n341) );
  XOR2_X1 U393 ( .A(G127GAT), .B(G155GAT), .Z(n419) );
  XNOR2_X1 U394 ( .A(G183GAT), .B(G211GAT), .ZN(n333) );
  XNOR2_X1 U395 ( .A(n333), .B(G8GAT), .ZN(n388) );
  XOR2_X1 U396 ( .A(n419), .B(n388), .Z(n335) );
  NAND2_X1 U397 ( .A1(G231GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U398 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U399 ( .A(n336), .B(KEYINPUT77), .Z(n339) );
  XNOR2_X1 U400 ( .A(G1GAT), .B(G15GAT), .ZN(n337) );
  XNOR2_X1 U401 ( .A(n337), .B(G22GAT), .ZN(n361) );
  XNOR2_X1 U402 ( .A(n361), .B(KEYINPUT14), .ZN(n338) );
  XNOR2_X1 U403 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U404 ( .A(n341), .B(n340), .ZN(n572) );
  XNOR2_X1 U405 ( .A(n572), .B(KEYINPUT105), .ZN(n557) );
  XOR2_X1 U406 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n343) );
  XNOR2_X1 U407 ( .A(G120GAT), .B(KEYINPUT72), .ZN(n342) );
  XNOR2_X1 U408 ( .A(n343), .B(n342), .ZN(n347) );
  NAND2_X1 U409 ( .A1(G230GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U410 ( .A(n291), .B(n345), .ZN(n346) );
  XOR2_X1 U411 ( .A(n347), .B(n346), .Z(n353) );
  XOR2_X1 U412 ( .A(KEYINPUT71), .B(G204GAT), .Z(n349) );
  XNOR2_X1 U413 ( .A(G92GAT), .B(G176GAT), .ZN(n348) );
  XNOR2_X1 U414 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U415 ( .A(G64GAT), .B(n350), .Z(n392) );
  XNOR2_X1 U416 ( .A(G148GAT), .B(G106GAT), .ZN(n351) );
  XNOR2_X1 U417 ( .A(n351), .B(KEYINPUT69), .ZN(n402) );
  XNOR2_X1 U418 ( .A(n392), .B(n402), .ZN(n352) );
  XNOR2_X1 U419 ( .A(n353), .B(n352), .ZN(n355) );
  INV_X1 U420 ( .A(n550), .ZN(n537) );
  XOR2_X1 U421 ( .A(G169GAT), .B(G113GAT), .Z(n357) );
  NAND2_X1 U422 ( .A1(G229GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U423 ( .A(n357), .B(n356), .ZN(n365) );
  XOR2_X1 U424 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n363) );
  XOR2_X1 U425 ( .A(KEYINPUT29), .B(G197GAT), .Z(n359) );
  XNOR2_X1 U426 ( .A(G141GAT), .B(G8GAT), .ZN(n358) );
  XNOR2_X1 U427 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U428 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U429 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n365), .B(n364), .ZN(n367) );
  XNOR2_X1 U431 ( .A(n367), .B(n366), .ZN(n563) );
  NAND2_X1 U432 ( .A1(n537), .A2(n563), .ZN(n369) );
  XOR2_X1 U433 ( .A(KEYINPUT106), .B(KEYINPUT46), .Z(n368) );
  XNOR2_X1 U434 ( .A(n369), .B(n368), .ZN(n370) );
  INV_X1 U435 ( .A(n528), .ZN(n544) );
  NOR2_X1 U436 ( .A1(n370), .A2(n544), .ZN(n371) );
  NAND2_X1 U437 ( .A1(n557), .A2(n371), .ZN(n374) );
  XNOR2_X1 U438 ( .A(KEYINPUT67), .B(n563), .ZN(n548) );
  XOR2_X1 U439 ( .A(KEYINPUT45), .B(KEYINPUT108), .Z(n376) );
  XOR2_X1 U440 ( .A(KEYINPUT36), .B(n528), .Z(n576) );
  NAND2_X1 U441 ( .A1(n572), .A2(n576), .ZN(n375) );
  XNOR2_X1 U442 ( .A(n376), .B(n375), .ZN(n377) );
  NAND2_X1 U443 ( .A1(n548), .A2(n377), .ZN(n378) );
  NOR2_X1 U444 ( .A1(n568), .A2(n378), .ZN(n379) );
  NOR2_X1 U445 ( .A1(n380), .A2(n379), .ZN(n383) );
  XOR2_X1 U446 ( .A(KEYINPUT64), .B(KEYINPUT109), .Z(n381) );
  XOR2_X1 U447 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n385) );
  NAND2_X1 U448 ( .A1(G226GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n385), .B(n384), .ZN(n387) );
  XOR2_X1 U450 ( .A(n387), .B(n386), .Z(n390) );
  XNOR2_X1 U451 ( .A(G36GAT), .B(n388), .ZN(n389) );
  XNOR2_X1 U452 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U453 ( .A(KEYINPUT21), .B(G197GAT), .Z(n408) );
  XOR2_X1 U454 ( .A(n391), .B(n408), .Z(n395) );
  XNOR2_X1 U455 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U456 ( .A(n395), .B(n394), .Z(n507) );
  NOR2_X1 U457 ( .A1(n516), .A2(n507), .ZN(n397) );
  XNOR2_X1 U458 ( .A(KEYINPUT118), .B(KEYINPUT54), .ZN(n396) );
  XNOR2_X1 U459 ( .A(n397), .B(n396), .ZN(n560) );
  XOR2_X1 U460 ( .A(KEYINPUT82), .B(KEYINPUT22), .Z(n399) );
  XNOR2_X1 U461 ( .A(G78GAT), .B(G22GAT), .ZN(n398) );
  XNOR2_X1 U462 ( .A(n399), .B(n398), .ZN(n417) );
  XOR2_X1 U463 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n401) );
  NAND2_X1 U464 ( .A1(G228GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U465 ( .A(n401), .B(n400), .ZN(n403) );
  XOR2_X1 U466 ( .A(n403), .B(n402), .Z(n407) );
  XOR2_X1 U467 ( .A(G141GAT), .B(KEYINPUT2), .Z(n405) );
  XNOR2_X1 U468 ( .A(KEYINPUT3), .B(KEYINPUT83), .ZN(n404) );
  XNOR2_X1 U469 ( .A(n405), .B(n404), .ZN(n418) );
  XNOR2_X1 U470 ( .A(n418), .B(G211GAT), .ZN(n406) );
  XNOR2_X1 U471 ( .A(n407), .B(n406), .ZN(n413) );
  XOR2_X1 U472 ( .A(n408), .B(G218GAT), .Z(n411) );
  XNOR2_X1 U473 ( .A(G50GAT), .B(n409), .ZN(n410) );
  XNOR2_X1 U474 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U475 ( .A(n413), .B(n412), .Z(n415) );
  XNOR2_X1 U476 ( .A(G155GAT), .B(G204GAT), .ZN(n414) );
  XNOR2_X1 U477 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U478 ( .A(n417), .B(n416), .Z(n443) );
  XOR2_X1 U479 ( .A(n419), .B(n418), .Z(n421) );
  XNOR2_X1 U480 ( .A(G29GAT), .B(G162GAT), .ZN(n420) );
  XNOR2_X1 U481 ( .A(n421), .B(n420), .ZN(n426) );
  XOR2_X1 U482 ( .A(n422), .B(G1GAT), .Z(n424) );
  NAND2_X1 U483 ( .A1(G225GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U484 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U485 ( .A(n426), .B(n425), .Z(n434) );
  XOR2_X1 U486 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n428) );
  XNOR2_X1 U487 ( .A(G85GAT), .B(G148GAT), .ZN(n427) );
  XNOR2_X1 U488 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U489 ( .A(G57GAT), .B(KEYINPUT84), .Z(n430) );
  XNOR2_X1 U490 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n429) );
  XNOR2_X1 U491 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U492 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U493 ( .A(n434), .B(n433), .Z(n472) );
  NOR2_X1 U494 ( .A1(n443), .A2(n472), .ZN(n435) );
  NAND2_X1 U495 ( .A1(n560), .A2(n435), .ZN(n436) );
  XNOR2_X1 U496 ( .A(n436), .B(n289), .ZN(n437) );
  NAND2_X1 U497 ( .A1(n478), .A2(n437), .ZN(n556) );
  NOR2_X1 U498 ( .A1(n528), .A2(n556), .ZN(n441) );
  XNOR2_X1 U499 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n439) );
  XOR2_X1 U500 ( .A(n507), .B(KEYINPUT87), .Z(n442) );
  XNOR2_X1 U501 ( .A(n442), .B(KEYINPUT27), .ZN(n453) );
  INV_X1 U502 ( .A(n443), .ZN(n452) );
  XOR2_X1 U503 ( .A(KEYINPUT26), .B(n444), .Z(n562) );
  NOR2_X1 U504 ( .A1(n453), .A2(n562), .ZN(n534) );
  INV_X1 U505 ( .A(n507), .ZN(n475) );
  NAND2_X1 U506 ( .A1(n475), .A2(n478), .ZN(n445) );
  NAND2_X1 U507 ( .A1(n445), .A2(n452), .ZN(n446) );
  XNOR2_X1 U508 ( .A(n446), .B(KEYINPUT25), .ZN(n447) );
  XNOR2_X1 U509 ( .A(n447), .B(KEYINPUT88), .ZN(n448) );
  XNOR2_X1 U510 ( .A(KEYINPUT89), .B(n449), .ZN(n450) );
  INV_X1 U511 ( .A(n472), .ZN(n559) );
  NAND2_X1 U512 ( .A1(n450), .A2(n559), .ZN(n451) );
  XOR2_X1 U513 ( .A(KEYINPUT90), .B(n451), .Z(n456) );
  XOR2_X1 U514 ( .A(n452), .B(KEYINPUT28), .Z(n489) );
  NOR2_X1 U515 ( .A1(n453), .A2(n489), .ZN(n517) );
  NAND2_X1 U516 ( .A1(n517), .A2(n472), .ZN(n454) );
  NOR2_X1 U517 ( .A1(n478), .A2(n454), .ZN(n455) );
  NOR2_X1 U518 ( .A1(n572), .A2(n468), .ZN(n457) );
  XNOR2_X1 U519 ( .A(KEYINPUT96), .B(n457), .ZN(n458) );
  NAND2_X1 U520 ( .A1(n458), .A2(n576), .ZN(n459) );
  XNOR2_X1 U521 ( .A(n459), .B(KEYINPUT37), .ZN(n505) );
  NOR2_X1 U522 ( .A1(n568), .A2(n548), .ZN(n470) );
  NAND2_X1 U523 ( .A1(n505), .A2(n470), .ZN(n460) );
  NOR2_X1 U524 ( .A1(n490), .A2(n519), .ZN(n464) );
  XNOR2_X1 U525 ( .A(KEYINPUT98), .B(KEYINPUT40), .ZN(n462) );
  NAND2_X1 U526 ( .A1(n528), .A2(n572), .ZN(n465) );
  XNOR2_X1 U527 ( .A(n465), .B(KEYINPUT16), .ZN(n466) );
  XNOR2_X1 U528 ( .A(n466), .B(KEYINPUT78), .ZN(n467) );
  NOR2_X1 U529 ( .A1(n468), .A2(n467), .ZN(n469) );
  XOR2_X1 U530 ( .A(KEYINPUT91), .B(n469), .Z(n493) );
  NAND2_X1 U531 ( .A1(n470), .A2(n493), .ZN(n471) );
  XOR2_X1 U532 ( .A(KEYINPUT92), .B(n471), .Z(n482) );
  NAND2_X1 U533 ( .A1(n482), .A2(n472), .ZN(n473) );
  XNOR2_X1 U534 ( .A(n473), .B(KEYINPUT34), .ZN(n474) );
  XNOR2_X1 U535 ( .A(G1GAT), .B(n474), .ZN(G1324GAT) );
  XOR2_X1 U536 ( .A(G8GAT), .B(KEYINPUT93), .Z(n477) );
  NAND2_X1 U537 ( .A1(n475), .A2(n482), .ZN(n476) );
  XNOR2_X1 U538 ( .A(n477), .B(n476), .ZN(G1325GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT94), .B(KEYINPUT35), .Z(n480) );
  NAND2_X1 U540 ( .A1(n478), .A2(n482), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U542 ( .A(G15GAT), .B(n481), .ZN(G1326GAT) );
  XOR2_X1 U543 ( .A(G22GAT), .B(KEYINPUT95), .Z(n484) );
  NAND2_X1 U544 ( .A1(n482), .A2(n489), .ZN(n483) );
  XNOR2_X1 U545 ( .A(n484), .B(n483), .ZN(G1327GAT) );
  NOR2_X1 U546 ( .A1(n559), .A2(n490), .ZN(n487) );
  XOR2_X1 U547 ( .A(G29GAT), .B(KEYINPUT97), .Z(n485) );
  XNOR2_X1 U548 ( .A(KEYINPUT39), .B(n485), .ZN(n486) );
  XNOR2_X1 U549 ( .A(n487), .B(n486), .ZN(G1328GAT) );
  NOR2_X1 U550 ( .A1(n490), .A2(n507), .ZN(n488) );
  XOR2_X1 U551 ( .A(G36GAT), .B(n488), .Z(G1329GAT) );
  XNOR2_X1 U552 ( .A(G50GAT), .B(KEYINPUT99), .ZN(n492) );
  INV_X1 U553 ( .A(n489), .ZN(n512) );
  NOR2_X1 U554 ( .A1(n512), .A2(n490), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(G1331GAT) );
  NOR2_X1 U556 ( .A1(n563), .A2(n550), .ZN(n504) );
  NAND2_X1 U557 ( .A1(n504), .A2(n493), .ZN(n499) );
  NOR2_X1 U558 ( .A1(n559), .A2(n499), .ZN(n495) );
  XNOR2_X1 U559 ( .A(KEYINPUT100), .B(KEYINPUT42), .ZN(n494) );
  XNOR2_X1 U560 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U561 ( .A(G57GAT), .B(n496), .Z(G1332GAT) );
  NOR2_X1 U562 ( .A1(n507), .A2(n499), .ZN(n497) );
  XOR2_X1 U563 ( .A(G64GAT), .B(n497), .Z(G1333GAT) );
  NOR2_X1 U564 ( .A1(n519), .A2(n499), .ZN(n498) );
  XOR2_X1 U565 ( .A(G71GAT), .B(n498), .Z(G1334GAT) );
  NOR2_X1 U566 ( .A1(n499), .A2(n512), .ZN(n503) );
  XOR2_X1 U567 ( .A(KEYINPUT101), .B(KEYINPUT43), .Z(n501) );
  XNOR2_X1 U568 ( .A(G78GAT), .B(KEYINPUT102), .ZN(n500) );
  XNOR2_X1 U569 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U570 ( .A(n503), .B(n502), .ZN(G1335GAT) );
  NAND2_X1 U571 ( .A1(n505), .A2(n504), .ZN(n511) );
  NOR2_X1 U572 ( .A1(n559), .A2(n511), .ZN(n506) );
  XOR2_X1 U573 ( .A(G85GAT), .B(n506), .Z(G1336GAT) );
  NOR2_X1 U574 ( .A1(n507), .A2(n511), .ZN(n509) );
  XNOR2_X1 U575 ( .A(G92GAT), .B(KEYINPUT103), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(n508), .ZN(G1337GAT) );
  NOR2_X1 U577 ( .A1(n519), .A2(n511), .ZN(n510) );
  XOR2_X1 U578 ( .A(G99GAT), .B(n510), .Z(G1338GAT) );
  NOR2_X1 U579 ( .A1(n512), .A2(n511), .ZN(n514) );
  XNOR2_X1 U580 ( .A(KEYINPUT104), .B(KEYINPUT44), .ZN(n513) );
  XNOR2_X1 U581 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U582 ( .A(G106GAT), .B(n515), .Z(G1339GAT) );
  NOR2_X1 U583 ( .A1(n559), .A2(n516), .ZN(n533) );
  NAND2_X1 U584 ( .A1(n517), .A2(n533), .ZN(n518) );
  NOR2_X1 U585 ( .A1(n519), .A2(n518), .ZN(n520) );
  XOR2_X1 U586 ( .A(KEYINPUT110), .B(n520), .Z(n529) );
  NOR2_X1 U587 ( .A1(n548), .A2(n529), .ZN(n521) );
  XOR2_X1 U588 ( .A(G113GAT), .B(n521), .Z(G1340GAT) );
  NOR2_X1 U589 ( .A1(n529), .A2(n550), .ZN(n523) );
  XNOR2_X1 U590 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n522) );
  XNOR2_X1 U591 ( .A(n523), .B(n522), .ZN(G1341GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT50), .B(KEYINPUT111), .Z(n525) );
  XNOR2_X1 U593 ( .A(G127GAT), .B(KEYINPUT112), .ZN(n524) );
  XNOR2_X1 U594 ( .A(n525), .B(n524), .ZN(n527) );
  NOR2_X1 U595 ( .A1(n529), .A2(n557), .ZN(n526) );
  XOR2_X1 U596 ( .A(n527), .B(n526), .Z(G1342GAT) );
  NOR2_X1 U597 ( .A1(n529), .A2(n528), .ZN(n531) );
  XNOR2_X1 U598 ( .A(KEYINPUT113), .B(KEYINPUT51), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U600 ( .A(G134GAT), .B(n532), .Z(G1343GAT) );
  AND2_X1 U601 ( .A1(n534), .A2(n533), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n545), .A2(n563), .ZN(n535) );
  XNOR2_X1 U603 ( .A(KEYINPUT114), .B(n535), .ZN(n536) );
  XNOR2_X1 U604 ( .A(G141GAT), .B(n536), .ZN(G1344GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT115), .B(KEYINPUT53), .Z(n539) );
  NAND2_X1 U606 ( .A1(n545), .A2(n537), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U608 ( .A(G148GAT), .B(KEYINPUT52), .Z(n540) );
  XNOR2_X1 U609 ( .A(n541), .B(n540), .ZN(G1345GAT) );
  NAND2_X1 U610 ( .A1(n545), .A2(n572), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n542), .B(KEYINPUT116), .ZN(n543) );
  XNOR2_X1 U612 ( .A(G155GAT), .B(n543), .ZN(G1346GAT) );
  XOR2_X1 U613 ( .A(G162GAT), .B(KEYINPUT117), .Z(n547) );
  NAND2_X1 U614 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(G1347GAT) );
  NOR2_X1 U616 ( .A1(n548), .A2(n556), .ZN(n549) );
  XOR2_X1 U617 ( .A(G169GAT), .B(n549), .Z(G1348GAT) );
  NOR2_X1 U618 ( .A1(n550), .A2(n556), .ZN(n555) );
  XOR2_X1 U619 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n552) );
  XNOR2_X1 U620 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n551) );
  XNOR2_X1 U621 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U622 ( .A(KEYINPUT120), .B(n553), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(G1349GAT) );
  NOR2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U625 ( .A(G183GAT), .B(n558), .Z(G1350GAT) );
  XOR2_X1 U626 ( .A(G197GAT), .B(KEYINPUT59), .Z(n565) );
  NAND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n577) );
  NAND2_X1 U629 ( .A1(n577), .A2(n563), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(n567) );
  XOR2_X1 U631 ( .A(KEYINPUT123), .B(KEYINPUT60), .Z(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1352GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n570) );
  NAND2_X1 U634 ( .A1(n577), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G204GAT), .B(n571), .ZN(G1353GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n574) );
  NAND2_X1 U638 ( .A1(n577), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G211GAT), .B(n575), .ZN(G1354GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n579) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

